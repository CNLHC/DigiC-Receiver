��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���������V�2���{�S���K~��FU�׹��]����ۙ��18P;qԁ��TS��e�mg�U�L��c��Y�u?�!�|�xT���0?�����[.�I��r��7k3��^;\��s֐-P�ȧ���1ez#�(y�wt�N@�fG�_�=6�X�vǙm)Z���;ȧ�4
�m��Ƞ6����*���rp�Z�/���s�,��:z5�t�����.i�#Ve�h�)ϰ��g�fxI������IA�>Pz_�1�L�h�GO�A�y���%�#�5D��	���/�I���,�� K7�1��B�٦-�@�4ӡ�������Y��Q*\�G��yi�=���g������w��"K^������jA>A�^�W�J�u��8O,��4K�q_�t���^���Q���q�)9�$7�i_�y��V��EU]GDl?~b����mȀ �Q����V���
���<>��8��iy���/�\�8S��Љ}_J"�'m��ꅚ��7U���u>^>K���Q-r��wP
 �%3��X5��o��vV�����?��vM�:kl�d�
���EV�,������&V����2J���_6߾]U�)4�{��"���3l-�b�2��խBH���Ta�Fq~{{��r��͙T���ƟZ�8�`�so�ŤK��#�~��cB�16�\���H;�:/��&���o��~]]ہhѹ�vr��gy�F�<�ȉ� ����#xz3�[��C	���A���ߓ!:u���0m���s���S���O�p�8%�OD�k#����w<v��&��q�e�0A�#�z�u@3��U%Fk+B����m!R��؝*����T�9�ˆ�;���̓��WH�<�9�9����5~<�
n���6m�c��[�p��.�CT�u���N�nZ8f�kJ֛�7�k��j�lH������FA�=$d�јH�` G����Fg;gF�;��v��RL���誂�>��&�t�!U��Ջ0�>F�f�vP~��n�c&Du�,�5Q�*�/0����s{Ě�-�+8t�S� ����S�`�c���d���␛f�)&2�����ܶ"�H*��Q��գhp��l�y�1�f� S0���KX����	�S����$>��	��Xf7���K�|�lVc�W��RP�Qpo���%�����Rͬ�T�,��}�?T�4��u7��˪#�m�o��R����q�'���0�z���$��Iʒ�l
�ɯ�}�M]�H����A]^zWf�8��f��dLO���NkT"Q�Y�3����mZX(��&�R� ��^�h!`�mFo*���,�=��r.�+�Ol�s$�0��ڗlC`�]�},��R�cm�Z�y�	�6�\�[ݶ�D��L4��$����������|��E�f�&���-�
�(/l�-�YZ���x�o��1!$�����+ş�J�t�e
�0�q$�	6d+�t���`b���'�%�W��?@�Y������k*dh4�3�d�U��3��B}�gD�J?2�`ކ���Y}m�b(R~~�K�d�)#)H)\�\��:�A$O���S$x��p��6KK� .�6<᚟��+����Ս)����]�N��#|TW���/m"O��j�u��#���Qg�vZ��+1�a�9�Vc�1`N���>�-��P��y��8h�� u˖l��Y\�~�� �Rכ@�5c)^���ϯ`ꕤ4%yJ*�2�kK4^�)X9f~*G�f�����(���>8q�pN q��Im$x���g��Â����F�����k��q�G�X�#�eh.A��Ps����\Z�-CTM�{4�N�k���?��b*7`�}O�G��?�Z0�
9���}B%�w�����\�QI�e�2�txT`D�D�=����"9`�Nd�DX��'��d�Z��E�e�`I.�t�3���x(�;5����"�*� ������i�]eS����j�ZFd=�\�h�>����o�-ւ��Й<��w��_4�B�`���5��rC��&�0��*�J��R��Q�Իq��� �q�\��4��&X� [���͵��h�p5X:���ܠr��ao��:5d���"r����
I.�ͮ\��<d�e#�/��Ω�t!i��^�+J�5
G�4q�<�N�	��@m��g��Jk�7T��/�"�@��jvʅ�(�"��S�%r;�t�_	D�̴+�CH�[Y���kcG�P �l^n�?2�·�?���)�VrD�j
�Ay��E�9��܆�����Ń��y�?�9ʜ3��=2�3SFq�y*��Y�N$Q�s�ohl:E�Ɋ��J�p��ńQ���!��ӵ1�}�Ɏ�`�ҚTˀYcG�c-5��"��$�P ��!�U��%�;/:�=̕�>0%����.�pLs[����b�<���>�~i��W0�f,�_�Vq���w{7<\9|l��[:L��0���p�3��C& ~T'2t��)�8��jk�B��d��%ýfj����ѷ�I�.N��%K��<=�87���L�Z��8�5��&Yn������ų����e�����U��"R>.���Y�@����0����Xi����G6[<�^ �.���(��mp��
Qزʝ"�G|��k�a�O��/��k�P�5������Gix��	��_��;�g�]5�~�z,Q�h�����"�N�:�R�xl�޽�����8=�����%��"Ű�(b�/��o��(:9�?wn�����*���H��r��۞x�8Im0T�X����v��LG{�}�H���>��}є�;sSC����$J���M1���l�z�^��T2x
����s��b-yey�M��ΜI`Kh&��I6�rl�]JԃfI�J���3�*k�k� ur�~�y��.Z��J�� Ӫ��s��g��!$3��h�tVtj���6:���50~l5���-��Ps\����39o2~-�!�b��u�.�h�Ņk�{���GK�,
I��P��Y�~�DW�G�������PfS�V�����Uq�������;��I��7*�����5����8	�2)��_�+�C��l� ���62��G���l�UY�3��`b�9�$��
�X.,�xӐ=ٵ�Z6���3����B��T.X�l���=lǹ=8��|�������x�;���2(OК�S���� J+gM��{!��2����9��ZL�k05�ݨ�0�o�{�y��rx���(�m���"6�!��+f��'&T7@!5�G�'�)����:����!�v;��y0%�,H5�(��x[��Իsw�^׹vӱ=�jK`�o��c��s/#&"����#{cZ����Z|���*CLj?�Ͼ��c�W��uȞhG0�Lb���T&ʼ�5ƻ:	���	�h����جz�S��oL�Uk�"/{�~��?����g�+w����X��5��1S菃����7��k6��� ���YOn��;���:R��|(=�L���uS���/���b�f�e���㲭p�i�$zݭ�����j�3=�o!��r��[ԩ9�/'��ј����o��1֧2�������S�X��K�ZQ�i͈�����)�-D�L�B�L��66��%D\Ȧ]��,E��>7�9���K3���k[qn���:c��.���W�����q='^%��/  j�����_�[ ʇ(:�y���I��ӌ-�o:�s�to�ه3�Ͽ�@��Z�7���C��f��n)�u�Rp\�r��/����̧]�K6�I����mhn��c��[9�yf&�w�% ��R���F���R/�G;�7��g
d8�6o,
�#���#�|"�t'�Cnx[ȍ��㢂�<g���+�,�_w�����5���ͯ���>-��p�kh���֒�[��o�Dq�2r޿�=B!��V�p���	�j��6�K	wx��Bj��R�ƽ�.^	�I.�8�Y�oV\\Yg�|�;�L{���P�Hl�4�2v.���Ń�Mv*����A��A����5�σ���C��X2��%�m�� ��0%3L)����!����*����G�-|�������0�447���O���������楧Dw�~3�&[�U�t����B�=٬�N���r�%~Wp�� @�A��E%�MZ��sGڠȻVR����i��5�[����R�֊����]ԵH �_��C��8[�m,�DL��V��U��(����\�w�l�M%�'��
�O����ݠs��������;�]�ǐ1�E�$"����}~�6����&�Tf1���V�j��||��C��Te�.2x!��� � b����?���ɜy��P/��(~�KF��4�4}�	X����?���
��Y�����aN&�s�UYB��B広'�+����I����0���,�Z��j;����!��z��#�ż���Zk�ԣ��`ދ]�[
��$�@�C��\��Ϗ~�Wk<�O]F�{
��~��ۜd%��r����'��Z�[��Ý����d�<��S�J�R]J<����\�
�|��3XA%s�G�7F焠���}�l�+���-��
�y��C;���Rn�r^x����i�_�i�b �7�y��������9�\�xje��:�!l�\���:��X�Q���h���%Y��?G��]��ozW�PtR�al�m ��pS�����7�0y�]����;1�ԛ���9�PS����n�D{�,��x˧��&�MD�1L�U��F�N��R�mUA3#3p�t��cLafO z�+���y���?`\pD�ww��`���m\���?z�+�H��-A�9ܲ�3�O8@Z�i�t�V:���/}n���V��G^�ڎ�7���1����-�Zr��{:UW�c�4Ū^?��ۤ�(�o�\��"/M�
�E;f�ۮ�W1坈��r��.#$5>cd��Ӟ�i"���x%���Yp�cᯧ��lOOu��J�}p����{h��2��3����i�@����.�s�m)�OoIjh��%Xm M�[ql�vZ�����m��N͗�b���E-N��O���FL*����z� ��P��q&�X�Dr�²�c�����a��,M�`���T��+袢:M�$YΧ�R4�T��� =��p��,�	�fBZ��v��4g��$�����'2���(}L���QM�)�v�T���4FW���$�=&7ß/TO6b�V8�᰹�����(��t���,TB�Ȫ@����n\ၽi��,�ݢ�*�Y�v|�n�껖 �����G7����=fwI����xy�v�?�)���28F�����硰Zc������٨��D��?V/�c�(b�y3����d*�Vcʈ���BA�m�{�����l��١���\�\��9�DE[)��eԩ��yR�r�l.�R7�L��#�l����>�B�(f(�e�L�df���+�O���Rp1]a��cګ������`����5�`m�8�dh
�wE$�ݵ�ͽ����I��U"�  �֯�ΕYC�\�-��H<?6%Q}��X����	��h%�e6N��>5W��f3�M�\�tn�Z�h�v�Ԍ@,�q��Yu��"(2��Έ%�MO���u��PG���-����4�`̍��k[,����� �-��eu9���:6�#�E�D���7�N��qSn�8=�D+.�b} �L3���t�z��}/�^�fé����l΄
%k^��6��	{�9ϒ+����&(ck��� ��HU�Ua�!�x�_I����"��uz�\�z�Λ��d�5��צ36�46��O.}J]�] ⢷�7%�I�5��q�@�|5���R'd`�'%��Эn�*v��3�[�j������A��%|!�H��������~�v73[34��HcK$��'�:c�-�/�5�2�I-�����,�	�m[��H��\���ND`JC�#q�?�ɳ�_�ɍ��ب�D��lȦ�	����l�J�m'�<Q"��|0�s����'9����%��@C�y�Y(��������Tl7�Qц�	�
�y�E�lُx�֔|H�]Q2F�ğ����d�DrI�%�Ȝڱܸ���jd�ْ�$��Q8+Nm`��� \�C9��~��Z��� t�

��y��a�s*m���w���g���}+h�<	�5��V���J�a�,I!���pZ[�x@-�w��'\/�8�ͥr-2����oL"RN$yϽ5�ɎO��V�1Tq_�y-������!2B����@�#Isl��Eu'^>mt������{6��!FV�!�����DG87|_�m3���<Tb����U{A�h�KwfͽI("��"�^P��9��^���Y�'�s�!�k�-F�SՓ���+�c��O9C���J��F�����Ô�K3.���6(�<�y�9c�������O�q����.�V�����)�?.N�� ��=P:�U��
���=&x���v�Ѡ	T��Ҙ3]�{����-���PI���޷tzPKиh��}�KYj�Ŋ��)���o��V���0���_~�aWx�V���B�z�{%��<pݚ����P+�g�W4�Bh6��XE�O���>ݯ̇�I�*(uӿV7����Q�^�}F�K�Dr׈�"�O�5G�}5�D�1��9�ī�?V�f�-�P\f�G�b�m�Yu���AJ�h�HH�=�9a�׏�&��C_�L�e���NQ���@�%2ҙ�Ɖ����t�g	�qE�G��:.�V��u$�HyO~����U�ٖ���5��Tᾏ�WB�FW��V]r�уw��xq�~�0�{���9q���Ud�����}�I��������쎲��6��K(
0Q��B���05W%1��n�y�Ӭ��� �6$ؾK�&P##�}����g���iLzK�k�g͍М�X`�O�DV����|����0��'7��I0���i�����cؐ�N�`���%�M����,�&�TV�2@��ZY:���Ƿ`x$�E볕V�5�v�7e��H��'��;㜔*�"N�_Qp��
0��с�1ȥ9��� �lo��T�*�T���O�tI �J��S��<d��
�ۅ�/��ҹ��1�aoZ��?B��bק�D�'� ���?�Z�9B
6�������-��|�N�^'��{;��o-@aY�[s8��X_[YQ�{�b��4u�0�O��UQ�����/v�U��AeX��f�bC��pv��[.�}a�yI�?/p}�A�����v�����'��}2%Ku��*9�ş؏��՞���T>Oh��9�緛�$�ϐ �e;
��)
��(�kY{vicS����T�y+@Vq6��ف��]+e����kJ��n8rYsv����@&9Hw�&�tǈz|�!Ϥ�W���Gح�m:9�Ҥ
<l>=�D��*��QA����SKɄ׆��7�M�xѰkdJr��Z
5��Z�>�����1�|_M4X��vY
� j��!�Պs�<���ɄPh�܊"�K:�n��BO�Q���J9�]�������a�N�M�ɂ����P,!d �+�7^����I���O�c.c��3�/p��m_�(��;',i�����m�����Z�@��Q���T��gZhY�w��;IT�Ebvx��r��.��Y1�}ܽ����8��_��؝mSF�Xa�����Q9���L_re&A�����9;�h�;�jd�	A+,�X\�b�h�B�����\ɩ���:	G9HD��uC��خ~ߊu�$�6��v�)�<)�� w�1n��`^���S��H��ú�,�,K��T�l��/�V�����ZrJ�c^u7�OҔ�R z"�3�A �HWU�by�mn�wmE�"F-�t�?�����5�?���	o�g��ߨ�����&rw���uЃu+���H�u5c�����-��D�5z_�"�����(.0���Q�O�pM�U��\�t�l􄮞0��d���P5�}���	Wcٜ}��q�K�[�F��J������k��xفX	\u��=�'�QU��u��	�v��I
�2���y8UG�o�0���\�����M���'p>$:!��N�c��ϱ��/���+"���>WMT�-�U��у�����we�w/ͤD��X��;
c���|j`����T�E8"������%l0�JD�9i�v����J*�Q�1\��m"��BR"�J�=��(�A|/������#V�)�����(�Jl�OY�e��%2p�+��#�e���h�Z�U�ʂU����㹱��|���,`,�\��J ��%BD'�w]P/[�o� g��v����!�i�=��Ig�D͞j�y$ZL��714�+'��*פ�1X���(:ʓB�'�@��9�3t���E��{*�>��t0�I�p��Kgm('L\�V�֫�U9ηt�7#��k�B�e:�DO3$27
<Tu��I�&���L��L����VZe�̻�
u�m�z�:V� �̚��ʆ�$W7_>&���(JS����D�|���į���¼�c��#7U�å���_�X�y��}��7��E�Q��e[�=�p������?]�s�m��G���F���tĭ ~��ؿ���#����L�&��bC���|l���U���ؤ������i�e�ijP*�oV�$d��Yހ0�V��F��i�na������>��`~=r�]�b��>DW��b�9��P�K�}e~�W�8PC2	��W�V�
Ҥ�V�t�㴝�J� .��
���j���!�{b���|�Ì�����264~c潎nry��-�vó��2�
-�U6i���M@������<�_�(@��c5�-M5����n�fR��Ze�`���fe��g����~+dCv�i��R�-����	�]���q���t[��1~���"��*:�����X�M,jw��"�gDm����$�M���_��j�)����>�ldRR�?M�8"��dq�\+�S�,�x����槾㺢�G��L�i���v�Ao�ޱܭ#����yo���� �x�n�Hvi-�ɲ����X>��^�謖&&?�c�+\�E
.�o ���q��Yp������Ŧ?��c�{�o��\�� ��{��pm�}�9�A[��m������S7�l��]N9Zݳ��ɴ1_Rx�>[��<2<-�{�!]��d_������0�I��^���X�\zd��.i�.�/f��X?�-�hO�'o��p�F�D��@����\޷u1����f哅g2��V�P��L����.��N��Һh�3-$��y�)10���!1,�]H���" +��P�}���q�����������hD�_�D�qrb�Y�_w��!O}<�2e��;�|F�b���-�l���Ͱ�i����X��f�J�
�*�{�ٖF�چJ�ѭ�`���:��+_:u�{/BA���&���6�
��8��3�;�[���=�r8.c�y��'�����3���֥�[L��&]	�~���.��0�G���T{.�dr�d��	'"�@Z�\�wFS�dw��u�
t[g?���l��B�w���zf�A�A>�O����#�Pe"��=��� 0 |��!�5�������7���.zt�a�4o����S%�h�*�����_K%�N\��S�5n0w�8���SY<���it��,��S���%
]9ώ�|�m?9Vߠ��1�Z���dX�4���a��v������9�ic�9�O���V�tƹe����ρ�MX�^��i,6�fex�x��\:���=��n;	 �֥�8�����"S���K�?,4�_��Â��vo�s�Eޗ�K����y�MIf�H��|#jʹel�kb6E��P��uU�JW��iG�}=ֻ���QCNY����(0����"f9�`ԛJ�� l]R�ʞ�-�1��#���s]֥i�C͆�jl�Q�ԝ2= ���8�h�"���[��O+Q�+�W%��;�><�G�R��wp� XK�q�0 � �r��k��c6T�����-�H&o��pM;{HL�N�SɎ.��<�$�Jn�w	xm�1��,�UG��G�kr��D�z�O6�(`˜�֙�[�b
l�<&���A�WIT�k���M+�mu����6g�E����} �S��},Q<|�<��������v�w�����Ym�9�0�$�)�|	��i���~%�|�W��I����h�ob~tgT�Dpb��
�]|��#\O�zvU��ʰ�#?8
T�gΣ�̋��>��PÞ�@�Q���$���>�4��L�Vؗ�q�n<��U��tU��/�(�1���da��VD��4�"a���'���]��Ϩdn�)�;�i�X���2-�;�����X��@M����lA��_)��X��U���J�Q�0��6������l.z(E)Ud��48o^+Oz�\Vn�{�	�8^����"���j#��[O7#؅��?st�C��4��Ü�5
�{+~7�I��~_3�W�5R�f�m�����S���)��9k8��|dҿC<5�Q&}Y�-]࢐�!o�`f��]����7S�����) ���[=Q&}9��} ��xy���w"_S�?�n�<%��y�PB(�s�[��+
���02�Σ�=ͻ:ͦh{U':�t�C��t�y��!���@��m�pC��x���gS��keK@�wʏW���w�rf���E�*V�0���A��h���ah��C�3ƿ�l9�t�l$��O���L���ל����
b�Tb���Յvlt.1�����S���j-G�6}��T���sl:ٕ<-�5m�&��u*���DV������v���I�z!qvNC�P�KΆsE�ce�ju�B�M�v� J�f�D�q$k�}��rK�Tǵ=DA4\'��!��i�I�]��D$$\�I�ӰN|J�.,�
G�+�۽��O�_t`�Ż�ٻV+��`؀�W�G=zՂ�q�uJ�'y����OҦ��#O�����~��Ԑ��jy�x�-��r{���2�F�u�L�>G�l�K �=E�>M���Er!�E27���pǡ;g����R3�ۙMz� �� ��)�5h�)7c}���ha���^�;�c��3
�Ķ;��٩�g�C�	D�9T������v�,��gJM���߼�_1�]�1p�%a��YDwFVS�g���,97ٲm��4X�9P�>�+�y@-	�{����k"_�o�M��X�uT�#������Уզ7��C��t4��q����3[�#=y������}�d��Wr55Ξ�������ݻ,�vI4��u_��8�X\⥓o�$	�g��Jɚ�놚�L�ar�e����
p��@�@t�6��TW��#\���mCK�"UG%����	:T���|��f�5Z�M����,���*��O�h��g��Y|�)_#���l�y,r�\?w�Bۀ���}죌
4��M�Y�=�s�01���Dz��!jN��Ul�`��~����Jm����w]�Pn4�絪}J���B�j��E��A#��@MG�^�n��~�0�R�ɾ-�J�m�� ���.�S�c�y�2!ʴ� `4<Sr!Z,KB�]��T~��jX���۶�2I7F2ef{ts���~�)�~��p��l_� ���� 9��xnF�3���}���wCzh�zp���$+~c��xC)��o��~츥�2�娢��q� ���UMh=�[Z3h���3�̄
���7/�x]?�A�4�fs��HbU�c�vS�ٕ	��g��,|���P&~��?�G�>���/1��k�8(���α�`Z�q���8Zb��w%v��g���䴉����L�WD'��|�����&m"|�l}����&�Ĭ�#�ۥya$�������:�muO�:ٷN���V�&���[$8d�'� �OT��+4M����E��td�{ DW1қM�Mv¼ W[&�e����
O���O�B��� �� ةB[�w��W�E�
��|D����K�)�/iSR�X|��㖂�ėF�3]�R��݋��U�� �{�W��R�)�x��z��Mks֌���s��������ˡC̝lHa��ϜrcFԂ����%��r���lO���3��[�Եs���6}gf=k��$a!�����Q]�[��iz�>���U�5��$עb-�{8t�r����72�s���G�ΐ��?CE��T�Dyr�MQ�NP�����uBZG��Wv���κ�F^���وd3�^��m�l�(�
DƄ�[�3{��qE���^�9ll/�#�Y2a�J�bO�]��ڥ�fq��s{�!���n�/{8|.�}-w�ۣ�\�w���T5����Ux���-����j$e)�p��z�����T�u�����O�x �)e�2�g�M�����%f���Q�ݮ�y��"2������^����^���(b�tJ��z8k��Zٮ��܅ikvqA1�ڣ�Hu,��j�ؖ%���*o�H�����a����X6�:�l����`=S4�����B���c?�ފ>�i�5���u��ir���K;��+� �^���卽���L�nd:�L$�AJ,﷋z2��A*<�"ج����{6��9ѥVB�M
:��V�?uUKwqH_��,�A�~��Cm I�.�Z�FW�ȸ1�=�m*A� ^e���5H��vWذ��hy^��5Hy#*���z\;w?��mI�ڼ�[�aу>�4�Ȋ�Y���ttH�)�$q�%Bߜ��D�t�txO��?R�+�����u��8�e����b�F��K����Ҋɥan9@ċ3��̘e��	@��Ϲn�d�}E�d?s����r*�I��Ec�~���`'��p�|�� >|����sG?��C��+sVD��+��!�����Ah�(���P����4²�[���#�)��Ј�n���εֺ�/��L�MJ��c`~d�Gfu<�&��;����h��'�}G�!�[�W����W=6��pb>7`DǪ��G���u�����'?�\\(�I�`���	%������c&$�P�V^!��{T�mK���D�3'�!�5$�ә麌u�cӨ�W:;�e�����(~Ѳw�T�W���`'_�j[���riR���l���*���7X"nݔ�xÝ���.>R��#HL���N�	���ĝOr�^��*8��e�` �7��k�Z9��j���X1���p�ȄY�7P
TU*$h9D9��K�U.�#q��4&^�k#|�oQ����idل�&�J���E�qȣ�g��� �*�Y�;'E������Z�i���4��+������Z�OK��7���F= �������P!�pm�Z�����rY����]�Kv5 ^���UG�ͱ�؟�mQ��8�p�T>x�l���$���M]6�Ct�.�cY�������s��ճ/j��1��m���-� ����k[d1�EI�]���k�ːm�Fv�&Z�P� ��:��{�ck��C�/D���yu������L�<-p�FaL�72B;���䉚i,԰�J���`��LH#�X2�-4�m��� fk�c��s��̃�X�V03�_��ᶐE����J^\Q^�H�B8����p����q�y��
&W��W(�["�`J�l_@d��x��{#�G��e�*�u�Ѵ5�b.�m�3����m���w!m\�\=���^%
s>)��-*u���U|g7l3@�IW$�ԅ#�np��ns(�f�#W�1llg8��Ҏ�?i6��I�����8d]��oV��q�J1�I���3��t,�3|`�3y�^�]����kJI�X��	��I�W�&��E[�l��P�H��e-#�8\�3Դ�WF$�Γ�"��zu��һ<�p~�����|+l���5���aN�1S���Q�$�0ڢ]�v����C9���`�:5�������=q�����c,�|�'��U1-L�f��x�y�Ŗ�e}28`_�O�����7C"�����k����ʣJ�u"n��w�8r0����x�-Q�xl���8�{�xb_܆{=_��|Hƴ��,7dO�t�ۦ
��"�	Ia^܋F^_�Nc{����̘�<@��Z��@⼋���v��:#r3�2s�l"��O�p�J)4��	Z���s�I2Ox�$H-|D(#�úJ�8A`�Sdm��Χ�Gš/����[��_�B(H5��bj�DCaշ�$#����v��>{�犓��h�o�f�"+�����܆Q!�%Q �W��FV���/F�w ܲ��`�̚�,>���F�s��;�A螂�]~�,��J5�{�R� ���83.ͮ�hL(=+������R$8�&�[� �ų��~��>�bȟ�'
�?��gNR�����po�P�!M�Ɯw��!�L���6g �
�;�R5;�*V	y���xT3<��I�eG������8?Sͩ���1�����'����>2wL����Dܯr?z3�$U����,vR
��`��%�!X�����xZd	��<�2W
��;	�P�hvwE�O�R\Ն�rj8̨������e��.��<+H-�/L�BD����I�5Ⱦ��L��
CN}��h��PՓ^�����������eނ�Y��0Q��J��7�Ջ~�V�]�������B�Da�y��z=���h����&~Ol�<�����[H��E�ޙm��Zq��Of����uW&6����Zd���J!�dt�� � �����ڦc��>�Z]��JL�Y�0rF@��8.�i���(N3�e:����C)��
���H���fl�uA[6ҋ>h�Em�����}ف�d������g� �WeDX�7PA�p.Fe��Q�%���W{�%&�Л���U���a��
-��f��ns��r�����iŐ�f�	�Ƴ���l!��eȮkg196���}r��.��_* B�8Ͷ#c�	�
�
0�E��fI=HнawK!��LJ�N��>����$g�D����=��[_���$��v��c�и_}|�.�DG�묭Ԣ-����pR���P��g�R8�c����T5Ҍ���>���)�U�c	t�����V����9i�C�o�>{�|8�9���� ����Giܽ��'c�^�����BE|���j@���5"IWrP�烳=ڡ����7<ɨ��m4�aH�]����%�1��,�
�^L ���NkD�&V��0�����4ye�X�O��IxZJʚ%�Q�B��djKu`��M'I�fP�T���2�1�h]fð�Q��IN:9�|9.j���P�]�b�s�p13��`��ތ�BЯd��#<<[|������d{)G�����n2��j�f*F�kQ�-�/<��<��az��)ɾT��t��W��h��f��#��d��nU�5; �Wz���`���
S;�y׮`F����`lLuQ�|���u|ʀӵ-��¦��N���F.Ɇ��oH��p�.��[�� O������� R^|E�qcj0d*�Ά���z���
�CG�Q�#�(���>�y�%;��G���0��2)�l����s%�-	�h�Y��@�(�ؒj�k����p?kƯM�V�En�ͺf������	0uDݧ!ç^y���/���E�j�t�)��0�`�'Q2�Υ`��ڱ�\�2�[}���]�����,�=�r�m� ��VE�d�&� ΟK�bmӈ�K>W$��|J�y-��/����w�n�09*6(s�lD�u��n`+eH��a��Q����/��&��>�KO@/[��	��D�'&�B�x�[IP�~���m��‐�t�6��<�������O=H����_T� �d�`���I����8����
`]���I	S��U����+t4�����%0n�I�$��z��<��{�K:�!M��à�3�c\�9��,��j'y{ #������5��_ҧ�y�\�9�A�$	�]����� E�����1�d4�$��h��"a�p��f�:yQ5�y�5�@�OW�V�x�|r8��@ԕ�l���t�Ŋi%�r�ݰt��*l�m5m�(�Kµ7��p3;���l����SR]8�4$47��t	��'l��O����X
������}�6��6�:m���� g�i�y�M�F����I�6槆M���2#��
"�A�����!��jٖbV���2��hx-��l�C���$0�B.5q4Gp�I��` o���y1k2�����O�x g�ޗ	-��C "4o�CR��_��1����9lQ�׷�P���+��E�&�w��aQX�-�$�ض^���{ҧ�bC���(rvf�(-'���㲂ִ|���p��-��3��/��l}
�l�kwLA��,F���΋[	7�T�&V�p�$Vr;}���e�����{Uq �V�ײ���N�m��A�}B-W�5�	�j
č��J���j[��������t%���X�7�嘿��D���6��;ČRTm�QM!��2%�A���y!Oy�j�R!(�(7 �;"hm��vҘ��#��;��|ť���n�׉�H&�[O-N�e��:1�1��z��"���LtK����6C,����y;�Cﮥ_�*ex�)�)G=G�����ah�+Lo���txh�F��Z\Km����ny�a��3�2�=�!�
SS��0%�*+�/A�bAlʟ�,�=\�:	|q� >�H�*���q�%t����^J<�撮�lX
Upp{$�T�[_�N����rN҄�3��K+P���8�/�O(���,����`���m�gU�{����h� ۄ5�ן���ЯZk_�=,��Vr_�]{H���ןS��WPWl��T��v�]fֺ��-0G�B�D>��ZU�p��4x�,� ٲ�eN^��w�j����m�ki��}�̃EU�����j���)U�JV�ݧA  Ǿ_���1D�;3bF���*�r��
��d�sRQ@�<��`o<���2^a� �2K��$�z`�^U<&�mG_�_ ��N�6G���8|��y�GL�#ϜB�"n�d���\+��(4�	��
IA]:��L3`@4$k��ˍ���MG�Up�޸��y�Yw��&�܇`��ε��$f�cp�����m\��WFYXm�q{�ג�*kT�+F��H�U�QY����O���e]F�6���tч[)��^@A�C�*p�C�e�&���ACn���g�b��J�������|���BZ��c8����f�x��~���4њ�%�F-� ]�s
���|�͙�a��_��?�y���gu#=6�6n��g_��,B)��Q�8��?-fF�$��Q�A��O����E%~�r �#�-ś�a�\���[�C�U��z08�"�``:�EL5S۞�W��{�����ڏR�����~�	tG u�%A�J!�B�7�����1%�:�����S��|X�]�4�RF�5�GW�p����!�5u�O�xP\��<W�H��+�b��;AN% ������-�AN)NY������}�*d��F�����Y���!$�J�˥�~@�vS��)q��/�>et�)jN��&�*TD|K�TE�;?s~��E
���-�v�q���j��f���ly�?'�NpV�Y2&�TD+�E�,��nj$��,��O����r��}�b�Ŵ���u����W冷�Cz}�c�`D�{j��Z�M��B]�F�Y,��´QNx�>ˑ�8e�Kq���}`���$�%�q9�	��z{
�����9X'Q�fCè-�	=� �W\`I��R��[v�T��)�������;��+]��F���4���3�ʼr�G$8�q��ݹagypZ�0tE�(7Z;�hE"�iO����s�D����Y�:��Trkџ�B�2.�7��Fb7#y�.Zm�D��\A��ol#{��&�cG��Ɯ�Ȍ1�O�P8AU���E1�޶E��q�m.i�3M�k)j�����,!�~	"2�F|�Jy�F�&� ՗r>A6Gr�����AE�׸X�<��!�R��������;�a7aeL
RU�{�O#ȝ�����㋜X�^{S��˒�c_�'��Hm�2@�h^9f,�2�d��oL�$�����O�|-����T7��,A��x�2�>Y��V\��R�=ԅ4)1�r��Hc_���]"�"�^\��Ge�747��[u���gꄂo��������l��Z��X���e�mЮ��l��M�p�y�\ث�Rj#�����@E��~4D|��EPm��.�;e�|�+��2d9R���4�#-+�k�n�U�Ҧ.�F�QP�J9奌���Q�a@Tʪ�`�s�r���Y��z!���5}FA>c@���春����&_�G��e�(�R��	2�p��Z��1����˧���W!���\�@yq=��mv,:�̱�Ç����fd�U|+p��s`�����ⱱ�_A�n3��Hh����k�_d������F���)G�g��#��<9]!wډPW�а\���nw%XXp]�pѯa��a�"Qp�oi��@-vI�Z�65�c�Zэ,n���C��G����]����7��=u�ܳ�ܦ`�O_`7�!�h���_��鰤LG�&D�c�� ��� %K&���T��_�c!������qysiO;��S�wϻ��t��-f8����,4ܜy��������2��b���j����PFQ̕���1�6����PG��jR�n$,�蔶LnY���I�KnMm̢珿6�����1�kJ�|��u�x��U7=2"-����-������B�~m�J��[>��Cey��.ٿ�Iz�9J;�5F��i�KKh.Jv�X^eMy���������P����K�-��/H˘c�h�g��r�[w8�#�.
$���ϡVTM<��%	*D��&g-�3�+蝾2�{��aޗ篕l��O��P��*�e8�_v��(P��ĕkw��b���Uh�p�I�G��2��zz�u�p���n��
$x7�ʐ75'�CUD��,� �Ǖ��g��!ϖ�'K���S�$7�]k0Ι��7OOQ��dD�YK�N��j��#��z��p�tM��jY���������_Q��l����5L҉8|T����t�Hr�O0�ܩpU:95���:�>�m'�Kz2˿��Kti�����{rɀ�����q&$:�%�1+�4�X�,C❂��_1+9�����4�-ٟK`~��\��3�����M�Q_�C[|�f�ZI�;MȦn�S4������U#�TT��{8N~�2ͶG�P"��D�k#�EC>�נ>����9��ـ032�Ӷ�K�b�����)�U0��,�B4;i�n��!S�b�V��m�s/�/��.���K���g��\R�ד���N���n�b�ڢ��_����D�X�X!t�������2P�)���e��ڱK�tMLj��hʹ�Y�9wI��~P��&�-�����N^�l"�S�Ң�T~_gدr�~����k���Z��a�_@�Pa��t���"q�S���WG �������՝�(�A�<Hrn'ڨ��y/�a��
3�zV)�}0{L�C���'�ȡ���/A3��ڄ�*=��d�s,A���_d�����Szd��]��5d��G�������zF'xsJ-T��,[����<(r ΣE�R��q�*hT1"��6�Bz�9�C2��֖���-�?0NX�'� ��7���8ͺ�UŖaв�E�7���AľB��^o=aEY<ۀ��U}v���b������ڈă"���ꥺ�ҳR������:h"����T{Z�@�l8�ٛۘi��y�Ʋf�����j(�y�x�0IHyYN��"��q(��I3�$Ц(̏ D�i�[�~� &��Vf˕��A�t�]��c�2�g�`|i�d1�}����N!2�c>Q�7.u����Zm��Vf��?IJ!�n��Di�� �������m�hGt����4D�_�q��{�#+���$%��
�fk����.r���	����fb�U[ώ��L.�Qn0�����1e�l�U�������Xu�o]0F`�QoG�"&�����A�jZ�s���P��*��7�S��Lj��T :����q[Y�neHŉ�s>����9{,瓓���f���
~}�qwY*����k#Ǖ	�(�� ���6�k�kC?V��������5�����K �>Q��w�dͼ���VH R&?���0&R�����ȩ��5UJ����b>g#?d�{��Ț���2t$���G���a�璲�u?T�]�[��V^�b(��z�5�w��M�%T� cR%N�Y|�L!*T�f9}0Z��۝��N L�[�3�
�Ӄ�s?����M�iB��o��O}�ND����%���C7�w���N� �@�ާ-MLx*j��*:�ܛ������q�zr�C�jj���l���V��ۛA����o��ss$� E��	ic�VhK��������R7Y3��pkd���n�N?_�r�$!���a��L0��^�4
z�1��"�_��y�s�ߊ9o['��u�9Ļ=+rf��¢b+55t˷���#�e�짅P8���@�[xLe5��1\����ew�Bq�ħ�n��#�����.�Gࢌ�8r�!=5Bu�DH�P+�)�䛼�e�CR �+�z�� �y���o�N+n;�ק%I�Rl�b��(��eơ~�h�i�O�y�bm�q��\_Bo'�z���%�g���Yٔ]V&�,"��$��mE��eHt L�Ӿ�� 8B7܀�嚊֦'&)95��=6�r6t�=��R�4LB5o��tlu����V��4��_3D��[���n&��:��&��y]�� �����0U�/
@��>4���b`��ZƬ���[� "˖���X�(�K�h�)���{b��u�ʿ7��[Hg!~�iF|�e��
 ���}��{֣~��>s�xo��E{���&g(Ƭ#}�z&x:�_c�P����8� ���VBE�fk%ɪ��${�#7�B�!Π�v:j��쒂ٵ�/�P�C<����Q6v�����o;Ԭ�?ߌ�R��ؠ,�W�)�e3P���-�5���F	��.,5�ƀ0��O�@&��3�@�>�v	�q&�UD�]XW�:�X�w�����^�����޸�����E����i���z��6aڟ�)�P�G^j���/^Ry[�@��y.i����la�R#.�ʭ`�1Ka�i�qw�%� {	��}��7���7toݲ؊��-��z?M��	�|u�����o��)�l>���6qV'%"���zT���I{�oA0�)Q�[�S"ۇ�>�n}�l���꭛R:�����}��ُ�?�A�Y	���M�@���i�F��;��j��J�ji�C�2˞ߏ��> ~ϧ��ϩ���GI@���p�yU�T�O�3w�Ay�XXHW�uC���zO����򚴸4I�/ ��.�!4Ґ)��]C�)�=* M��V���ظw�����%c_	4�Y���X�OS�,�d��Qf�/ց��bM��4��&bK��~�ZU��ZX��$��D���7T�#H������%�*3q�o m"wѦ�L����`���9b�8��{��r�͔%�g^�����p}�?"�/}O��)G[Z�=��X�V�/ʠ��Y
�(���+jV)����>�ή-YU�\�I�=8Ya�� �R͌��	X�<͑���s�D@��2�4>�j�?dX�J5inE�þ�LRC/n�S�CZ�џ�}�C��������)���T&w��@�f0��h.6��� �|N/2��Rj�`M����(D$�_�5�:iء��x_@Nܦ�K�!Te�d�:����y���Q$̌��[crm�*�&xIiA���� �,g��|�74��λ<��6����$���(V+T_|�)k�U�����=I�͡�J	�g˒�Zf������l~b.Y63��Qe��}d��*�T9Y|�J�+��5��W��+�	�4����E�`�F��z����^M���ԟK���a�8��h���U�f)'G�{���_���K�q�kO��޾fC��� 4Q�e۷��ל�� ��2M>2�;6ؗiW�g��{c�5_�g�:N��ӣ[��{�7�h�@ׯ�8rP�S��ve8rM�x�Kչ��_���D�o�a>^u���Cc.��hb�9�y�]� �O-��$�c�d�H�߹�t�#���f�-�|lH��|��\�XG�͵v���S�M����t��*�5�����B�p+p(�E�b�ɢ�D�]���|����	�+����!��mA��;d��c���W��T0�Y����V�}��M�)N(��n�}������Й/�
�Drfg
�	�-A������E�ϩ�n�Њ�>��(���"��^���s�
�1�B������� ���SȢ/�_O���P����,�eI�5~����.KN(�B<�g69��"�d 앇ie|�g�6���7l�.5��D����.րE�Aז��Ē猠�'�gԤT��m�0�6�,t�N���T!���ק�!���J�SH�/>�]�r˥��pӛ���e��q��C��5��>I$ZĨj_$�ײh�V��Gd��|�9�7A1���Ut�$��9�*��N�XL�4a���'^�^+��T�-^]s���`�|��s�3��藙q0��l���csyw!�3<���Wo��;�����n������ն�i��6Y�������܎����z�iW_�y��,w^��=��E)_��N�*	�W��Y����d���@�S�b��)�]�Y��S��&=��Q8�Df�&i�?�ج43�W?QTF���/������h^vQ
�ӓ �lӥ=G؄3'aYw�ߡJJ��(��=�6�L�t��N"~�-�p�Ũ��	�����|�F��-�k5">ц�9#i�㑹x�|g�uI[�<a8�
��ҧ�����FpoT�+�W�.�r/M��m|��R��%'����XpB�l��� f��Q��ǅ�O=��'|}�� �iW� �|�04E�&
�i����`�����g�/ ���E�o��1�*5�?ª�=�)t��Cu'jE��*޷6�
hG��W�ONo�lS�c��ʨ�/e�ߺ:��/�V�ܜ���n�D
��M������9�Î�{�������i\��a�� �	�@F�a��f���qo���m�<�D�[J,d��Q-�s�'��y��I�.��Ǘ����%[AE�EL�	�"k���5H�Z�p����������5�^�Ò~;~�OJ5��D�ё=���*\��m�k��,��V�a'�B�����ʺ���3�h�*$%�Ci�F6�[2���w�ۯoV�F F�r+m�q)PLL=c���e1C��7�˚�]�j��S���%k�/�DlɔZӡ;�� E^KǙ;v�G^��}|��l+�6��l&�V�x��n��R*`�6S�}�S;�t��0f$�Eq�ǿ�˩����CC����ڔJ�/ٯ�9٥(���6m{ H�MAZ̇�h�Gؠ��4�b���
Gn	v�n�����;-ۣ3Q�j#k��#��  n�4��y1|���<�¢7������9�c���B@7{P��q�q�-����6J-�q�.�,��i�G�z�[{�4��9�,=���dҕ#��z/nN(}^&��ʮ&���$�F�QFA���&�X��~�HѥM�ғt�X$���ξCe�}E������[��Są/"Ҿ�cj�ڧU�|j�4j)c���İ.39�zu����pT1ྐ�ѥ�(-|��F^���)4���5�\�d�. ��
��۟��C
�m�.HE�NپX22�<QCӐ�WL�>�Z}�i�k��s���#��5�J��p����1<���)Zj��<�ɒ�����sW/R�GK�'-��dç:���yt�#��K�4m�b�����P��S�W5g�[�?%�n|P��oY�6`d��U�q�}QE�X+2;��9�Y�[&�O���(��`�/�Kڅr�I��:�?��댯P��9	q��;�P=Hr�R4P0��zN���V<�H5���r��5�$^�;5oH��k�x�`�X�Y��(Vr�͒���a�$T�:k��V�)/�m]���g�3c�1�:G�� ���p�!�R�_�%��}��'���N��*��� ��$҂���7y�7}U�9	���gL��������;�?�+L��4������BQ���\+V�������~��_I��wJ��5p,UY�����-�O���Ư��"z�L��v�����/7������W.b͵z��/1�&�5Q1�f�e� �`GF�N�_u����3)�ȅ)-]!jx;_.t��1� ���C��4�x�� ^ �QYOb�ʀ�G�,�n��7)*��s���R�Sh�CS��c�ؖ9&�࿉�'ë�;�>���m�SK��f%���p3ƞk�S�΂����&?��z0["a$ZF-y7f����J��ڜ����Y@֨�R�����ŋ,�ca�=��ibg3C�e�
1���bT�=b��"F�ݡm�z@Q�Si0+P�%�G�{�bQ���ڝ�·t����y�[�Wݟ��{yɯEe{��ң��OQ�	]�]�qxX��*�.��]��`���CK6ٯ_/�^u��"$'9k,>v�.b����UdtcϘ�K j���+��x+ �f[�i��p��-��n���޿5D"&���wUۀ���6�v��ck{q�z��-���W*�fn�jp�`�d7���
���ĝ�&S�H0����ێl�e�UA���1C��`q�N��ĭC��(�P���͓��ԉ�yA�Z�����w#�lsȆ��
�U��J�f���b�s���!&�-������,4��gC�8�K6��9/���6Й�PhSdM k�e$@׳Q̘� �0���9�zn���{����7�tD���d�I�*"�b7�b5�"+v�˅�~B�M1�X�%��?��?�0ٌR�nT���e���|���J�_�l:K:�9�x���2mT*�+D��/7Ěٯ�'�?���#eIG(��=��[�L�|�%d#i��^��� ]s�K���º���>�w�C]�(��_�F���T�e��Ϲ5� w:݅�B����Ǫ�ט؇��e[
�j�m�� ���D���3u��b e�Z)��1e�R����c���jd	6+����� DQ��	�׆�t�v�����<�H �W��ΰ����r;8o��4P��Z��q3��>�0B��@�0Gu�TO��s��h�)!x�}AcRq:HP��i-|b̩'f����J��M&Ǵ�),M�˰�J�8�~*GjE�蜀�5��@I��W4�(U:��i*��c:HE���0`
m]��BE��� %����_@����&�"�*X�e��}�ߧ�='}Y@�aS����'���Wx5���G�5���l1_<6�䩗+�6�8��x�  ��&>��7,�zP��_�,�q�=�F �ݽ�-d鼺q�A��K�b��W�ꏣ�\����$Bp�_��]����V��ӠMo%4�#	�W��H�B�_v�N�0ŤH��2P(y��
Z݆o���͢~�� 0��ˆ�*@I�>��'���f�$e��6�m_���¹�(YQ�e����wOa~��u[z�A�[J���Gw�}kbe����j��V"�X~��*����������xHΌe�/� �af�0%�.4���O`*v}�*���I
_;)�鲉<ɱ������@j��ܧ��z�gY�9$?�"D	�������9�Q�ZR�0����`����`F�W{q��>��
K�Xj�I)�5*�!��A]vx���c _ha���T;�p� }��˸3�f5XW�!Įi����
������l��#g��N�u�}v֐Y�5R����Hi��D'����e�<u'��Z'�f��H�'⼓�T��jߦ7K�[�����U!�*L*��P�|n`zH���/�;�.���JB�A�0��έ&v���fnB0!�A������H)��H;�ߵ �?��z�>\)���I�u�]t���y	^u�����^7>�և؝��u��eV-�|���N�N�����bW������[k�gu̕�6��Z�����&�-ZN��O<�ބx�\��bw�u����ëS�7�=�����pw�(<� L;KG)����LN��Q0�%D)K�	�<2N_�]Bض�)`���˾�e� ��ifaU;����9�����~I�<�\�֞�&�Fr�����4~�_���7���H1!#��JKT�*��1>&=^�%�U�6�t��e��V��1�^@c�ݥ#GS�!�{����Ջ}�M�H��&@����0Q�ۍ���G|Jz�#WVMw-πu+��S�$
�X�8V,���x��u>�,�#��*� ���J�ЋA���'���T=fϤrLT���mg?&�̮ɴ�s����i�5W��1�4���Env���
8�ǖ��	Rrc����
r��.loӳ_
�� V���Ou�^�������F���]�IȲ���EM��cۍ���r�2-��p��w�o����-�|G(vϙ4����m�����0�=�p������Q3�AÄ���'5�-8�GWn�Fk�[m<�����>`���v��<�~R��~����-,e��a��J��
q,��3�Cf3��z��xg?j2q8��Y�]������E|� ���%�\��<H�̟N�T��\�1��d҈��dӻ-��K%�D]a� � ��ů%QY�iQ �P0E;�L�w���^le�."�����i�V�a��H}�;e���b;�V�"�(m�X=��=��`N��.��#�!G�D(�b񍘌5m*"g?Bs�����F��w��-��<$���:6�}�c�d>6OI܋!:ƴ�A�Zi]tc�D��i	 �N��\��؜�t��p�v�l"��觤��}����H����D�g��}Kf����M:Ç�J��k?~��0f"�G�H���'^c���~�"4��A3����/}3P�E�-��eL4�KT�!{�Cg�
�6��z���rSoK�'�n��0��F��:l�_��N�N�O!Ъ�u�0���q���#��W��q�TyFe/���\\?)~+1�ȸ��.�O_���q�]e�A�/;|�������S������F0kX��}m]@͡�K��cМqy7$�0�D�HT�!��T��:)�<�
�a{�ط��9U��xt�BR	�����ƻ���털��߂��(����6��$&�KT�*�4��:����ʼ;�;[�a�&�m^f�����6m�+���nR��r��])&/Q�8�� ߨyn��ӴT��aI� �]��7�����xRoG���\�\GK�M�a֢T䵿d� `�G�K\�����8�r}ː�����l�@��H�Ct��wq����Urk�u\䒔|̽��!yh0U}�+È��*'�2��ζY�m�{�\L����i�`�^�3d0���bt;�	|��r<���W��+_c�L[�}|���,���?�S���6r�zPO�B?U]��������k����=D�\�7�::*Ҙ�{�tYmx��b�ؽ���1����H$���e���^x�y���+�7�� ��g|��f�qe5�׶����!~�ntх}�,���Vg!�F�&�Q�2�}X%!P��e�WDr'QQ���8�D�:�t�J��My�Y��*3���a{�k	"_UPD�W��o��).��!^F�&8Z��1̒N��'m�(�ټ��8Kk5�q��N<�U��ac�O�ɶ#�"�T}c}�{H3>�h���n��o�A7�x����V����4��?_�9,5�>�ڕJ�z�+�9�i&�z�>I8d�D�<��NN�J�����M�+!1�p|��]̺�������T��G��>AXD暺V(�������G�(?�K6\b_���^fo�n-w���#ۤ������b$�'�v�D�g�65t"M��?�r]���RܫGP}-n��uX�v�;f��"~��p½�xM�o�o��Y�?�u^$���3�Tp��}�֔���i4�����?Ҍ�S.U~�t�R��t�����q��ă44���ȏ�&��E����`�Khc���.WӍ<W��ɼ���ڡn�'������j����d�#� G���^D:#}�/œ3�/69&�`~�z��81��:t���T"�޾3�.s[���,n�������ؿ�u�RU�UA[�-��͖�����U���q*��?��zMN�ִ�J�@�LA�Y�</�ãT$;K_믃H��
X҄܅�Y�!�-{�?�n���`
���Qr>��Z��(�  b�c�)F�I[^S���<�����l�S��>�#� ��� �Ӊ�sK���CҾ&���~;J�ՆОA}7���#�`NJvOY�IX}v�_=������i�p�j����}F��SK%0Y�<'��)գvǫ�����XUq�q�S ���،�>�$�*�&��3:q����]�S�]w��k"�,b���
J��Z���d��ߟ2�����H���9'��{�]"E�(�zs�TH�@w���oYeSs��5�\S�R�����eg�<Z#?3���*BlG��ܘ�q{`@F�@�)�aY�9H��.�r�S�^��Ի�L"���4�|�)����?i��	�f�C_�~@�N��p�tADDƲ��w�W�Sɮ�F��D۱
��%��ډ#��N�{i�ޟ�Գ�m�l��߀Z"�� �O�~�֢3��ۗ��o ���7"vW�[�5&`H�t|�-���V�Nu4��cS��^=�?f�`�q^�����1��2{^��Է���}u$p`��'M��q��?~.��[4��]b.�&�_���|,���yG���n�^������z	oB�f����,����xd�;S�W�?���c�^mY6�!�7&bZF�����L�O�"=���Y*�������U>�5�;��$�43}��q<�\���̋��
p���=��x�`�ůj5`9�^�B�b6���e�Gq�/��q�����] -�+��L�鼍�_(�}���T=۶�m�rS�.�I�"�=�f9�4R�v��*� d�F"o@_(�EG|����J�/�[�V ��{qq�����EQ�̍�o_!��#.V�����k��S$|�%�tG3�Id(�[����{݈푑�OO�[.�˞�[5�\��,�����lj�$�OP�ȼ��YcNO�#��;X	�~DtCS]b�"O� '<W��*%U���YY���Qec(�u������x�v� �/2��&���y��N<��W��h��_��Rӑ�.V�g|��9��ҽ��i�Am�<ͧ(v�N4U�(���Z��t��%V䂪G<��#g�of`i_�}�*�p�M���R�h�&�m���y�q����sƼ��Hp)���<l���8��ә����c>�B����?:�?���K�W����3c�q6�p(k���&]�K���Iy���.'�.����y��QtI1I��������ycٝv%��2V�WY�=�t�,I�_����O��=`VJ���
�)�Sj�uY��LK*#�E!�g;'-n�jxw��s�H��X����"}�����0_���'�u���@rX�r � yH#_J��&%����+�B�i��,�XQVX�,:5����w"_��_R����Pq>t41nO������4[,���������xE��������{���Yx�:亗/� g4�5�6�Q�ʀ�0���v�c$��nd�g�v-e3G�>D�=wP�^�/3ٚ����(� a5Չ��9ܓ1ʇ"O�	  ����j�ڎ-�	]��䦜����rK���[1�lx�I��v���(p*H��gG��=z�C�\5�.�Ζm�;v��W �Vw'��#����>`:? ��F�δ��H�Y��G�O��F,Q *�2� �1F+����������<���j̽,�C���9�g��6�p����r�����/��'?��d�l��=#%-��;��{X�h��`�N�g���["��4��j�Yfs���gw=s��ԗ��Pf���e�{b.��Cj5����3.x
4\O믻6B2�l��xAﳌ므�Q���S6��4OG8�^˕�l")��S8P��|=2d�꣌v�����g�Z�|�F���c�y]���g��_�FI�č(TSъ{ ���3�r�GG�B�����p�,� ��"�n�p!���o��nB��:;��-���Q"_�8d#K	�������K��wMm����!��O�O�Ɣ��¸�����"�M�E���t�Hj�R?L�ɕS�b_���z�y�e��_�Hd���8��{W`kT
��A��N������	��Ӎ���?�w�]i~��qͳ�W�]�k=�4Q��7����B����	��Sg�����io���� �r��.{ʬ�<����w"�/�+�ɰ{ص��g��hs�7�	�[��`,s�/Ψ�1��q�u\ƺ6�T)����>�e��FЬHd� ]���iU�L��\�Q��]5<A�3��b�JEnO���wJ�G+ΎkqёS?8]A�?�>�n���(6�Lx͍�]K1�]=��p`	�~W�Kz���'��c'o�5��ԅ�޵dM��p��50L'f^c��wn����G�s�8��t�F) H�9b&��|�f�5�H�e*V5�]��d�޼>r���޶d��c	8Lӄr��Vvn8�Έ�e�p�l	�mM��A�v�FBtσ�W%�=�e�I�T�����='���:6�P����8��(I[�XI��;n㙑Y(m�^�H��z������a�pi�Q��f>�N-��x|��J� �����L5ïη(V��=�1����e[�%��Sa��Q|��s��t���?�r�s�{�O6��;[�gr�߫�e�kի�ux��
4���"�1�R9���t5�����^1㠲�뢩*�\�CN[�P�X����"� AHy���j�&�����՗�Jh�tO
�q=ґ�S��U�
�z��.��[�^�T����l?Ѥ���h�Yhp-���2�@i�x.7��˩�� b���sg��Q�#X�k�M��i^+�Ȧ$��TF�����(ƽO#X���d^}!���g�����w?�i��>����&E�x�������	'rk�h\?Q��(aN{=�#��r�W�<�zG$����Sd���(����h�1 a�(-��D�*���Ҕ����ݭCA;)�Uj�^����t�9��o� �ܑ8h�EJ�)������]NKX�dhB����ݒ^�SbEba�!�kd��q����Q�����?(������!-Ռ�H�>��_�&��+w,˨�M�E欯>�{-}��D�3g���Ze6��f�㚲z�}��A4�ż�G`9RT��T�B
r��+����>�>��p,Tx�[�%���N��O+�������#�2������zPR�<�
�Ig��o��u��2k��UX���z�pJV�P�jJ�k��ʕGs*eh���&��'�}��4G��y@f���?�m@�5݄��V)�2J���\�.��-8=�)Lf�9�����om�8Dh�������λ�S`T��tw'��hG�M�QA!���=�aﳻG@\���0�/�3N*5|��U��.O)F���Ɋ-t�,�o����ќa�2}aJ�*��[T;;72�E��!�b,�9t�$�����!��� �k����V��ki�⮭���KD�����e���ۀ�3�3�Xg�+&���Z���n�:/~ 1Ϡ�1�:�*��F4ol�P��h��g��P]��(M�/���{�ۡR|ٹ�![˙z�r#-�����k�}�&�o#LZ=��_6�[�	�iD +�-#G��\���$�K8a��%;�$H ���~+��j��K����ܮؤ�F~�Á�Em�s^�^`�h��`���%��OC؞��EE�x?�/͍.]�s�(Z0�r�;�[������@�'V���\V�g�g.���e]k�,�0E
6˞�o��s�������N�;hD$-�)l�F R��qϝ���Ċ��pFHŶ�/I�֕Ы�Q�P�:��	#8�6Ɋ���:��?�9�٣�-(�>��ݙ�F)vR)�.�v-�e��Xӹ�B�)�K�Ȗ�q�ٌ}�kM���.+s��毐HsI��3�26��H$�G�� _.��d_���v屔/�]������s�'����[ƛv�]f��Y�|��s��Ɖܑ�I��|�1k��ޑ��If�TZ�4L�����B�ۓ�w���	�U��}SƳ�m9x�1�����BB���o�5'c@�H�����)��f6�0�����Ú�OX�t�Ư�^��������d�tc�ao�,?P�G�^p�`BF��v��ͧ�g��wd3��j;:�i6�[��$�J$,�xo�fi{E��E ��P�`�1ɳ��K�1-Xh7?���Y(�^Y�Qi$,�͋##O��L�G2�q�E�Tu��gJ��\����Y���y��%(`Z�[#\7��b�$H��Ym�������]��~�U���I��~fh�A�F�,��T$z���+�a�c@��WQ�&\m�m3���s�
Ѳ��Tny6���x�z��=��%6�d�w��M<�Y��O��Q=�$G�b*��A4�kqċ��f�,�]��y�I�W:YsBG%ZY4U=>	Q�O�R��ή���B) Fr�1�=X�Hqv��q�p��El����7����H�m�����������i�N>�C���O�`0]|�E�]v�7L��39�]W8ίK�qL� ������<�B! �lE�j4D-��%���r�oX4dQ���@`��m��g���j��u
c����.���.�q ��$'�9:�ã�@�2d1�'/�T�y��v-8�G�[�q[�6?�~�}t�iL̶���i���<�qp�a,�xT�-I���O#�Î��/�9���?U��}A�����9ql6�x#hV�;r���X��b~!��h�C���>��ๆ[�[�P�|;p�Z21^���O���#
W��> �Fء����@W�>�낆����6�o��̪&H>����(4��	��I ^��[v~%�ĥ��v#��ٶ���$��2)�t(�6���e�P��6�$PG\;��N��:
��2NA�b/��:�(�H�aܤ4	C��ͻ��g��N�B��H8G5-�ǯns�����f��ҁ[Jf�b��0u�;�5}��Us�^��$��m�^Ѐ^5�4گ/�uyL����ff3k���ꡅ�Mۖ��L>JC���B
q�٫Ԇ���1�D\��z�H�\h����I���ܮ�����\}���+jr��V��X�/я�Ű3�>�}Qr���8vb���]/wiS���ĭP���� ���7���
KRH˜�K3�i�Jl�|#/+]|�D����5ɜ^���hO4J=��DT��Ȟal�#YD[~Ґ���"yw�hw`�դ6��|�V�Ǳ'��8�/����1�P�u�ȉ�)K;�-|2D���8��`�l�7���7uB=zJXqo��U�FեxL�J���c�b���F� %�/g�_Tᤖ9O��F�t!�hrߢ�@Q�h��oȢB �c��%�-���=���S�i�:���B�TH�Wv�Į���jI��C#�}E����J��V4�A}�Y�!���K3m�J�'�4LB��ct(5�|
��b���9Տjb�bU��!He���xzh�SO���w��vm\���O���n�j���%�Ze�`��`�^����ӀZ�+�>'��7<��=f�?��K���8-�Sq�t{���h�QV����W�r6d���G���/��ɹ��}@��bK�+��b[T�Eq;���0�2Vc���*CN�
��?��Y���T��8zf�k��K�	<	���bt��������:	��z>d�+�g�]�=����ç^jr��5��k��'��E(�>���+2
�8Ѫ�݃w���y(^e�H��"+m�cc��)��zWc8�b�Y�\>r�"���U$P��j��ͻ`hؑd^?E�ē�X#��R�~�T[�g�Y$�ң�x���یPӟ��c0�0�2��RK�m'���V=(����g	<�K��j���O�/�����le��Rl��6G�:J�}�F�[,*�k�~mW�LU@^���˸�b�إc��� ɒM�����b_�9���D�>o��1i�U?p�ʒ,�"W�:�H��j�忇&o��eݎ��<�A�\�1N_b�uaS#9�W���a&�8��.�?1WaZ��K�T��n1JQ�`����������?�(qiö;�2N�2k{jAb��u�a=�C������ۆ��}��z;��*�<��4@����}��T���`��v��|c=�2U!�P�l��Ա�S��у<sgPﱍ��ⱨ���!V�/��GL?�m1�����v�!I�o�� G.ϡ��I���J��^��%�̓>����w�_�ޡDMv"�.�h�.$ v���c�!	)?��87��b�e#�r�	��oǺ�?��k�|��F3��o�v���>�!�,Y��
���m���*C�բ(�3�O�/�Itan}�MY������!��i�;��,@<�X��r�t�\y��vNf?:�s�:m����x"{�<b���t)���0�D�1�Y ���@\�BjS.���/a�%T�dU����GII�6aE��XTbǇ�=7�!_���Ф��*t:���������iQ3��%k!�D/�BWS��A=����Usb�%0��7�v�.g�}S�6Ŏw�^pC�$�q��)B_�'r���Ns����d�]V�ʏ"x:� ]rh K���-���yV����3A��5���.
:=T:wO��Y�`�v���������g�e˔�P����a�R،��е8B����p2�pɐ��\Z��XPr�L�01�~o��^�`Rэ�a�~PЛeU�Q�L�
���K��t[���RR�H��_��oI��������,HxW�ľ�L��zY'<1�tV�.���ܯ/?Eb�ň�;F�/c|&SOP6���#^�C;\�Ģ�g�E�����l,uBv��R��]����=䷎7���͕{
K��x�� e֜o�>NKqQ� �ЬBdA�m�,�0�6����a�<k��IW6�?��ŋL�z���ʈ�A���H���F��Ǹ��q�ĵ�EH�?��;�ߣ껢�@�1��K0$s��Ӎ���S��E�N\�����]Kzy���fۈm�Ǟ�c��Yt�g�������k���-�`�4)�NYaE_N2T�t���/�˿��������^�5���>WϮ�C_����#J|��J_'��|"��O���칾V�f�f�'Hf�?~c�����d��J���)O����z���}�*�U� D����/��]����,�fe�kt�6�|�N�����J�;� 1��I˪s���.�O�d~57U�������N��kN/Jt���a)8�;8Ya�\�t'I�9s%D�0��W�h�|�ѿ�{oB��Y�~N������v��S�g?u�/8�붍d��:�B�[U�M���~��0ʡ8�
9���xh��$����K�0����y����	�է��Ν�I�7���%�S��w�.�pM�0�[�PM܅r9�[����j��߯��(��@�qZ�r�٤������m������8�*u��9d~�1Gn���Fa�^��5��f�bK�۞��-�_��6���0�Z�uf��-�����iM(QJ��� hY_S���1L�<��z\�K���{noh���F��^�5����OG���Ŕs��{�򘛛Sm[�� �E�dc��ҝL�F��A8߱P��owp�~��!�����S��� �E% 
oD;���+�eO�"�~q�a���f�����;Tw��A���s�*��=`0D�ҽ|k����u�XI-�:�O�0ή�Gԡ��f����@�t&G'�f��f2%��&�������JZ�A�m�L��s�	�
��m�N!<��HZ��e�5i���rX,�x���p��������;"�%@tO5�al��+�G)�P���h�I��<3����L��4�aNUF�6�S� C 4�7�-Lb���"L;}�C����3r�7tS�dt�I4��8�z�^��7n0 \e�ऽ�L���.cq��?�����J�s�>s�k�T�ɾ/� �al�����M.�-��X��;�r̓3{��c,HL��2�C6\���w�ć��S�=���4�ZEUA�4Ο'IR�T�D���}��P^6�𦎄��W�t�xH �X�.��<�85�:�h1S9>}�"���/���P��?NNm�ƶ�cJ����K��0�N ���~jKg(���s �ٹ\�JQ����T�[o��R��x��(�#F�Iq�?�+�o<���%���7���G\���Ĳ�Z}�E(~�?`�5"��\Yg[bXB [�OM��	\�2��� upZ�ŕ5�yIT<ڸ�r5!���q<jZD+�Z*0����Elu	�du�����n�M�+�K��d�^�՞��*f�G�A`�Fb��er�jW(�C��<��0G�+~ˠ�K�n�0zށ1�������y��O���,(Q|���w�4Ϡ^S^��ߴ��u�Dķ�\&[����>��i8�b�kX�9��r���4u����C������������h@�S�z"˼��8��};��Qw�� �C�0#.���IO�\\C`}.Y��K9���Q��D��&�JZtf�C�����#$�i���h�X7�5
�D�p�V>�
B�\��Q������2�^���`-�h �{���k�x�s�Ϻ)�t�����������z�:,���FN��wI�3�G�^Y�֮pq�J<��`�� U(�1�YW0�P|�{�ЊV��Ͼ�Q>��VF�S��t*�Ʃ8S&�s��{�:�;.tu�#�X�l{�@j�!�g�s��0��M�>��[T��8���s���{�'����71쫐0x����|��7�Ft������
2�e|��ߖ�\�st��4��]�g)I�gED�LO�E�wr�I;lb~��Z�{w\��M�@��XE�GJI+!���KoT�nf���7T�$�T_��r0ǀ��+����"��)����c�)�a~��DC}o�	��0���X(�-�1|�a��͹["K�Bu�P��׭TD�p��ϱEU�����vHč��B��E�����"�x��5B�(��n��/��4D�!}�p����1y*�[<K`�Bo5��C]y����};. �����H/�6r$�Q��?!�����d�n wu���y�8m�����o�<rHp����J�;�����k�0��`�N/�ݺID�h�i>](�����N(��Y?��T�:���v����<��wt�v�N�ԃ�CzUY/0.���tmW��$��"u�ɹ��鬏��R��l�0�f`��$U1EF����kĹ��M6�5�\�ο����'1�'b4���$#��;��}���7�i� �	��lE��v�"El��M8r��Z�F]KQ���ٰ�AP�6��f�::~2�=#,+/ӎ���m�(J}A��M�i����Ӛ��u�$<���z�R�CӅv�����G���3��P��(�p�\{����P�)T�;���ptq��+(�|�x[4�Q��N�P����n��2�:.�_�'�=2l�o�d�k��q��`s���Pz��'Y�>U�<x
��~���qp<�w�x�~*c��tTw�Z��Ͱ�-�Ϩ4ێy���I��a>���GL���N\���E"��|�#���7�ʡ/�W�5j.8#s4����1�;֫ݎ�Uʲy_���O�7 ��D%,�-:N�1�#��ޫa�X�@�KB�&n89�IJi�k@�RL�,�o����^�����M��߆^\�
�;��*m�9�ٞ�HO�݅0Z<���(}��m4�&,N.0��V�C\�d�[�r��6q9O�N�)�I������a���)l�Es4 ��O�?���<E	�d`�p0���%��̪�1J��$̤���x��ӷ��#^	^��j��R�w5�����T��8Rt,!���uw����SNr�bө��I�zx���s]�����
����#��`U2��U�J�ȞnU兔}��wL$�5G�����v��
����M�G���)�R_ꩀV��HU, J~�e�3����bgp��G^�D�x��$��]r���V7+�@�1'�/;�}��qdcHĨ��؅55��Yٞu�Z�J�ɬfȃ������(q�{ ���P����.p�I�T�euc��D�ev?e������7��������Ž��P÷	�������f~kRD���+gE�#u�Y-]�/�.T��Y��K9�P߭ZZ*�=�=�q*��dP��T��Q�S٤E�Yr�y��P�L�LƖ��0~2̙�8ԣ�lb+�cm
#�8��H�Ü9�\>�X�8�n/IE	+&.��=��[ܵEV�v[l�ǐם�&몀�z�g,'�O+�M���H4跽JA�}��~���5-M��~�XG�#0+[�8�=�d%��Bd-qؐw0O��i�g�?h��g��R_�%>�r4�l��c~�_��5M�׊�w�;2,=�b�?�-C���wT�3~1�l#�=����8�J��T@�M��%�d
T�Ԅ��o�J������4����/S?�ӣb��M>�.��n��b��2����o���[>�{ ?���U/�-�R��&{]����:c=�����MOʐ��b�	h��n�΃U��UI���cC�n�o��q��9������бP1��@����2΍3��,�c^/y�6le�Q9��Us֊v�$<��5���̯:!Ko�UZV9H�x���U��,�a�\�O��5{���x �Lu�A���J�s��� '���O�q�^�6M�W_|R<Ifx|Pj��B�ü#�!��6F^7��fN�:���������hUTW����<ٺbbM6z� i4�Sv��I�6mj�3��J��u:����*��;�������Ѻ��\�)5`�T�i�j������s�l���Б*�W���edjF���f׆�%(�0`=���rY:���}n�Zj�뗾q�_�J�^�8�~���L�A�@4�#4r\�Ե�q�S��K�����V�Q�L�c�\=X����j|���H_��E� �r�x�� ;޽�-6�&!�Nl�]rG5� �	���X��9��si"t��OE�Lm��@(lr�}�ۓ*�w�������w���{h�@�y]�K���-��j���P?���_�C��į�?��m��J��*��o��T������G��=?���m��0�	C7�IX3���rd%\�Re{J:d�ڽM�|�c�7��\j�=ΙBx(��$�
���`�8͘_����ɘ��\�%��z���+�|)z[��]]�0ڃ}�I�2�)�(�g���_���v�b,��18tL� ;ݖP<,���LdmG:~il���P���r�Kd��M �68��Y�n�e�kT�����Bu	27����U���a\\%���/�H�������t�-�'����z=O?���+����̧��PD���PH��=����
hi�@"A(k��L�Ly��xW�o�m�$p�����Ȓ�4��F�K�׬ퟎCg�G-�u�;h�K��P��q�Yh?�(��R~OW;�gWBh>*���_K,����΋Z$%�q�>,���傩ϯ*k������ʬ�U�;��j$�Bn��u\z��͇�$IŢR� Q]���a|d��Y2-���iuk"1yk#�Q0�&��>�leK؀�q���9Ժ��T���pi�j�N�痾�c5���$r�J�,���픮]��=3���Lz�V�c�(Z��t��2K]X�|(�Tz|=�_����q��������q�8��t�����V��Uu�Ukq�>�� �"P��X��d�r��oǕ���ێn��X
bc�û����v�+Q���<��"��(�:�6o��A�M�Q�8ʆ������	�\t���v���4�vW6���/�sui���i�ϣ{�qSb��Yϕ���E��gb��#�ɤ�(�h"|ĬMW���2���%�~e���T3��6iektV\���>�j*�3'] HƉ%�������)2�.�@�#K��`u�*����C�l�h'^���W�(!)Kg��O�Ц�ѓ���
���9�D���	K�6靟�t��Va����(x�ߌZ�Fkh`������\�Kx
��ߡ(�B�F@�G��NZ=j�]*�`�>�k���!�O}�$� c�{\���ߐa��9����G<o���p_w���������*R�;J�d����`��P�	-I�9��>�e�n�	�n�wH�`'���[f�1��x4�O�F�588͝J��~ߋ�rW(0}Z��3vΊѤ�sc���˲���;T�7�``�G�?n��5�G*OQ�:�=��u�}b^kvvKv�2ڌe?l�L�2�YZ-��#�l:��~v��V��b+�Pq��}Y�����Vz��j�t��9n�:�\_�0g���e	����![��ڻ��T��_{'��R�z9��j��ޤ�A��w�d46������{�_�Wv�<��.ޙ�ٵ �Q9��vs铠 �p�	�72�nvI�?lc&�g�ۭC����	\Ʊ��HׁR���6�;::�i聤O-��s6S`�i��X�hS2T;�|�R�ڶRWV_�2�.:�pG�t�;�I�@�1�I[7<�J�Yu������6��j������@�8����R�Ռ���̖��K� 0�^�nP��� �G�R������7��;I8wY ��f2F�x�@����N�B�]�Ҹ��y�Ţn��M�J�� n�QQ����ڠa���s9������c"+J�����:��h��/ԗN�o���$��� XK"��O3���o7�z'��@�m�ո�w�{���Ȉ��Ü����M�변g^�	.�Pj���ŮT�߮r5w�Y�?��s��)�>1���H�l�{^����1/�mq��>��^�g�F`��)2�Tj>�r������!�l�h*��J��ɕ��@��a�xZ����nU�>܎�N䂎���Sנ(m֪����c�g�q[���G��=��v���:�%��8v���T�BM�pw�vG�j>���{�Z/,����%�t T��#J�OT�Z?q2��n���E�(ÆE#�}��e����EG�>��]���@���|yVu���7??�E����rT������l��6	��$�I""v���!L������Y��+Z�f��6��0()�̭�,�g��z+|��s]�E��l~6S'��X ��#�ێ���$X.:�g���hO��\����sF1ာ"�s?��� D:�U�1��{�����wĶ?�\�nK��2�Ę{�$��x!�D>R/Dܜ�\��$n��ًSW^�H�K��{Gx���}��1/��K70r08������c:1<�}�� u�9�9<�=�>j�AO����z�W2pm-�]���12��~p%c��vޗ��1H���6y��J��9�˝C�D;I���)��z���<�_��mW����l�Z�=�(����M�G�)���_�0Q#����E�V��E��cb ~�#񉌥�c6р��2J�R��x�������@�F�����9������U����+��@��0#f�����b���qH"��y�N��{7믎!���H]�miQ,T�.�{v�>b�5���IL&�i�� �>�Aw(J��osQ<�%�	�� e!����v���Hp�^� ��lK �fl�;Ü�����7}���}O�Z���dr�9�E�S�lސ��2WO�]�rx�
�R<᠃�'�%�Ѳ^(H���I�)M���U��:04��)1��p�Xc�X��iȸ�Y�����$����o9,�V5��xZ��m��L7.X�c�D(T�B�	cC9�����ȴ��M1���T���qm"�F��H����У1����
]�z�{`{�,Þt�g�ѭ��Xz}'�Z�����卍o��� ]�r'&���  �sӈ3��B��[uuGl~JH�lt��ّ��@�Q��oƭ���\�����[i�ZRr�9볉 
N%.���&u!Ʒ�x��^(,�ب?�JC�A�B��}���3e���x0@�T�wP�� �-�9�o����ಘ��N*��T�qBDEI�ޖg^��P`�u�/�Zg48r��� ONj����g���N�A4�c��y��skv)1Z ������-	��[8��e-Z³d5ak�Gg��K�����s&��JH�ئ-we�$��.CwV1���ۥ೤.�K"O�Q���۸'U	�A�22=�C0�ϩ�- 7��l�N�j�Yx�%zף9$�=����K8"v��㐩��[�%���8
ƙ��|�j+}��f�I�gJ��ZJ/2�8�Ќf�Lf��k��q/o���ui&��Z���`�s��'H��j[��*�����6�xY����cSOQ�F�j���y�)��N��9��r���I�8�*�������	�p�l��e�@��1[{ LX	��6^�Y![#���RO^s��8��|�j�����<
�HZ'a�`������v�³7#/Z?ȵ�m�ؗ\VJ8����t,]��z��O>�O��W��/���P�_������p���'��?����Mx}�OX����I�Vܻ�W*Q��[;�������U@7����깮���^�=>2�<���pTb���	%����(S;�p����J��2�ZGb~*�F/�3w(��E	ZM��j�����!����ܾ���� JVG�kx �`sLĿ��p�
���kr������a]�d������M��h$�=���wc��p1�2�S�"��2vo�[=d��o(,�����j�?�_cmNhk�u�i�$�~�7������f�C
'�ߠ~��3bRܼY�z��0�����S	�O�t����S?��+���n�i�#�Pʤ?Y.}_���ci◘=z��h��]M��V�Qy���z)��T.#������(�ĹIU���� KS�G-�G|�4&�X��7�:'0�۷G[�D��EAzd��C�C��U�eFg�'�J��4"��n�V�!����(��N��y�o��%�@ٻ<ܔ@��;��`�#37�G�{J�ގl����_��#.�p�nMǰ����^R��n0wQ�&��o$���/�:�L�Q��d��hu9	��Z[�/��G��iu�IB0��X�"�mڌ%w�BeI
X�pS{W��?OQ�!��o�.J/�}�_dm@[ߨ�-҅t�;؏)SO���%QU�-_���φխ��
��$�;f�|�Ӟ���r��/�ǠX��}h.cs$�dK�+*_v&�;��G(bX�<t�rE6���xFW�{�P've+]�(�W�9�q1�3H��t)rAo����g�qiĞ�(�<t�X�&+�8�bPs��t��j�=�ål	��|��;���/F��Gʡ���uu��%��-M��>7���8$���)����F-f	�n���ٕ��`%Kn*�#���o�-p	�5̌ķuk���t.�:�IG9|d�b�g�! ¶̚ �AL hj��sc�w
��������b�,�Q�9|7;h��'�����VF��@��E�O�x䖼��t�K@T-?�/����^���X���C1��.�V��0J9��0�
�w�x�����MS��ʦuSb�׾^t�N�ux��I��p"ܹ���FK*拏˖�6�ԭ>��H�2��4���>d�#l��T��~��;n�Y8�	#A�z���%����Uk+VM�o-����*��Qs�z��+�F�Qi2s�S�q����Ԫ)�Rk�u.2@!m|�Eԭ"�`�nߕ[��۶j���ũ���+���������aP"K}��)�-�3�Ӟ�#��(3G>�Z_����k(��a���V�	���B�F�]:O:��>`e`Nj����,c0���~��I���D�`�I���Du����6�=��y`@)}�^��z<���r4�
g4�j��k���Q�)����Y�yk��Y�qr���Dݦ�����<�p�\Nۡ(h�4g�Ƙ.N��tQ�U�
�DD���,�TO\A� �{A�w����s M�I��H@�A�w���H���{#gYO ]����K=�S��"ț���9�1�H00�V�=��:�!�ɴ�����@xǶ۷��A�%t�T�N�'t�p�p:�p���6��/l�̵����ho�50� ����ޠ3����Á7���+戻{�[��#庅ԁs�t�6LA/>���,�(wk�Y��c\��j�w%�Ca�R�v������xV�7b�{_���$����>S�ލ2�-@s���*�;���>U-��e���Z�8�Ժ=V<T�5��2��n�%�>�{UF"�� o�R$���P������Һ����4�d�U���{^�z���� ���X�Y���+ܜ��wwWsQ���%��F�ocb������`"],�Y��}�E*ɴv,�Bw�9@�$p��-�����/�!u�0��ɖZv(p�Z
C�����H��PЙ�4��V��� ��q��AF�H��E҆�����0��Z.�X��Y����o��>tB��rB`�ΊG���]d*Z4���;`֖Y0FF�C�R����v�Ӄ�/��uU�3{�X�'�;�@��99u��|��Fu�qoq�<.�_)��a��z�WT�j2Կ3��z��ꎲ�EhN�J5AA���2�"52�hǤ��C݌�17�@��O��R����Q7ؽ|���`�Z��$��ƥ(~I��B�M���2K��Α��=[\]ȃi��P.��7q�n�;KȚIr�!'�5�#��._��5���v����{��;�-�*I���X �T =���c'v<[%`�d֩1H���'JG��^d��Y�I�8�0\�!�-�R���$S�<�:�y�gCܻ/��F��|i*tU�}>oA���,�o���z[�q�E���W���)q5�8g����-��-����H�8�<�G��sV<|� ��]�񟋇(hg���(5 :C�d���p�"�Bm@��(�5�Y����"\zʺ�P�^�D&��'���
O�+ :e%��8	�~_��C� �%F�h�y�B�Kf���e�qKǅ�W�ޝ����d�L�������x�G���7콌"���\�15��ѯ�3���R���������.��V��> ���c�C+ո���r��H���E.�"��T���.�u��ɩ=X2tD\����gtmP��1^d���m;R��ϣ��FOF�֪�nY_նO����	3UH���8c	:���^{�l'-�3@|��^�Ժs� ���|������&��ݬ��P���w��J�_�Z��n�H#�Y8��
�<�`�g��F�~�a h��_p	��D�*.'o���_d��yM�&7�朿h�=O�{����CD@�E3��З��>���j8�)!i&L/�Nt_0��q�gM���H��X"9�ҡ%��σ��0�Is7�p*u1mQ�I�F�xYQ�D�ւ	�}��Q�%��Lb�>����u�����:�����$6e"X��n6�@�.�{�.���$g_	�L�DM~�"��w���Ss����S&VH}��FHr������xo�z�MϾF7t��7q�qo�Ə-�#X�ƥ9P�4�ދ�vd��`�6<�2���GE.͟+^�lbx�p�9pA�57fV�/h����N�)vst�s��|R���=K�G>K(}��KW�	�m�lѹꋑ��������e�����/����c�t3q'H��y�r{���,�~��e�38�����C�'Cq�8#R�.ʬ� ����Ә8��С�0Z^�:ub�Z��7�gH����6�ز����,b�Y���X�h��w���4?+�;s��t�J� /W��fK�(��Mξ��D9��ˡ���-N��X���(�	��16�*�E�"u�1R=�a[�5�'���5�h 6BCF��!V%�S�y $�(�!�W�ib�1bZ��;��I��l�.����C��@,�]i�F����5�q�+B��-�x^1�����ި�e� ���X�P���Dw宀��.�D`���A�C�dd %5�~H\��Rꪊ�,���-%Bd����+��k��=���NKG�`s���s�
�S8�,�k{*�9�3����;�b�[�>���g�9:�#��qeD-v�_�|p�ҳ5�Xi��7b�w�} ���s��	�S�79��@�=�7�z0!P߄7���ȐR�S�N�B�8�u_��h!�F��"e�oɛMj��j������En�M�����l� 1�����sA��T��_392 Ϛ�=h��/�W��p��Q�Emxy���
�2�"��{Z�g,�0�%gm�q�u���ʬ���c�^�MR��J�ی̢))��\%�yɃ2O�-S?z�o�2ۃ*���E��q8Upߣ�~��p�&�Ea�ȹ�h��T��B�q��/�����������C�^��� �0G����r�2L����8X��,�$����j���K�����g�/�y'KGd4h�).Ar�@Z��M[�p��e��n���k�Y�����{�ەkj'T#`.?���}�LqO�^��m�Q�ƙ#lP� Y'W�#���A��g��q�O�p��F�E`���t3��l�y���أ/�B���a�Ҕ�.�������k�?[�)�d��O��	�Q �[
�q�j�6���н��)vJV��c"{��eY��ȫҏӻ�	�}}
0L���WjX�R!��m)Va��rV%ě��<�L6����(��Z�v�����"=gz�4�8g]ݼ��r��G�7dճFT����WB%��-8�j-h��+�0@-�*��<oL�f�����,O��7C0�1��naS��}���혓�u4<8��EKēAk�@�ʚX$9��x\a�Z��
C�@dۨ犊�D�%s��Y�a3r%u��� �d��P�%��D�]�]��Mu6U�5u���`���A�
��=���c��s�+r���9o���ͩ�J�X]E���h99����dBx
���FX�x��@,%�vck� u�����1t&#��d�5�Ѩ,� �[��v�}�%�`��5O^��U�k3(EmJosؔdh�:3d`}İ������+�AW�7%��*/��\�`���A�xQ�J��-�a�*�h�{��Vez+�z�wv��)��K�K�#�YE��1~���ji#��;�%ۣ\Ѽp��1^���z�Wa��P���R �U�%�2rE��|�N:��:�2����"y�W~�Dm�
��;
]L1Hѹ�A��{�{�3`I�)���@b���k�����c�e�R�Nj�R1-6�&$���'�/�3�1�8)���엀>������Re�����sǃkX�H��R,�]� �W��
w[c^MT��3� @�G�;?�2yoXc#�[��@N�5��R2�����;F�؎�fWIdPM�>0��{��qk��h���T
L
��@�������[q�*�@_������cR���tEjBh��>c재��'˭ow��;\�n i��������3q�S'�݁�9X��}v�r��1���	�=z����ۡYgS��
�\η����wr�	� mWX�`�Yԩ[�|pxiܲ'{'�%̎�>�[@PIkt��̲l��k�;�#��J��ah�{��ג��OSq���2xbg���J�u��<Zr�ц����hʛ���aX�=�<T^ac+.�Qh�%�1�a�� 1�!5� `m6O���ɫ��z���M;�����=��!3Ȣ���.��BWN�1��n;���T�Q�Q�jW�RO �}���:⊻�������~��p�!�Ȫ=��S6�X�n@^ǉ��UVd�b����X3������7�@�T�L�,,KJ���1�4Q��!���0}Bf_���q���a�ބ�'��;5-<k�w���B������0Of�3b��*����!aU
R�Z�9m��v��s���ER��R�yY�������T
L$�x!����0�1EV֫O#v6��٭��T�"�"*!�k��GR�Z X�s�����&��}�ؤN�5�v�Vj/�}b����{��YDƠ'� ��7���hJ�T���XO9���
�*� ��iۈ^#ܐ�逭�m�X3q_A�Q �E�!��W��@�bkx]�q���AI���k1�.k[i{vݢ&��>M��7�Q�z�'�~q����^G�iRҗ~9+r�$��)O�@G�$�����o�n� ����d��m��; �/�/5T3,d��ؖX)�d'˪��ܸ�?�`!�C��=�[��&x~;&
�>M5Xv���F��}	؈I2e"�d�����KD�x��;b?�'x�~jR�� �
C��@�(�ú�o7[��L�@�}�Z��[�W���hg��\c%�W� �B�f�L'FuF�M�{}M�5�9���&�W�=3)6�QI�nd?����u̙����m��O��a		�V��u��CS����T�T�?�4��:�R٘�]3� ]��H�fW=<E���Ӯ�a</0�ѳ�����b�s�v����3!���L�i�x5�*l�s\g회���&�y:��׈�9�N��vzb�DsIJW*T�#��.a�،��p����g7��;���W���G[��]5/g4�%���\���+��d�t���*��M���켲?���"nYT!��#��x5_����h<�Z��&Mi�_~u������S��̀�ɧZ����_,�n��85���<���ҝ��y�n��6 _�`QG��죸�"U����C{������-�8����K~
�v�&T��o,U�gE�e:ud��p҄�$-b��_V{�����(>�y*��:�1T��:,��lv��'R��G��u_d����?����"ǁ�CI���R�����3�j��Tl��ӂ��M���$u��C��۝�1ӝ:����H ��%B���v@���uU�e�>|��ѵD����<��:��M���u(dyv�b܌�;d0�ڜ^�����q�6	���4��.�T��ۥ��+�����4�u�9�4_����q�=	��]��u��퇐l֫�?�D��/�x�^A�7%�b��?=;X$^=�_ ���O:g�-S��$Lr eZ]2�ӛDA�g:Jk�@i�F`�X���e�伊I`��7��M��M�Ӓ��K)��𒢪�2k��C�ߥ�e�� �Ʃ-��(���x�O���u���B�F K��(������i��ı�a���*�՘XTQ7��#D��.4-��N��v��W(qmH2=�`�<�<��IO~�tLNR�s(�EY�M���Sz"t%��i2�*΁���T�I&�e"��D�p��9�@�r &¯�k���G��
*�-X�=���9�ǒV�38k�����LN{�Uت�HJC���|�p�����cmN[�p�>�zD�!�]���<b'�f��gJ4^���Fac��E����7��D�yN�I"d�X=(�W%�Հ��þ��bѬK_h���R����μ�_��0�� �)�v����VU�ʉ�(�_�y����)� �/��:/��:��Q�>��+j�,c��U5��Z�S�3��^m[^y c�&��#M��d��T���r755�� IGM��.�2��P4Ey�.K��Z���ʘ	W�]��$�x��3��+p���)��6�2ɦ@/*i?E��PG�PE��b�3�`��)x��v�;�uW>#g�{]�R�S� �(ւV;	]D������Z���}.-���`T�,��bD�.�U\�<�0�V����-;��2\/�l!����Q:̚����
��\���]�Uy:��ųG\��\Q������/*� ��c�6��@��yK2d�� �[B��ޘOLν�j/�jR���؅���ǧί�[m
A!Mɭ@z����Ƙ>/F!1`{(xh+���9��Аx�d���5����1WԐ�+1K�тp���.��P�ai�Jd��*��̘�~��2Ozǣ�+	�e'��P�f<�A�(Bfi��	��jgy�/�u|g�.��h����v��! �����A��4����j+.�H]Ϡ$\��n7W���:U�wkl#��Q[E�� np&�x���bH?�rc�_��.n��Ȋ��qn�c����z{���]������)���ld�1ucYF��?s~�]�v�G=T��)\��mK�����yr�I��z��?��K
�F61����}|�C��n�*��~�2�ޓ�F	&�=ҡb�A�����ُ{8[�vC����b�����w �����;:��;��A -^"����y	;��Q�������V ;�Ej�?|�|��#n׹xX��ƸM"�-�s���kq�p~���>t��y� _�����I2�.���l��z�-��b�Wl�6y�^��2+����?+  ��_�������hL�zsj�B\�B}:ߴ�q)�co�{�$��R�N��g��|u�n��N��g�R<rM��^�������e.�E|�ME�^TJ�&�HԳ&o�ҳ�-J����s��V�Q���Đв��d���ۏ�`�p������g5D���^C)�+��=��8i»�qh�i�̮F\XY4�޻���Ea�q��}���Ik0�s4�����߽y�S���ծ��ŧ�+#\��Y���zOS�C�eG�#�����nV� �����!E^5 ��Z�Է`3T}.�G=#3@;I.Ԝc�^���#�pLK�.P���ұ5��Q!�7[.[�;
����򤆍���mnҪ0�,i���� �j.ͷ\ã��T���ZbZq�����K�@N�����rX�s�����"աa�Ox
d���Fs��%��R+�o�wFZ��f��� �W��xh�ڰ�����ۅ+sޥ��jh��>s��g�xdO3��I��ʊ_uG1�h��	C��'� ��k*|:�r`},��������2f9R���,廀�[l��IX��&b�I��>W������s�ޙF�H����9�D�O4�ak��������<7�[��$N� �b�Eԣ+���2��h�S[p��ǭ�?2VuZ�Z��a��@�����D4u{��/�Q�ɁV���0�z�9�e�]��>���$�Q� �հz
𽄑d!�r]��.����R�E��:cRƪ'����8=�T�U�_6����c�6J|�3�gϖ��{}ps�S�ŕ�Ѣծ*9�g�������Z��k�3b�4��>�ǝ���ED�dj�R|X���N>%�!�� \�`/�((�өz4���G���Q�	���mN�I}9hB�AG�rT֐Z+=^�'��\�r���W��÷�PqDU>)(fw�c����&�2)�/��&���!n1E�-���Ѕ��jϛfch-P�V��uzZ��ձ�~�4��%����2s׀m]��e�[3ѨVh�ۚM�"��~�É��N�+���
���p��6�0QZ���;�xz_�\�n�Ȇ<��������b�٣B�"���)MƆ�Ǭ�����6�ׅFϯ��Q����R�{��8hY:Nf������ON�����P�Â���s�2�ƣ��eHYc����پ�H�SI�ϴ'��C��Q�T�$&VH��Ɵ������m1d���u����F�X�M�P5z��V�T!8-�c�Z���!�ƞ���;�𷥴�a�g��x/���4��n�[�-�E�֡6
l?��Qʕ���u������i�AG�z=��]�Bw�kv��l���;�N�0��I���U��������M{�����<�Hͨ*��:z�1�]���4�Z�:�y��&G�eg��Lo?���?TH!H��~b2P����oW�2�� ����l��<��������\!�k��2�@N�^)ū��T,U�n4��՗��,2SJ����c�e��� x�l���TO�g��F����'���%���{)w͕��[��������!�`�|�4�eٮ�qǭ[��x2̐�;�Ze�O�{���a�E� �(V��ep�7����(�g8���hN�)ِ1p&�Δ�U��jRTtib�{��~�� �ǜ\!�^d�l�]��7�&=���X�j��]E|�ud:٩��Y��ي�����W��!��+��=��\H总���CB���:�~�����|��̂��cm��n��p��6��K�?l��8b[���.;��Z���SL�jȥkڜݖr;%�6xn�O�#��(L@{�&�wz�C�4ԅ���}�RK^U:�^�ȁt (��2��؈��ӄ��'�����)w��?�.75@.NN"�k��X��D�#-r4�UJa.a!!]�]�{����\�����T�3���ͳYx���u��TF���C��^i�*0ApR����T��B�ˇTU��յ���#�y�Q-��)�j����m�L`�"F�����[ן��d�̝�������bF�������Z�vTSn�ws�v���J�_��vNj~|*�P[�%u7"��D�,Ū���z�6�B��(8˭{yΊ����7
�gg��z-|�z_bm
3?�x���"�*�������.����5���0`�+��8U�5^�'��9x~�+��ɬ^��5g���'�5KLM:S /fl�`�/!w��/���wu�gSEK������d̔�I�w��5�r���.N�O�2�'�x�8e*^���>	�U}K����R�TCv/.�0����'��w�j��W��Nb݋$����H��w?$�ʥ���J7]���κa��%��0�T�F�RnXϿxr���xS���V`��(?s�K<��=�I]6�{���/���3�ܮ��]�y�����>�c4+�r235�i�
��Z��D�?��2��	g�
c�Nqљ8���<�(��R���Gꔻ���<#�ʓ���Y���b�3 �Gi�O7���5C�9�">Z��P`�����A�e�_Zm�=��ĺ+ڌ__��j��?�D�g�?����sS�f���|���1 ������7Jd�艴���rUc-�"�<��7�@t��B����)N�~@I^�5��Mt���"e�,�2�r�AN�/����$R�XJ��6�d��0��9L���~.P�+%���	9ލ�AÎJ �;&���z�I��{!��X�Zh#G���i�ycvT���5����T�k���]�Ɠ��FW��v�Ύ\��8e��-��aR�A-?��Ld�ks��"�У9/�L��K0W�76R��DԲ��I����,�%9{1u/^��-�o�Wmv/�u��#Oc�cI�Ϸ:}]=��<�EP�3�ZIV�!��~� j�"�Y��8�uܤ��xU`)e*��6�QkyR�n�D������,�[��T�'!/>q�6kdMި���(פ��r����-Z|��&����hs�6�[��GL��k��}�U��½��j�a�K��g;��M���b����mwcAhw`#�#��(��h�3�x%�����L�l������{���X���uM+/#(mr뵂�J�q0(�Yn�8�,�u��F�����j�8��#� wn|y�NRM#7��M���Ȫ:����K���f�������}
�	,����䭐C�ε����.
�K-�is��^��Ur	F��i���?~5�_��f��{{9UF{�q�Lm�����A϶(?gӅk�ڦK��b��ácKp/��3S��77�v,�Np�W�M����Y���	��o��)�/>ui76v��c�W�(��J`��e�3\w���r?a�U��B^���LV�	��=��W�߶X��NG*��������z�.��8��W+i����7\��in�OO#�3��(�����P����g��v��:���El5�W�C�v�E)>|���Ue%K����Ku�W���߫XL����57����t8�q,���j�3t�?��d�����8���Ɯ-���jd^���rE�W-�헩��R��8ԃ(��[P#�G��@bn��4���Rk�?�B ��$�Ms2ߊM�������yDɷ��?����S+׾�e~����}K.�֞E7�J*�Y_��	|��W��$Z�08x��~���H_3��9L٣:�>����Q�@�#��=�q�EA�-�RCA��VG|�8�+WI���zl����c�E�D;ەy�
G'z�����d�va�dÞ�Q�[l��u��|��6^g��+�r��'�ŊȜ.�����{�$���|�
�BI��{sh�؇�꜈~���nO.�D|,���������ܖg��rJ�⼍e��U�?�-��w���s n�x?S	�E�Dz�zw|0�:��aJj����BJ��)����*�k��rG��#��Ƴ4Ҿw���"�wq�̀~�ʄ��I�2���Ɨ����5��%��H\�E]!�Dpb��G�Q1����UJ!t�4��>�Ƥ"y5 %W��;��Br��l���]@���0UG��|c)' T��~�
�{	z�A�rq2����S�ia}�0�W�yC@���K�¶�KiIB�f}��?eL)���--��^��`,Z�y�(��`4�Y e�ܭ�S�@gfa��8S�S�!"��H���}�i/ѣ짶�=zo�Yr�GK,�8|�NUM��+�l�z$�^Sr�KՑ�T_d�h�#d��{[����|՗����pjt����e��3Q�>>*�1��tK�n�̊�]�kb�5zf�;&n�"K߈$A�i��;bmUw	{��^Zu���eC~]9�UODu�����;`����n����&=o.��*����`�����Uw�
%}T��}�\+%]�_��+X́�q�*���:�������g�(S�>B�E"Wt�Stm&7�:��}ZǔP���e���D�yc�Qo��<d	�!u�9@g��>Aơ�\,�Rs�O�$��X�q_g#����B�o~c~'|Pe�~pBa?��s�r�_��gv2p&�wP��c�GP&4��g���6��14)�����eK��1?�	�F�N���v�o,��	):���D&,)9�@�����k����>㻝��$
��Hh&��S�$J�t�WE9m*E�l�X��'�6����i%��s��g��]�.����4n�i�)o�P��D���Ip���M�Y�y��������5x�ӭ&` �^���Xbt�y ]�!�G٩���4Hhv�<���l¡-&�DWY��]C��o�ΰ�"a��/Z^�6����5�5�+,=���R�TG'8�o}�qk�)p\YW�|&#��lvP�7?Y|��(�1oG��X������nl�e�rAg�-1�y,sAhw���v��d�~���5w���W����,�!��;V�C�ه\__��B�Z�-�����A
�#�*$0"9nVZ�&�A�Bq7Q[�����
�U��!�,�oz~��g����f͕���[%���d�¯�������^��p�24�rg� a��b�;�ྱ���wik�����+����/w�^�z��L�}����m�4(�"|Y�K�	[Rp��MxɸI��j%��²��00����2�ߎbN!4�@�y��0s��=�s�)bSi��&r���׊dg;�o� ���T�q���e�L�� CBHfP;�p���	X���dS��_ӕ\��PQ,��P��Z�7<c�����V/����> �5g=}B����VwqlA'��ů{���tp���,�6���Y։=����̰F�'�_W��x�@�	&�K�j�$��*�	ك��o�-!�����v��l��J3�w�
MxRq�޷ٸ� ��(@��[~�$/��[��(?�m��7gI�h�e�̥.����ߡ)�!%*	h��f�~�����d���Y�7�<��� ��1��_l%t6�O,���K�-�G���- ؖD
?h�ݴf���vuǣЫD0�R�P>A��ݫ(җ:0�a|4Fy\O�θ/ƨ��pG�[T:�P���e`����t�IKG��=�#�Ҕ�Ow��� �j�}b�A ��U\����h��m���0ZB��l���1k% )��sFa�7U~|Lr4��!��L��W�3O�`^�G;��Tt*&�<Tt�\/���,�;���n������������
��Q�)�Trô����U�L�Γ��5x B��� ��8��R�}�����j<̳5��� ��~Z�
R�'���Z�� t�<7���|ED�@]F|	4�77L� Mb�T�,K� ����2��G����j'|*�#?@V��%=��
!��}�!\�?��6:a�<��=������y�nQ_B��_���_�������i���L�HZf���N� �6��H��|p�Ԍ0�'MٕY�����( ��^��5ɱ9aip�'�IA���50���Эr�ݎ.�5��:�7��ڨ��3�%�O"��	�Q}�]�sp�=>ߴ�ţQ6��h����jU~�-5om.�&n[�D���~���#G�x�K��� �d,F����Ee��?�+�H2�[�T̪�&�uӜ+����(4af��n���iNY���\`ݩYCSLT�xZPɶ��J�$���B�+��0����>ҹ�+�"���|O��U�[ �!��@��Q�p޳�ƅUo�" ����" �vߕ=��s�Ӓ$�m��)�Vs~�Z������w��GXLM> O�ۣʌ�O����`���A ����'zt$G�C��RQ!P��nr�?���.���Iآ�u���,n+���E��X�5��ħ���sLp�-* Y���:���Y���?�`�x�H��YU��c�ݰ5̖F�#$�?[�ZW�æ�H�*(!�{��=J_ś|6r�9��{��,�aY�������w���_F#)�����U�lp#��d��"G�b��`X��tN)Յ����u������<1|FUs,���%k��
�}Q�=Y�c��b��۟lӵ4G�-޵!z�.�o��'��w�a�����H�0���i�r
�����(�~�t$m���ޯ���H�s�ɹ�e�(Nb^"�c @�q�,d����K$9DR��zX��Z(�ll� W��ie=�m�.+�{f�My�k�_�2�ƙ�z��bb���V��4�;��ƪ>.�C||]��}�Ƒ��.r4a�3��e�:�?�����)7����o��O<��ނ��7����I�`R}K�t���͟|�3�l|�����2tYI�n�ތ�!�K�Ү�(p���Dk-p;MD������٧]��1�fX�/��%�L(��q{�|�l((�!μa���i�4�_E8t}�x�A�%�Pz:�ݢ>��QC����z�af�*~��Q�O��.f�����!���,��Y����ްaba� N�Tw�/fA-�3P~����w�<�*j@}��l���K$�g�]XaZc���IuyW)s]�܏� �a��d����Դ��J�3y��������A]�[�(��慌�R����;1�z�r�l�F��A'��^8�u�b�M����̲ƇG�ǆ��j(�T?׭�A�oi����5�	b"�A�f��1	,����o�����w�$Һ.<s����er�W�@��)��=���a���N᝕�d��)�ǽ&��P 6S��C��=@���RС;�JC B���Dx�"�p{:��;��_�2G��.�kl��n�i;ì�����KWb������c�V,!��N��ڳp�C=.��\�<d@Ĝ<�ك ͨ�6���8`�@�I���\��
��n�f�����:?!g�G��0	x��N��-��s��~w�/4�[ڴ��J��s��� �\��W  �pb^�WX I�̤�����v�}�z*���w���SIOw��:K�u�'��n��40Ѝx*⮻
�8��_!���+~�R���0>Gw-�.�W�����n���/D�P3����c�b3��v���}P���y/���{Dd
7� *Nc	_��{�k��N���I����6h�%�p�(\D�J�i �ũ1JhS
ް��@T��H�K�A����Y�(cC�s�M�|�/1�Q܋��e�:^�z��ιKd2�Ç��E��M��t��9#���0���홁�)�M���U��_aE�2Q3ZB/�OUc"E(;��쒙b���u&�! u��ly�;�����cX��2=��!;��\�<BX<U|�˭��h�Do��I��ax/�8y��W�ȶ����Pv���X�!�E�^q�rO�8ݹ��xI.O�[5�Oyg�qD?d��9N
�#�����rn�[5vO�9�S3�-�1������9`����{B��0)�RxgY��ɣ����o
X5�%�� �����hK�f�Z�?�m��5$e.�1�1 v:r&��Ld�[�޶����8|��A+�r���G�?:SR�/�@��p�Y/a.r-��V�{�7��#��LK�����x���7�݇�R��|��`����@��2�>I^Ӷ�z����M��L�r5
��~t���0�h8�ि��z�]ph��@3���ُ��?78|�#�)��+A �CF�gv&�TN�q���3;���0�V��9R�B*��y?�ѿ�pR?�^����:E���"R|�'�[yE
I��1Z�I!�I@3��|��0���:���,>�UliJQm!�f)ɷ]�O����𓌢�2���#D�S�1�&�?�}�X�{&)��--vǬg������BI*�SM�Ӡ�)m]ϲ}��#|����e�I��E%��k�&^�8����L��逵��'��L<�6��|�-!P&}�5��^�tI��cgK�-��!H�BV���
1)奇������zkܦV��8�9%Tj��h(���9W��N�մ�%/�=8���,��
�_��<4D�Y44Ñ��S�Jͧ0����B��m9���R�9x\&ұMxX� �,����2��I��`�p�4�e\��ǩ���Ĺp;�����`�ad�k� ���OB���V�W|T`���z�5(Ia{N��GZ�=�_$���]�"8���*~+Q^ ��K'�'E�V:-F�C�}�p �S�Yk򯦽�t$����C+���d��7��;��+�]a�a��
'r�rY�l�(����jn̑�Ieϲ'� ��K�	�E�,��&ˌܜ��sl
m��i��������|0�9������2G�Gf>�����B�m1&��k1&�9">&S��7n���3�#+�R�ҩ����|�>��i�<��*�g�����+<$�d<��X��8�4n�O��}�]:�V�����d$Ʒn�G� E�	F d����2Q骺�R��/������2�H�F6-����������#�J�Z15���*�a���>~R�� �ۢ�#��<��~I� ;�,n�?6������oS��j��&��e�*3���w�3�N����b[�.ceѹ5�#��2�q܅���T��&$�&��p��l��;����u�A�K�t��h?�Ci`80j.<8璿�;z�6r:���cU�V�>�&
��f�;-�
����ť��j�O1&�q�V��!��4�9�|��m�]j�����u���(,��ӗ������y���J]#�D��X���"^�Z��0�x�'����Y:]�,�B�o��Ͱvv}�p���Ś�&P��(�<�X�	�ΐ9���%�e76��??J�k��k��X�]@%�n�DqJ�r�Ø�Q��;G:�C�2q��/���;��`�s��s4�D�:��k��UB2N(���� ���l!�Q��&�h�j�]��zK���%]YF�Jh2�ob��Φ���;��8�܅&���~ѼD�4�9���;a� �"��ΪE]bUJ���e�$.ۥ���x	Uܚ!�eBN�����M���)���RIW�^�K9��T��h�S(�V��?E&3�z�x��G�����߶$�u���UtU/�����V�q�-M-Y����"�\��[8KtZ�����ӟb��e�e;1+Y쬑9�n�Iͩe�i��Y�ˁel�U!ch[爍<�gJ�d5+Yj�spS����1�I�;AߩԚ�|#Iޛ�#1���!�+ ����]E����P�cp��s�����rl�Gs~�}�::k^���?7�'���YA���Il����>z���b���ë��̹�욅H�������-�,�٩a��b��Y�z�&����cOl�,w�kKu�u�'����yL�������l��A%�sG)&1.d�D����i��M�)\�P����T��A�Χ��,�gS����̐���+BL��Z?�S,4�`P�+����mX
�}D�
�#{dYqVF�#�Uv3�G�:�5�Tޑ!�A4�)q箈˻�Wm����g
�U7Cƣ�j�`�RxmH��Y;F�	����)�&�ˇ\H���l����f��^��c�3.(�:Ӹ���v�6 �@T4,r�bҢmp�J�"S~\���	�iT$u�uQ���Q�<?��o�z��uv����i�}��I0��"���}L OL�Ü���;Y��A�]b�^	�#R�R㤿.��>������
n�eI��ث�S�+Ub���]��h�<I����t�@[#���.$�����ӊ�x��A�^�H3��'zn�~f�����P8Fi��x�;��H���!�@�H�B�Hٸ/P���u&M��	FϔIޚ���R��9C4��:s¾
k�T稑,�G<���jd��G�3Ely�7:��b��~�Y��7������s`�,��Z(|8w���I�vT�[�/�ê%.6O������6~�W��*W�÷o2"i��ϰ��8M�����
��$���ߜ,�H�遇��7�{��cv{��H���c����~v����W�W���0g#�1ǰ�|�YXι��Q��^��ʏîI˰v�P5WCS�U��Ú���\y�r��E��ި���C��[�Wn	���_��z >{N�_��7T,a�k$���nwm�\�_=~�2� ;�P��.��������𿲤h��{�eB)v����D��s����G��i1���
;ZD�Y���+	�!�RW
h���f��a�}?ܙn��B���93�jg������4��� �|	�Z�u�?ڗ��
zb�OCVFw�Y����6c�u4S�+�ߡ�`�!`k���`¯<-��N������`�
8^2\t�ao3�'\�{`|�QZ��9���A�By�[��jƂ��qh��vjy<���m<��,
Å�nAH�`|��kE���sQ��0����"��Mb����	E���M3�ʑǡ xgy�1/o;ճ������Sё�rt=�jŝ&LC�2����!r����a�-�`3��'�� �Z��[s��z%3�̷w�\���ܩ����2P/�OZ)�c4
#ŹS����-�2�V� 1����} F�����+���n����Z<wwh�
�
���9u)�8X����	b��A`8�L�ߢ�5`��8QZNq25��c�A�_@��Q�� "�mYa_\���i��Z��,���<n���ĺ17�a$�D��X7K����	�y�=z��.W��r����z	�|\ӗ����^�C�s�ل�i��UCn�,%O�����;b��*ceJ?Pv�����8h���)q,��������R�)�V���S�?y��M���b��9O�)�������2�]�׬�,]��b&��X���y�|����۩�KlAǙ:|eM�IE�����!^5�X��Nݩ}�g�B���'.=R��S�6/VR�Q迓��'7j	�M�T[���@I��������.(T�27�9\�#c9S��,��v�:!`�}'~s��=<9G�x�g+����u����&�S�8��3zƪ���/i���o���kV���ȃ�DE֗�u���\���6N���aWC�k�9?�dDc�{�r��BǛ��G̵���ԉ���O���ƍ�, V��"��9���_q�*��6�h��lm�P�8�W�d�ו9��+�&���`�Q�`��:sk�Ui쁕�ݙl��H�,�)�p^_������7�nF�Ş�"��_�:�x�t(֏�I	a�p�G�G8�-b�ѳ�Y�2�, q�W�=�R.v��>M���'��*����~���5'!�y�X3!����¼��0kܜf�m,X��i=E�ҭ�C��C3>���z�JG���8��V���1w��}��ec��ӷ����Ȇk�����@�&sK�ݯz��Է¦2��9��0B�+@S>�˗���*��v��$�nf-���rA��$�����z�s��7����s�78>�;�Ţ�����h������1o�4�ɇM�����N����O!����#��5]����1)5�)X�:H��kz#����~U5�$�� �嵷Y�0�i���Ya��2t���⑧W����0nQ�j=�s����� ��>ӛ�.ЄC�1�eFϤ�a䕿|�6���'F�dWـ��V��g}��p�m޼�t%�E�ph��!�6}����~1���B��,�3C.��h�2�.f����<Q��j!�Kv{YWu7�4�#��ݽ/���>C��~vW�B24�� ��XfJ�9%(�K�ƈF���&}��dP�c�q��!.�3�&�	�D��8�·_�Т�0w�W�sO��Է*R��)K����DQ�-����L�7�.��c@��b�v�8U
����DۗVi-
�J���]{��qA
T��� �W��ٶ?��_G�"@N�Òk���I�	�Zq��B��~,�Lļ����,ĺ)���1�t��?�j�:>���I�x�(8KZ����;Ȥ7��$���|� ��~���G��~���1�l���0�\���%Kǋ����'(�	O3��'.�6-u$ky�A�3G�;�!�nrvE�����Z�T�xWO���������}�9u10^A�oG�7�8�#2�����9t�ª�5��Wt�A��!S<�N8�s&I�|T=b5dڭ�=�	�'�l���� �jc5t8��J�0�j����Ҝ@�K��$r��O/+���i���
v���.�]p`�i���]}�Aρ$Z�s�hZ��Pk�L�#��*]$s�"*���a�cӟ��&/�cG5wQK��� ��;uiG|B����Ū6���Fe��0l�<mP6R\������1��q:��D';�S�D���&p�ɀ��۰�QC������	:�?��A��:��j���h���?=
¤	�&I~|�e[B5�-�$��ql'�UدN$�I�w�S�q�jS3�}xbId��.e�ԑ��d&\��AwmO�F����Hh�E
�L3�jj��}����xp����P�I?��$����$�A�ev�����Y���xl?E=����NA�T���S=���8�GTB�xN�|�3/�=,\ Վ�T�9:d��Ʒ�d���Egn1�+Gs��Xn7�K*B͇It��J���R�/g�J� ���~ō��%�=ofD�s2C�4�A�V��ǒo8��i7�W��	���_���$[�j�x��+���K���`(��~S���ر+���>@F����f;!�ϐ_�[-�Y�0'������B��@�"�V�C�l�XW�y�A��4�yc��+#c��L�a�/њϫ~?���C *��2����/B�q���Y�=M�NgY�������������8��}�H�y��k�g<���v��i�p����0���N�Vn%�,��{#��x�69���/��Y�nN��2�n�+���i�d9�bK�(_����ZŨ|R�ńA�j��2��0,Ofw^N��0tǁ��O(�����oj���d��S5�o�^P�}�HA)���tX�q��o�-ޭ*�xj�j����W�O�\�_DWS'R7c�` ��/z�%��#N2�O��S�������B%��ƀ���t;l�t�t-�fK��(���m�eLhWɁρ�H��v�7 �,�S�a��<��6Y�h��x()2�/{@��>z���G5�(�W�њo��g���S��<���'�̧`~��M�rF>K|����"�����#�<R䱟�胹mw���{^�Y����A(X03ǖ��J.�'F1��*
Sk%����px��u7ɒ�8�G�Z�i�f^�r�ٴ	���ȋW'�<�%�LB�\=�h/�a8�w6p�q��Ϙ�j-��Y�l@��w{_�\����D��	,�Pܟ��e�0�sPqػ�˫���f�/��M�yra*]�� 2����Mx�"�����B}�i��g�.�S.8D����ʅ�}��w��3���N�"`�.��W���'���{-
��D��N|}0Rf*��!���xgM�lڀ�6����f�@�E������b&=Ui
�C�>��LD�׶�fu{w�%����1�RCJ��	a.��f��MV��S��n+�x�v�7M�xj+I�ᴵPY�H�m��x�!"��5��i���ux�$v�0���8���TT?S˻Ʌ��ᇽւ=LZ|��
�R綢��3�1U�7��ޔ���ci��w�k�&���A�{�D*��^����b �W��J+�S_���,b*&Cz�e�d��e�T�²q�x�4����-J�4UF�vם��q���=�O�� us�,��h�Φ��C�G�Ձ�[e	({�~*���M���#1\c��ɲz2���Z�k����z�dȟ$���8��$�4W����A������(��;�t��D���(|鱘�w�o��;	r�m��Sj�\ /a��@����Ea7�������&�t�y�",C���D��,f*�4��4~*[��S�y󴳰3���&j�Nf7v�Ú�"A �O2��=Y��{���YG���o����s�#1,{������0]���z3a^�bL3�D�[\�7����`ӫwV�Ho�̦��J�0+}\��(ъ���~X�^~8oOSY�9
|���jP�YL����v�����!�.�X����Ǯ������_�yN�W��Y�`f�1'�]�� M�w^=%�h]|���p{[���/��Fl�,q�h���1eBx�ض��ʄoh����Gt�x}S�	�yK��s]���^:}�e	�!ciu�����i�9�����?J�bPX�1٫gN��s+`�YR`�B\SJ�˽Z��I�O}�7�zJ3#�d��>�gJ$S3�k�}�\{r�����pbb�Hˎ��d��?�'*��8����d�ß�ܩؑuE1]7��J8caĠkM�Tr*�H��;�>`L��j�"Bwj��`���	%5ǝ��мW��w�s0�	��A����w��4Z�*>E`d!���O79��Rg-�Z{�Uq���δ�q�g����gB��pU`_�зpD���k���غ�Jp���.�B#�V��yW�^�L5���\��x����(�[`<���@�}/�"�^A���z��j�5�C�4*�
o"�ף�W�v��D_̚�a����鉏K
��&��c�����?�����B1�r���72�� �j��7���ub*W�JOםG�I�r�A�/NR� �����#p�&H�){]@��q���P��H,Q�f���a˲���w0*Q�7��k�`�;�G^�M����pF0���y����md��A��1�@��	�j"v<Vۢ�/̌U͟V�#���μ1\VD9l�K[�XR��:��6�3��PFv�^r�aɬY}�=4Z�'�u��&�#T"�/g�����ǏZ�)������8���h?�5 cBJF�i�\�E����*��`QG�{,�|���{P�rӽ���o�Y�����ʤ<XZ�'����z誃���F�}n��X�����4C��˄S����ϳH<XN�����u����B�F|�r��F���PhF5�"'�T�/�qB��i� X�U���y���j���Cz[�y��(L��a�HC���+Do�Y��m�੹�=�1؆%uur'��~?H�l N��>��R�o�T���nR!4B��*���Qj�9�Vv����yC����Dִ��T^��G0v�5�BN�i�F�3��0�Sֺg�(1�n3�_��㟔�(��R��I j���k��+5�o_$r�;6���J���#�&(�Y���@l���YԐӓ�"D�*�\X�fq�|�^�
�;�B�3����cൾ-K�F_;�V.���D���q����g]�p��b��/���A�ҷΐ�b