��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��S??Gl��4�͌^����>��͡7h�`H����a�.����a��bFj֗3p"��@�{�@]{���U�F8LK���L�׶��(-,T
Py!ҫz�������7C�t嶂)�>=?��M8���9���6�F�sm;��H	g�58
���<�#v� �'�FF���on�_y�ͨ Z	� ��ˣ��B�1�:ϲt�r8��-FЙ����؟q|u��=�-�F��G�g.:1��O~'`:��bZ�^�0��Q-��<�ϭ>Z���^�J�/����:.�p�C�0
�l�:1w��"�`ށs�$����dt}Z��w���^��M�
2h7n����+1�oM�O�Y�t�O��	Q^�bh\x=�.P��4�2���8�c$R{�>8�ϧ�&A%k�Wk=ml��,2�.��t��^�R��m�����z�v��r"��R���T+"W����'�h��7��:�e$��J�4t961�������N�v=4J3q����r�߯����6ak�W���%(���+HAk0��vᠱ���V����(a8�7�gíp=��J�vc�.2���#�'�&��������,�����?�`		��@?��lp��E�3��b�b~�.q�J����d���ju���	�m���9��& ]�0���)���z1�����e�g��3�yʧ�춵�	�y��e�B��6	�h��3^��q�\�"6�ٙ)e��6޲"�՚�L�+$Ʀ�_�������"�-��Q����1	�%?��d���T�j^�M#��3��fD'��Hy)l`�g����^�[��Yw@v��EAY�-G�goa���2;����F�`�jvC#f]��H�tc�U;�^[G`��wX$|˸Y�6n�u�u�\[;���#�W{��U��v��������#�̾�:,D�.U��㷗�j���T����ۡ��j{^nO�y(	s�dwΉ�}��}U��ϰp9�hBz��r�K,@��և�1_�+���LF"��Xs��O��0S=
'�ܾd/��wq>.F�E�=k)%I|�����򧊋��kf���.z% ��#N#�g��K�g�&Q����b�q6w֥���m��F���6�l�1�}0���Sܶ��x˹��	Y��57���g��f���d�Z�ÖP��4b/&���%JN������8�emy<Ix�0Ǹ��Ą �芷^�.�MD�Bxe�~[� �`\�\����ϊ � @0K������}H���^���\�aR��Z�D$� y�C-�sŒa���aD.;6]�-,�wŘ�Q�Y^�!~��QL$��Z���VvE.o{�M���KhE�8�c�:��nȀY�J��@�����E�K8U9{Px��CC����(�+�t>��Cf5
�L$����� ��=Ssy��z�߈:�V�C���X�
���²�$��3�r�~�����Iq�
1��y�b�L��F�ua�q�7��$���2�aS�qr�E\k�^*]��2{�-Ȅ�y�P�y��H�[���Q���2>ԍY�"_릉X̅g�қ����U1],�OPUGP	,�������>���>� �|1�`v��f�d%p2^�'!w��/"�!9ЏV�
����p_Q�
�WI�1تB�9�"���a��x1������'�$̫b��:���d�*�m�E;f�u�U�a˴и�u�"�����1�'�X��s��S��	�2_B����OI������O�B �M�,4yaN;�pv@��l���yR��,}���$�T���L����=jւKb��3O�E�|������z��+��d�W[����G��*� *E��f�J��	���-Ti�2TmT�i�&��S6Ռ��9J�E�Z��b��Y� ��D��e��+��kX��59v��3���v�➬'n�>�?��qF��˸������1$7YB3c/Q<��}��U�n2��v :��4he�d���=��M9�ws'f�6U%����lM"*j�%�:��6�8h�I��z���ܶ������b�Ҙӱ��� 4�YϨ��x8��BJ�����K�}D��*�1O ����7�u�*+����`�3ƻ(�]�;�3��G]3�ф�6@xv�n	[���đ ҩ��^�wTD�����*d��=���	�H�I�����7��-|)o�?(�cQ�Hm�e����Of�LY���B��P�9|$��n�
0�l1�j�Ȇb�|ˍ�{�q�+��#�/��}�C"������c��bOx"�r������s�Պ��A�Q�𸾥U�w�Ж��p	�7���n4W$VΧ�!�-�Z��u��>�!&+�4V�]jl��l�Vom��f�Ǭ�_�G��,^�� ��� ZV��?���AC�[��s.�I�gSuǟ�a��U�6�JX;���8�y��(���b��r�'05�,X.�̗��B��d��ݱ�	�'��S��H���h�ܾ�p*t^��y 2����H°iw�U�ǏE� �T%��
7���:��F㭽K||�ݔ�9K�Q"���{�}�ˮG� \�GK8��[>�l ~ϓw-��♵��]MQ�{�����*"�k5.�y)gM���c�Gª;�VV���rsT�oKҼ#�;�Ĵ�e��yNn�b��x!}	T��
j�T�d�y��l6MqUֱ�C'���ǎ r4gV�[p�g޺�L�BN������Sè�����8O0��C���͝�x������ms���.C�ݠ�3�Ҽi���(�Qo~���<�>�KVD�����	8Z���y���k%i������CKW�o܈����UK�4����gּ� @ߙ��z�#F�W�~N��=s�_����na�E�h9�*ia;<ɶ����D>oz-�IÁ��WԒ7�0�ĥ<�*�7�)!��u2KK�*�m��3h�M�hߗhQ��0�}8��6��U�0��T9���$q�_�+-����@��"�������`����!c��U�~Ax��L�IgQO�M��
�;��<oGc`�����S�+ӕ�yA
��މ7jj`�zi
?�(��c�>LS�l��u�cV�F<��U�s��Dw4w�C�'3�4�����-[k��S�~k���y*���q��%�*QYQ$���A� IJ3��V�L��v3�C�8��XT���3=���(���ߢ���6�-{p&�Vl�����oT��<zgAh�'�U�8���6��J"=/ּKW��!�EKZ�P�h�9��P�PIZ�ZGo����,4+O�F.��=�p������Y��?m�E�p�Df���:��3$�Mns�0���f��txv�a�O�H>�	 A�ؘK><�މ.4hik_�Egyy��*Q��+��u��Ja������k��\�G�z�e�2@��{��Dh�����y����P���~ʈ�<=��5=�)��ؙU�è8�>���y'�&i�䄪�ّ�?��Uf����
�㾧U1�
�m,̻V��� ���P �������{�'Z���/���[2l�\�a�9����6��%(�>M!��V�@�	K�-~Y�ဍ^?=� �Z �C#%�z�������1��hm��a��w�-��/\��7���3!4l����z_��G���E�����Àk��&`�R9��8�N������^��)�� `<d��}6*_�!Y�U�"e`���(���k��'׶�����!|J��2���f�	v���p�1T{9êU�){)|���}�����Y��Ǳ��)�v�tT�9�걹o��R�;�ã;�=�Q[��Q/�k��#h�;k$�u�#���V7�"xG���Q��j	��(1(79�q���{o������-"Q��ܞإn�
��ڃ�w���f��暭����y�\xɎTaK6ּ��D<�\������r9����y$]�*���'��5 4X�����yO����LU��Z_�ɨT��`�c��I(�`b���|>s ����H���{�5eg�wЀ�I���2Յ��u}�/X�}C�3�.�l��b$�([N����y��ڭ�������
�Q{G�n- ��Cf�O--W�7Jtg�ί��T�������~HD�6*����JJ����D���aP�R}��
C��mM��R��B�E�$5��/7�w�cQ�DEhmBv�Kh.����,�÷�@��[x���ye��%���Hw����8O�#���
�r-��K{>����ܵ��u�7L'_�֗#G��Ӫbm�=�O|y�����q;�֦��vf����6�ھ�14�va!��k��~�$�n �?�N��Ǒk2�c��WKL�E;�3+�V�6m�ݩ���~k�_�q�y2�@=V:k�̝���Y]~�vG�3�}��Px*O|����Vm��h�־��1�ʉ�0l���6�)l�Qr�]I�:���n�a�l?�m��# � �-���o�dBe5 �Ӻ�g�/���hl�=�׻ny��@�T�v7xFgC��Msn^��FX۝#�ȹ���`����<W_v&��"6�^�6���"�Bc
!o�vK��؎%j�(��颵�?]z��P��pN��s�4�$[в��`$��d��L	�dCM{Vzmk�ܤ���ұ�M����8g��
��2|Pgr&r&�{��́j�*��7��O!	r�\`�a�)�-��.�h,]�*a(^B��7چ+����4�x���~�Zgت�F�]_��}�9]@����1ުiu�� ��`Cntm�a�[��?X�⫸�z�İuqm�ՖGB�U�>�̛�X\��x���#� ��d��"��̊��R�҄�_�O1�~�z@�K�_-���^�,��&�x֭쩖����?��+ns1�ƚ�zQK�b� ��i_؟p}y"��w��`HV�/e���=F �W�1���ھ�O�ohS*��ijY�#ɬ����f��A�5$D�+c�#!ڹ~�{�q >�|K�x�m|��f����5�daQ5o2ޓ�����7�7�Gq�&{��5���t,���c�����}K�ҨA�����,��q��a�2G*��~�BÙ}�ļL������qq�@�i�%��5��l�0��f��Q��H����<�>�L4���O��u��ߗZ��"�����)N��5�>w�?W	ٮÔt��D�D�<�`dc١�������c0
W�U4�O ]���mޗ�b[�3(���d:R^��E:h����Km�50f[���=Ό+�g)|7Tz���2q��6M^H��ݑps�v�)�����^��wM�4��O�=��{x��g��s�]�>t�*��_v�i�_�v����A<tf!���d	5��ìO����$�	�c���!��#��M�!�pQ-���$�g��I���㕻q���f�h�Π�G|"�aC�{�Y��v������r���yEU�ۉɋ.�E�_��#��C3���˚����2P	�_�
���ۢUgA����1�J�J�6x�
�}��[�[����g��t�o�G��Q�nX
 �zz�6!���Y�}�����+��|���eD{W;�-����6��D0��mJԧ1-�7�UVNM+0�
���	��I�k�6	 ��2�:C�������ſ�冶��!P�}h��sI�0��ڛb��-�^]%����M1��o�@	�&�M���G��H[o߇�����-FJ�H�u۠��Ր�(�\�̂�#R�ܤ�7Z��#0�ۉ�+�G��Jo�@8��|�Y���8��K=����a�U�U"�3c̱V�]Tm�[���7ǆ8�mu|_�K�"7r����V�s �v�������|Y���8
li��5��������;1�W�l%���l�0�[�Q�66��_���������uq���e�T h����������i���lA<L� ����_J��dZ��x��yVta��`�iJ�K�V�����POnZ�ޕo�K�g�(|�DA���$�xY�UL}!�2d���
f:޽�f����Ɍ�fٱ�G*W>�"�2�>.B�#�mȀ�kqĢ��P(?2�W�$����R �~S��at\�)TjlbQn�UW���N�}e>���v���
Yȯ�*�rZ��)�D'�d������a�O�Tc��3��&�Lڤ����u�\��懹��A_�͠7�X��b`��kV��mH�6��/wc+y�ւ^=�%�)�spdg�b��Ld趆[ �t�GBΛ���6�֦���|��35<	P���J�I:*&��eM�	���NKz�,<f�M�U����Φm@6__~%۝�ֽ}���̘`s$ɍ��(p��E����<��3D�����\�ꦸ2��"�i��
�{��������ў%�����zC�{uߗ��8��ӷd!��9h0��� �m���d��^w�7���|���WɬTx
�5�F����dZ}����n�%�}7�<��+�c�a,�h�`�m��_���5�0䩂�3�	%������+R��t���$n������O�ߤ��/n�b/��P��Ыg����3# p�vd���_�mS�DP�����½ş�Q���bkSRy�{Ddt@�#�9�}����h�ʃ�컂�RK�Y	���$q
ex��<�
W� �����h��E/�Rj"<[O#ݼX���g�*�e��6 �H�03�$��i@H��|$�o�|	�#�oqC�5G��4���_�U�� �3/Ā����g1Y(���t�6ƴ)y���TZ�-zV�b���p�]�6��s+�ic��
�M!�gA�2y��E�u�ç���LB�9`z:D͙U��z�޳��x*/�Sՙ����|��B�s��Mj..-<�lg�Æ��jV)ʺ���ɮ�?�E �ള�1��@Mr�ō�Grm�ߑ	�v꘵Q�TC���ؠ��f�*,F�#����4���T��~��Bbf��������.hW��̚�Ψ��I�ڰ+_X���q	I��A��PL�%��v�o�Q���j3��N�������;o-���0��C�B,�b����f�A�E���e!��$t�8ya���_�a ���T���W��6O1}I�!��^�F6�3�%�죷�mH�Ƴ�w��D�	"MFyW�{Ϡq!���&�q���������*�B��͛����a$�@P_�ʈ���P1�-ޣ�wa8����-�i�XP씳36�Z�O7&h�|���d�g�:�r���1�ɥː��ɬǳ�t�#W�M�[׏�h�L���f��U��񅽊�3����]]Hh�5��D�y`C.��%����M�AqB<���M��P��	�B��cPċ&�U�4t|��n���89��ڟ{iҾd�uU#��}�d�1�/Ă�bY	�[XY��WK�ͯ],@:�Ji������]����OSc>��V3�SwG%W�J��V��
@.�A&]�=O�߻��C��+�3�Z�gd�_�l�����Dkj@��鿦��d��FVJ����I��j�J�463����vn���Y_Y�t���������,j,�ɂ�x�h���b�mzL	�e�Om�HsNE�N����o�Ȣ ��k�g�Ytf�w�>�_��R�w4�WY�8��	%}a�1{��!��_�*K����>��� ��y����f����oΉP�o$��e�'h+9���ӏc(XMT���+ݯ��x>Ѯ` W�C9Z����LHm';�ۼ�i���0�D�7����O����mdjpe�//���X-��T��hw}���u��_3��A��
'�����S0��:#�$x}����b�j��Ɯ�4�\&>+��wWٝ�Y��}��ғ�y)),$a�0�?)h,Q�Γ��Z�� �7	6`�����X7�"(p3�4Zh��X�<\̩*�h�;�&l�q��1��,�(�;?��R_��g�n']7�n*�m#+��n�s4ӊ�^�p+��ȝ�	�E�r�������iKqn�(ή��[�������I^��I��w��Xƙ�&.jlw*[�T`g-�㲛�,,%�O;_�Q��R�ic�>�	��@�zY���O�C!�lʓf�
�nx&2��3<�@��&۔��T�=� f��"����wLi\Vu敬�:�!R���Eb����VJK�6f��w?��` ��A NM\�}��S��B�5��y?֋�-}���ڳ�WA�s����զ���$j�t���y'��k7��_>oW ?���GC"	�}�5�u��u��7+��\T�WX}H�<��,"_�՘p�1.������C��E���su���"��K�Q���8ظH��-�+q���x\Kѱ,��j�t�[PB��\�$A����p�N�9��$F=8��?qM��X�. *D�e�.���>	y��ȍ��a��n�E-;�7V�L$�c���|D�5���'�.��h1�_*J<�φԕ���'TR߬2��~���=:8��-1�\����K��/��|hG��˵m7�tPlMa]��~�uQ֚�r�4p���)_ c�s�3o18���@�N�Gc��z+�1������ʗu�iC�x�;���#����ĬN���V��Ā�S��sV����'�zy��E���|Mv:���uB@
Sz� �6v@��rC��d[�{x�������X#�k!z�z�1=��q��~>Z�p�!��z�H@�`oDE��Y�i�y-Pt�P ���S1qo��hu���z�ִC��N����fw}�G��%�r�yB��p�q�}^J�\�	��0��!��o�%�V�U7�qE���Y�o&F=��B�:��P��߫z��f�'�/���bk��ҕʮOH�)�2�*	OP��:��,E���]Ɏ{�x�"�ȳ�u��ǣ������Z�9�y/(�2���<�h}é���U4��9���ݦy�@���ŵ�r��z���!����^h>�7��ͬc~�h�Qn�ƙi��U wZ�G�wt�l<@�H��͏n��\�I:3[����`Bc�G�� $ZZ��]OM��K�I�z��1Ex[��+�u_d����,��)����uv3��� �^}\_�<�r��!�L���ȼu�(Ц�Bf��������'s����E�xH�!1����aol_�'���a3&B�[=Jk�+����p<D7[��艼�r��֭�j�jNIN��1���o��!ľ1hTI�)(_�5ɿX���&��&�������㋕V���픣?��y� ��,弽�\�o!��35�b+d�	�r��F��5�#6!{��H�aB[���PQ�5�a�z=������� ��J��iLHW�Dsr(� TZBu+�A#�q���FuDC�%S3z?"G}��O����^!��Mhl"8\B��t��� �w���h�i���`$6��N~99v�&�V}~����B�J��T��`V���_�I��@� һ?P�<��Jd�ŵo։ �TXj2M�#?$�A��ω�lߥ�$/��C�[�9�p ;{��c��D�"�����(�����ү�z`l$NA/�����K~)/!\,)j��BA���n���R5��(/�X����7O�?CK�ҏZ�}�6P�%��$Kmٱ�k�gvg{�7����&��j���"s����̖���k��H}���a!Q��h��s�|�ei �X\�ґP�7t���]��U�2Y`l�Zk����C���,����b˅�
�24:V� ��<��!G����y��9��ԃ�M�<e���Z�M5��!��uz��D*a!���1��=
r��z�ƞV�fk{�
[geXi�a�P�X�+��-�?V�m7׉,c�N�hm��oZ+p�����Hcڎ~.Z��̍˽uq��j���/�4�Yꍧ��I)ʰ6�@d�{�H����d_B)��M���nջ�����)?蟜Rc*�C?Mzo���_7�s>5ܓ����9݋K�l.�5y9�vDP�C�J<MC�0��f��.���&,�R�P��=Q<��:���2`#z�x����6�e���r��Ӻ���݋�绎.j�>0�v��[uABF
7W���4��J/V�HF�R^��;�l��d��pT�X��2��B��J�8�fI�y5^PEN{��K���_I�8�0��ؒ��Y[�.{7�3��l�i}���şc_��F"��ޯ?g�ҷ�
-b\�];��UP���h������#�R� #:�0��2]g(ˎY��A�4*��v��G��˒%�W��1�2�+0���}��9����]~�0X�§�F� )¨#x���ɵ�N��5�����ĉ�Aw=^��d�S���^>h3
�a ����eB��uRv��^pR�QE�4�s$^���K�:Nf�⬆�W�|�pC�A����y"�`W�L�wX�F�0��e{�{=�?(�<��P2�g\S������U����pE������n�]��p�P�;Pp]����ZI�찍;X��f�����|�F�EcI{��5��~}&���*�e��%'��Dܢ>�i#�Cq�La|.c^�j9�J�,ь:����&(��{|&ԇ�g�I������v ��#�B`z�bڝ
	�b��{���ԓ��0O.Є���
zm6��'��2�Gb	ᒹW?�w��I��u��	]b	cT��:#]������d��������pe�ib]�,��y���S���;UVw�S����T;��Ԟ�F�o�g�,����/�~�pq�%�t'e7%@Y@�OX�4g�������ݢL���N�r��^���DTNB��Nku;Ħ�ٳ/]�Y����`f� �c�E����v�G�:��� ��š��-W>��hE�w���s1ќ�J�K`A��nbȄ�/�c��+V�J�(n ҏo��]ǻ�ӭ�V�c��<7vDC&�7E��%�ylXJ@��bI��M ��B���L��r�&�c�s�0B:7����a����r�W�2�BIR�2�s����d�������)�4�ԝ�AT�<&fd��M����8�S��&O�?
���Lɳ�Gx��Ch���$�1�{���ï�T����G<�[蹣����C��W�z���sQ�~�1�Lu�g��IVA��Qߣu�HɘXA&�F��R팤��%�R�󙽟�b��)��]l�&v����9�1ɒҡ�-����Ig�=REfO��U��F]��y&2����؏r�J������ծ��*��g�س��/[�e7��� V� �_�� 6�k����!���)I���<�fTl[CO�4zS�xY�e���q灑}��tk�r�9�`�����AZA�g�e�w�1�s���%��b�]��zgG�0��0��W,���r����^�4fw�x�2��a*��F]�W��7k����;6˫㝤�FuI5�k�l�X	��=���� ���z��l�-�
e�me���a�)�k\��!-A,h"ʯ�x�4Њs���Cw8	��jM%N~�2K8HJ� ����Fd��N�]�2n�hI�	���q*F�J)�`q9v=�J��4�'����)$w������?Q��K�ـ(6�f©��s+��4v1�`�z��C�[v�!|p̈.yH�v��%��I����e;�[�8����g�t�8Ɠ�r42�����h�mE5w�m3u�P�'�Nu�~M�OOr'ކ��i�/����,�߱�Eˈ��bD oN�Y���ر��~����I��b ���Rk�����M�9d�z�O�XXc}�<$����@B7#Փc��YDa`��z'�K����V���h�O�\�ŉ��3���$��(h�!��{�m�]��6P2�� ��ҖrMg��+�\o��Z�}�NHB�qk��/�	]��p���;�d���і�; ��x���bb9�'� -Ļ!��ȁ�O�3@m�(D�	\a����z�1,}vs.H�T;Iǌ;_�I�i�O��uHP��Tӿ��A�^^�Q�''/�c}�7WA�`>ITD��㨊���t����U	wy3v��Hm�-�m&<H5T���Ci���MR5�P�[ؠIO?0�`�-xvآ+bm�h�M,��H�+���
�a
r�?�q���X+�E?����,���ؑc����.�J�;��W��Ijh���h��r�%���T������r�`ȧ(��y�\] Ÿ��rŒ�X�{�m&{��٤�l֍v�	C�}�"nz��PYkLg��9����1AE�Ύ�;k2�pez�8��������R�EKGGt�l�s�K��s��|@C�m�8����'�7"��)�$�#����}b,8�gIEE�P�y@R,�9T����`�XM��[���������+�5TU��z�a��l�A9�i�H�NF&�q5=�D�Go_~i"]a�<���m�H�F�r��c$K���}�t���*�V�y�<|2����C���~��}���r��J�4���7 J���\�[F2����J���@$�5VU�2YϲE��70�x{=Fw]q͆|����c־YQ ������y��W�Y`����pOђqX�s_;�=�o��9(ɸ���OKٳOB��|1��͑�C��]t�I�����Kë~kX���T�G�.O�msx���{�����G|�8��L��%΍M"���O0u���Lu7��S����!����{�x��I5�w������b�Œ���T3g�A��v���Bp+I�0��o:��B�4�[���|RRh%�=K� 6:(c�~�ƬO<��5D��@ِWpo�p`@�@%�L¹�`��#@Jr�sG� ���S/�
����Ⱦc�=�_�����a����B!V�\��A�]���AG�M(���y�W�3�H�R ��pf>o����~�3$
���9I	���|�4�Ȝ�ɿ2k��u��}���䜣�$�8r��GO�#�`r9�z�R�V���g&}�R)KMw������l�@�!A�y	I��'��Y�ʹπ4�Ud�l0:XS�n?�����������sS���TD�q"�+u�B�y�{��JeR�H���l`�]r�E�Zsnw;����w�8y쿿=��Z�?�~�|�u⓶�����ق� �c�+mܵ�eK4�
L��;���n`.�i��׌`|��0��z [C��*�\d�U�Yo%�(;��k�;O��}��Q�f�����ߘՐF���a"�-�J��O�@;UJ���U��@�7�ZͬO�l�##������ż���XD|�EͲY�)���+���b����b*[0Ņ�s�_\��&���u�ر��o_jߪ��WӞ0��7 �h��;���|/5+dn�������<}�GT~�	� ^���e��R�]Tb�W�˯�-_V�TW�������f	���m"�jh7�z&o�N/n���ȣ+ᯢ��߸������N(�Ȗ��XNF���N���&�|�BW�PE�9�"���Zb$$���k�s��QP�h�{U���p�O�	��E��P�]���])�(���FY8�~��f�������KC� 1��G.GG]WrT�n,v�)p�)��.���%�q������}��]f�<����"���&6��BSr#�p�:��΁����r�E��
�O�bM���RT����E"G9��(���r�;���4ް�����
����%Ño,�uɍG:3�?fsM?iW�_��.(�O���)����#�[��&�S���i��ص�`7fT��?������6��j�.e������	�Q�>�e��n���ݥi���#퉣-9{�ޟO����E��v��~�󸥲eg������^���?�9�e�8��ӰO�0���bqԶw��#�ݜ(eQWZ��qc���YH�h��k��M��u��5"��z�-yih	)�~����L-C��S��z��QȘi�l���M-�� :H>��AC�בtg�p~��1}�NC�����.�/G�����c�^����&>�lߌ2Xx+A` ��V�j��g(��Ӷ���P��OJ�l���v�U��h���)���������̈�U@���n�U!���*�o�W>4�׿&�	d���FNe��i,p����xs3aY`uhZ��Lh�_?g����_d��2���y=$�5>�l��ݨH��M�Fcb���r��dQ��K<������W�H*�����/4���`���j��G��S�u�~\F����Ǉ]�( �a��P7�6֌[I�K�@X�� k�˙!���P_���?(4HEP���t/��׽�C�-�Pf��{w��y8DS��'G$Μ�Y��>��M%�y|;ĳ�O�<���]�SV��c�D]���i�i�S`z���^��<��lt�uK$;�6�RA� �y2�WÑr�`�@�W��MyW�u��4�(=�L������儁T[�<jH��0H1M�"�J�Mw��~�G�D��s�$5?s|�ߒν��V�7����I��/��,�6_�D����`w��K8Ґ1a<�$��	�Y�hQ�o��' �la������a����� ���N�����<��H����f@u��Sr10�}��O������R��6��2㉪�'�&�w�kLm��-��� -{F
��t!���d���-��9� �x�Lĥ��Mrd�CuCD@�_��㺅�%�R��c86|N��^���@�š���e�5/V@E�L��l�!�o��N�(݁�_�ّ�FVO���X�,������d8h��ؼ�~�e��c=o'���Ɛ��voW�C����C"� Q�%j?��I�^&��6V��5w�mǿkø[C�٬o4
��`ב�q
D���>�IG��`y�@4y;
�@���ɦ���٧`��Z�	ϖ�E�ng��o���!��9Abj0��0/�H�e�(�|�yvM�el���1�FX��n���t���b�s0;p�����C�����	���P�`(�h�8znGQ� �4�C���A&�y�À���1�X+YQ�O`y� m+�ho�fTm��h�q`(��P�\��DD�tf�[��:}P�	�)�E���RT^!e���4�B���SK�Gc�EkI��q�ҙl��1pr��^��H-j��F��!�G �\!���P�;_�AS�?�����?���eS�p����H�:��(kX��-�/9��q�L��{����n��!=i9^��5�2e���Lb@KZ/��P���;�����U�֕�lҝX���!�{r� ���ٲ�4q�N;$��g��r���o*�����Ch&o�%l���O����X鱗�<R�3ﱹ�Q!Q���<Fr�x����e�/{D�k�/hjh�t_����C�L���ۿ���>K�7�(F�x�@xw,Y�К�ߧ?]Pp�6(��)��_��Y�7�43�,0H�J�{4Θ3s�C�l&_�Fآ��J��gZ��Wn�Q���1�0��\�_�C���{�Mk�v�oC8�h>C��v�l~׫4��ф ��r�P�h7��R�a��?&�����ըF�RN��-��'����Lm2�;�mB����R�d}K�oz3+D�GnW���d���{�y�b�I3Os�X7��Nn��݄�)3;��`G�w��^=�����(Vɛ����M9*ٽ&S�
!K�߽��<^`�9H	5i8Xe�w0��̄]WN0�_����8�5q�?!8���M^�c+|Y���c���N�w�ʛ���2c�paMꤰ�ĩ0f8F%��u%0�~sh�e�H����R���#�5��Hs��)��/Y�e�?��"��F�Aci���J9 $�{�1��n����{}�4�d} ����Wy�Z���[�"yS�~��oZoY!��"�ko���[;	
((�<��ɂ�=X2���6�\<_	z�Ό��X����m���U�i�p��j��&;���@ ����*C�?��og!W�(��/fP䙨h�tj���`�{R�l��DͶ�z"��&·�@���<���u� XV��H���d���t���ў��h������\�������YrzOנ!s�E���)��A�E}+kG�z�ZﰅTNL0�$!��tc;J��º���٭��VpQ�@�B�3E��5�vj�CY���F�*��[�e�'�?=+@����֮��RG�P���_��z�|��47�2w�%����S�3t�K*u���-1��EEh@��r���Ϊ`�Rl���Ոg�>��a�J=eO�,"Xg8��O���p�]\F>6�i�V�GҲf��9��)�##ǟ� ���Jd>�hpc�$�IJ8sQ�B�v���l�oNM��]��+�8<��ncv���Ƣ� �<Z�D@j-F1��}��ƙ7��Ud��߇8S0���'����`8ch܄����6Rn��6	��O�J�r{XP~!Dv�%�K��o��=m��E�����M�0�DR���U�Ͳ���F]e�r����>��!�b�5uO��Y��_�X�+8�Bg�.�t���jZ�4M�f�W]%�{�	�
�@�Ss=֦s�o�����d�c�2M�Ϳ��w�ֲ5�������+��}q�U]�_0g��,��L(\���k�{w	��L��oj�����TWD/;O��?(�=�Y��I�����J�����W^�T��
�� bp@R�����{ݮ��>[���>2#[�W��U`�e�� ���6S��F�����Zm(3�ݐ)����>-���e��f4
����[��\�}U�{9����tGl��ȕP��宼�/�h���)��x��Z�2K�`�X�u��ժ'��[1��(�K��p��r�g�3��Hw�,�}����CГ�h�����D�Sn��΅ߤ�r��E���������]/�T!9E�iEN����pi�↬���3�E7V������XNO	��]�U�Z���Ɠ[4#��Q�ג��ȵ�r\���z}��2$��<�5�Z�4K���&�}��p�06Cp�*����p�<�R������$�m��c���ݣ��j�-3[\U.�р��$�;軖l��?�^�v�¥rn�=�摿�#�k�C27xZ0��p�a6��x�z�*(��}��b�R0�nI�@��}��r�#�uK��������eR謚�gn�U+�5@Bp�1Ł�zn�H�&םɼ����m����,� Q㡉���:X��
<�{��V�{ؑG�+3I���y�s/"��:��n���/wIy��d��F�x���C�,#_��V*w��h��m���a�j��D!�4��u`JvJq�+,61�O�y9����k�X�-�/�d�hJ��ma�^ǫc�;��}�3�u�.�3�"睃�%�H��灗�z*�q�#��O�����?o`�I'Ԏ��C��حi�	�:$x��W�`�49S��3���!�4'��؜>�  Gr�q��"�Y�P�n<�BIE�xSno)ȟE�����JAL��G
NG�Di�����U_�6�P�]�b*���)�d��=]�]�(ƪm�$��H(�S��!�̈́���7Xt�������>r5~����n(�qB���H��QL�N���?u����*���h�n3o��[ϱ��{��~�1K�Rp^�tY�vө�&˯u�K��a�f~�g���*S�Kp7�rwR'����k3ts~��֓ŕ�"�kM�8!5�0F�k�v=O0,�3��J�q�F
�p2��y�{|��WIA�Nn�|uj!�������<*�h�����w�v�Y��xM�32����<����'�������.��\��?��s��>���Y)�h��}o����϶�=�vBתX�Eb�|B�E	������j�I�&��U�X>�}L�Yk�I����T�ycF"�E@Pg�5�W�)u)��c���U��|BXI�^?��(�g����(�H�V�RS�et"���N�E��H�!:m�O�"�$�M�V>�O[��XI%��*.�>�b$�1��	����eܢ�:� �1�Bv�i)����X�ZQ�י�(U���������bc9M��ԟ�8l���;��4@Kp�w�����%0��yؔ9�v�{{4�}��Zҝ#��9kbh;�2�Օ��a�������Ab���&[v?�������S"�� _�i�ۻ!�>`%۾=�h�$<�����ZS�E	�	;���W��令%��v���t/̉���gn|H|p�<ENUr%�k�V�@)E�#�*J�=����4d�y�%�C1�i�
(0�V����cU#4d"=g�f1���J�9 xOj�Z���۠��j����`��V�N��1�~�y�J���G	�����c� %�\�q�>�y \N	-�_��RW�P��)KV��i�?<���*��w�/ .J���i8�Ȼ��}�i��Y�*6�L!���$�'���<h�Si@GA��\塇*N~��R�J�w��_:�<賉a�|�nQ�ςp2�,;Lܢ��։���{z��
��zyqP���"���*5}����c~�9'�y	:P8܀�g�טL����MÞ-C
��ii$���H>�.e�Zf�)������L&���, 8d3�N���}���x)&�t�|Ra���,��"HYZM�jVmY�w�~��ד�������02�w[O�J"���X�ӑU�:6u��<\D��"Is�!	�6� rc�|qҭzLq ��u��U���l�	\ad���sȆi��'u&R8Uz��}�h�J�D#E��K��Z���8��%��v��H�������r(Ʀc`�ϰ<��x-�Y��	L�o���}t�<OF�?� 6�qX_G/�x�f�U���$Ћ�0I��_9!6�!�