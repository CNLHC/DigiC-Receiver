// ReceiverTopQsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module ReceiverTopQsys (
		input  wire        clk_clk,                           //                         clk.clk
		input  wire        hps_0_f2h_cold_reset_req_reset_n,  //    hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n, //   hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_warm_reset_req_reset_n,  //    hps_0_f2h_warm_reset_req.reset_n
		output wire [14:0] memory_mem_a,                      //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                     //                            .mem_ba
		output wire        memory_mem_ck,                     //                            .mem_ck
		output wire        memory_mem_ck_n,                   //                            .mem_ck_n
		output wire        memory_mem_cke,                    //                            .mem_cke
		output wire        memory_mem_cs_n,                   //                            .mem_cs_n
		output wire        memory_mem_ras_n,                  //                            .mem_ras_n
		output wire        memory_mem_cas_n,                  //                            .mem_cas_n
		output wire        memory_mem_we_n,                   //                            .mem_we_n
		output wire        memory_mem_reset_n,                //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                     //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                    //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                  //                            .mem_dqs_n
		output wire        memory_mem_odt,                    //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                     //                            .mem_dm
		input  wire        memory_oct_rzqin,                  //                            .oct_rzqin
		input  wire [13:0] ofdmadccontrol_external_adc_data,  // ofdmadccontrol_external_adc.data
		input  wire        reset_reset_n                      //                       reset.reset_n
	);

	wire         ofdmsymbolsync_aso_out0_valid;                    // OFDMSymbolSync:aso_out0_valid -> OFDMPrefixWipeer:asi_in0_valid
	wire  [31:0] ofdmsymbolsync_aso_out0_data;                     // OFDMSymbolSync:aso_out0_data -> OFDMPrefixWipeer:asi_in0_data
	wire         ofdmsymbolsync_aso_out0_ready;                    // OFDMPrefixWipeer:asi_in0_ready -> OFDMSymbolSync:aso_out0_ready
	wire         ofdmsymbolsync_aso_out0_startofpacket;            // OFDMSymbolSync:aso_out0_startofpacket -> OFDMPrefixWipeer:asi_in0_startofpacket
	wire         ofdmsymbolsync_aso_out0_endofpacket;              // OFDMSymbolSync:aso_out0_endofpacket -> OFDMPrefixWipeer:asi_in0_endofpacket
	wire         ofdmchannelequalization_aso_out0_valid;           // OFDMChannelEqualization:aso_out0_valid -> QAMDemodulation:asi_in0_valid
	wire  [31:0] ofdmchannelequalization_aso_out0_data;            // OFDMChannelEqualization:aso_out0_data -> QAMDemodulation:asi_in0_data
	wire         ofdmchannelequalization_aso_out0_ready;           // QAMDemodulation:asi_in0_ready -> OFDMChannelEqualization:aso_out0_ready
	wire         ofdmchannelequalization_aso_out0_startofpacket;   // OFDMChannelEqualization:aso_out0_startofpacket -> QAMDemodulation:asi_in0_startofpacket
	wire         ofdmchannelequalization_aso_out0_endofpacket;     // OFDMChannelEqualization:aso_out0_endofpacket -> QAMDemodulation:asi_in0_endofpacket
	wire         pllsampleclock_outclk0_clk;                       // PLLSampleClock:outclk_0 -> [OFDMADCControl:sampling_clk, avalon_st_adapter_001:in_clk_0_clk, dc_fifo_0:in_clk, rst_controller_001:clk, rst_controller_002:clk]
	wire         ofdmsymbolsync_sample_control_pre_sample_control; // OFDMSymbolSync:pre_sampling -> OFDMADCControl:pre_sampling
	wire         ofdmsymbolsync_reset_source_reset;                // OFDMSymbolSync:reset_source_reset_req -> [PLLSampleClock:rst, rst_controller_002:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                  // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                    // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                    // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                   // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                    // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                      // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                  // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                   // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                   // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                   // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                   // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                    // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                  // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                  // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                     // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                   // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                   // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                   // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                  // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                   // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                   // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                    // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                     // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                   // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                  // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_mmbridge_s0_readdata;           // MMBridge:s0_readdata -> mm_interconnect_0:MMBridge_s0_readdata
	wire         mm_interconnect_0_mmbridge_s0_waitrequest;        // MMBridge:s0_waitrequest -> mm_interconnect_0:MMBridge_s0_waitrequest
	wire         mm_interconnect_0_mmbridge_s0_debugaccess;        // mm_interconnect_0:MMBridge_s0_debugaccess -> MMBridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mmbridge_s0_address;            // mm_interconnect_0:MMBridge_s0_address -> MMBridge:s0_address
	wire         mm_interconnect_0_mmbridge_s0_read;               // mm_interconnect_0:MMBridge_s0_read -> MMBridge:s0_read
	wire   [3:0] mm_interconnect_0_mmbridge_s0_byteenable;         // mm_interconnect_0:MMBridge_s0_byteenable -> MMBridge:s0_byteenable
	wire         mm_interconnect_0_mmbridge_s0_readdatavalid;      // MMBridge:s0_readdatavalid -> mm_interconnect_0:MMBridge_s0_readdatavalid
	wire         mm_interconnect_0_mmbridge_s0_write;              // mm_interconnect_0:MMBridge_s0_write -> MMBridge:s0_write
	wire  [31:0] mm_interconnect_0_mmbridge_s0_writedata;          // mm_interconnect_0:MMBridge_s0_writedata -> MMBridge:s0_writedata
	wire   [0:0] mm_interconnect_0_mmbridge_s0_burstcount;         // mm_interconnect_0:MMBridge_s0_burstcount -> MMBridge:s0_burstcount
	wire         mmbridge_m0_waitrequest;                          // mm_interconnect_1:MMBridge_m0_waitrequest -> MMBridge:m0_waitrequest
	wire  [31:0] mmbridge_m0_readdata;                             // mm_interconnect_1:MMBridge_m0_readdata -> MMBridge:m0_readdata
	wire         mmbridge_m0_debugaccess;                          // MMBridge:m0_debugaccess -> mm_interconnect_1:MMBridge_m0_debugaccess
	wire   [9:0] mmbridge_m0_address;                              // MMBridge:m0_address -> mm_interconnect_1:MMBridge_m0_address
	wire         mmbridge_m0_read;                                 // MMBridge:m0_read -> mm_interconnect_1:MMBridge_m0_read
	wire   [3:0] mmbridge_m0_byteenable;                           // MMBridge:m0_byteenable -> mm_interconnect_1:MMBridge_m0_byteenable
	wire         mmbridge_m0_readdatavalid;                        // mm_interconnect_1:MMBridge_m0_readdatavalid -> MMBridge:m0_readdatavalid
	wire  [31:0] mmbridge_m0_writedata;                            // MMBridge:m0_writedata -> mm_interconnect_1:MMBridge_m0_writedata
	wire         mmbridge_m0_write;                                // MMBridge:m0_write -> mm_interconnect_1:MMBridge_m0_write
	wire   [0:0] mmbridge_m0_burstcount;                           // MMBridge:m0_burstcount -> mm_interconnect_1:MMBridge_m0_burstcount
	wire  [31:0] mm_interconnect_1_avalonfifo_out_readdata;        // AvalonFIFO:avalonmm_read_slave_readdata -> mm_interconnect_1:AvalonFIFO_out_readdata
	wire         mm_interconnect_1_avalonfifo_out_waitrequest;     // AvalonFIFO:avalonmm_read_slave_waitrequest -> mm_interconnect_1:AvalonFIFO_out_waitrequest
	wire   [0:0] mm_interconnect_1_avalonfifo_out_address;         // mm_interconnect_1:AvalonFIFO_out_address -> AvalonFIFO:avalonmm_read_slave_address
	wire         mm_interconnect_1_avalonfifo_out_read;            // mm_interconnect_1:AvalonFIFO_out_read -> AvalonFIFO:avalonmm_read_slave_read
	wire  [31:0] hps_0_f2h_irq0_irq;                               // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                               // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         qamdemodulation_aso_out0_valid;                   // QAMDemodulation:aso_out0_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] qamdemodulation_aso_out0_data;                    // QAMDemodulation:aso_out0_data -> avalon_st_adapter:in_0_data
	wire         qamdemodulation_aso_out0_ready;                   // avalon_st_adapter:in_0_ready -> QAMDemodulation:aso_out0_ready
	wire         qamdemodulation_aso_out0_startofpacket;           // QAMDemodulation:aso_out0_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         qamdemodulation_aso_out0_endofpacket;             // QAMDemodulation:aso_out0_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                    // avalon_st_adapter:out_0_valid -> AvalonFIFO:avalonst_sink_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                     // avalon_st_adapter:out_0_data -> AvalonFIFO:avalonst_sink_data
	wire         avalon_st_adapter_out_0_ready;                    // AvalonFIFO:avalonst_sink_ready -> avalon_st_adapter:out_0_ready
	wire   [7:0] avalon_st_adapter_out_0_channel;                  // avalon_st_adapter:out_0_channel -> AvalonFIFO:avalonst_sink_channel
	wire         avalon_st_adapter_out_0_startofpacket;            // avalon_st_adapter:out_0_startofpacket -> AvalonFIFO:avalonst_sink_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;              // avalon_st_adapter:out_0_endofpacket -> AvalonFIFO:avalonst_sink_endofpacket
	wire   [7:0] avalon_st_adapter_out_0_error;                    // avalon_st_adapter:out_0_error -> AvalonFIFO:avalonst_sink_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                    // avalon_st_adapter:out_0_empty -> AvalonFIFO:avalonst_sink_empty
	wire         ofdmadccontrol_aso_out0_valid;                    // OFDMADCControl:aso_out0_valid -> avalon_st_adapter_001:in_0_valid
	wire  [31:0] ofdmadccontrol_aso_out0_data;                     // OFDMADCControl:aso_out0_data -> avalon_st_adapter_001:in_0_data
	wire         ofdmadccontrol_aso_out0_startofpacket;            // OFDMADCControl:aso_out0_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire         ofdmadccontrol_aso_out0_endofpacket;              // OFDMADCControl:aso_out0_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire         ofdmadccontrol_aso_out0_empty;                    // OFDMADCControl:aso_out0_empty -> avalon_st_adapter_001:in_0_empty
	wire         avalon_st_adapter_001_out_0_valid;                // avalon_st_adapter_001:out_0_valid -> dc_fifo_0:in_valid
	wire   [7:0] avalon_st_adapter_001_out_0_data;                 // avalon_st_adapter_001:out_0_data -> dc_fifo_0:in_data
	wire         avalon_st_adapter_001_out_0_ready;                // dc_fifo_0:in_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;        // avalon_st_adapter_001:out_0_startofpacket -> dc_fifo_0:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;          // avalon_st_adapter_001:out_0_endofpacket -> dc_fifo_0:in_endofpacket
	wire         ofdmprefixwipeer_aso_out0_1_valid;                // OFDMPrefixWipeer:aso_out0_valid -> avalon_st_adapter_002:in_0_valid
	wire  [32:0] ofdmprefixwipeer_aso_out0_1_data;                 // OFDMPrefixWipeer:aso_out0_data -> avalon_st_adapter_002:in_0_data
	wire         ofdmprefixwipeer_aso_out0_1_ready;                // avalon_st_adapter_002:in_0_ready -> OFDMPrefixWipeer:aso_out0_ready
	wire         ofdmprefixwipeer_aso_out0_1_startofpacket;        // OFDMPrefixWipeer:aso_out0_startofpacket -> avalon_st_adapter_002:in_0_startofpacket
	wire         ofdmprefixwipeer_aso_out0_1_endofpacket;          // OFDMPrefixWipeer:aso_out0_endofpacket -> avalon_st_adapter_002:in_0_endofpacket
	wire         avalon_st_adapter_002_out_0_valid;                // avalon_st_adapter_002:out_0_valid -> IFFT:sink_valid
	wire  [32:0] avalon_st_adapter_002_out_0_data;                 // avalon_st_adapter_002:out_0_data -> IFFT:sink_data
	wire         avalon_st_adapter_002_out_0_ready;                // IFFT:sink_ready -> avalon_st_adapter_002:out_0_ready
	wire         avalon_st_adapter_002_out_0_startofpacket;        // avalon_st_adapter_002:out_0_startofpacket -> IFFT:sink_sop
	wire         avalon_st_adapter_002_out_0_endofpacket;          // avalon_st_adapter_002:out_0_endofpacket -> IFFT:sink_eop
	wire   [1:0] avalon_st_adapter_002_out_0_error;                // avalon_st_adapter_002:out_0_error -> IFFT:sink_error
	wire         dc_fifo_0_out_valid;                              // dc_fifo_0:out_valid -> avalon_st_adapter_003:in_0_valid
	wire   [7:0] dc_fifo_0_out_data;                               // dc_fifo_0:out_data -> avalon_st_adapter_003:in_0_data
	wire         dc_fifo_0_out_ready;                              // avalon_st_adapter_003:in_0_ready -> dc_fifo_0:out_ready
	wire         dc_fifo_0_out_startofpacket;                      // dc_fifo_0:out_startofpacket -> avalon_st_adapter_003:in_0_startofpacket
	wire         dc_fifo_0_out_endofpacket;                        // dc_fifo_0:out_endofpacket -> avalon_st_adapter_003:in_0_endofpacket
	wire         avalon_st_adapter_003_out_0_valid;                // avalon_st_adapter_003:out_0_valid -> OFDMSymbolSync:asi_in0_valid
	wire  [31:0] avalon_st_adapter_003_out_0_data;                 // avalon_st_adapter_003:out_0_data -> OFDMSymbolSync:asi_in0_data
	wire         avalon_st_adapter_003_out_0_ready;                // OFDMSymbolSync:asi_in0_ready -> avalon_st_adapter_003:out_0_ready
	wire         avalon_st_adapter_003_out_0_startofpacket;        // avalon_st_adapter_003:out_0_startofpacket -> OFDMSymbolSync:asi_in0_startofpacket
	wire         avalon_st_adapter_003_out_0_endofpacket;          // avalon_st_adapter_003:out_0_endofpacket -> OFDMSymbolSync:asi_in0_endofpacket
	wire   [1:0] avalon_st_adapter_003_out_0_empty;                // avalon_st_adapter_003:out_0_empty -> OFDMSymbolSync:asi_in0_empty
	wire         ifft_source_valid;                                // IFFT:source_valid -> avalon_st_adapter_004:in_0_valid
	wire  [37:0] ifft_source_data;                                 // IFFT:source_data -> avalon_st_adapter_004:in_0_data
	wire         ifft_source_ready;                                // avalon_st_adapter_004:in_0_ready -> IFFT:source_ready
	wire         ifft_source_startofpacket;                        // IFFT:source_sop -> avalon_st_adapter_004:in_0_startofpacket
	wire   [1:0] ifft_source_error;                                // IFFT:source_error -> avalon_st_adapter_004:in_0_error
	wire         ifft_source_endofpacket;                          // IFFT:source_eop -> avalon_st_adapter_004:in_0_endofpacket
	wire         avalon_st_adapter_004_out_0_valid;                // avalon_st_adapter_004:out_0_valid -> OFDMChannelEqualization:asi_in0_valid
	wire  [37:0] avalon_st_adapter_004_out_0_data;                 // avalon_st_adapter_004:out_0_data -> OFDMChannelEqualization:asi_in0_data
	wire         avalon_st_adapter_004_out_0_ready;                // OFDMChannelEqualization:asi_in0_ready -> avalon_st_adapter_004:out_0_ready
	wire         avalon_st_adapter_004_out_0_startofpacket;        // avalon_st_adapter_004:out_0_startofpacket -> OFDMChannelEqualization:asi_in0_startofpacket
	wire         avalon_st_adapter_004_out_0_endofpacket;          // avalon_st_adapter_004:out_0_endofpacket -> OFDMChannelEqualization:asi_in0_endofpacket
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [AvalonFIFO:reset_n, IFFT:reset_n, MMBridge:reset, OFDMChannelEqualization:reset_reset, OFDMPrefixWipeer:reset_reset, QAMDemodulation:reset_reset, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, avalon_st_adapter_004:in_rst_0_reset, dc_fifo_0:out_reset_n, mm_interconnect_0:MMBridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:MMBridge_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;               // rst_controller_001:reset_out -> [OFDMADCControl:reset_reset, avalon_st_adapter_001:in_rst_0_reset]
	wire         rst_controller_002_reset_out_reset;               // rst_controller_002:reset_out -> dc_fifo_0:in_reset_n
	wire         rst_controller_003_reset_out_reset;               // rst_controller_003:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                            // hps_0:h2f_rst_n -> rst_controller_003:reset_in0
	wire  [15:0] ifft_source_imag;                                 // port fragment
	wire  [15:0] ifft_source_real;                                 // port fragment
	wire   [5:0] ifft_source_exp;                                  // port fragment

	ReceiverTopQsys_AvalonFIFO avalonfifo (
		.wrclock                         (clk_clk),                                      //   clk_in.clk
		.reset_n                         (~rst_controller_reset_out_reset),              // reset_in.reset_n
		.avalonst_sink_valid             (avalon_st_adapter_out_0_valid),                //       in.valid
		.avalonst_sink_data              (avalon_st_adapter_out_0_data),                 //         .data
		.avalonst_sink_channel           (avalon_st_adapter_out_0_channel),              //         .channel
		.avalonst_sink_error             (avalon_st_adapter_out_0_error),                //         .error
		.avalonst_sink_startofpacket     (avalon_st_adapter_out_0_startofpacket),        //         .startofpacket
		.avalonst_sink_endofpacket       (avalon_st_adapter_out_0_endofpacket),          //         .endofpacket
		.avalonst_sink_empty             (avalon_st_adapter_out_0_empty),                //         .empty
		.avalonst_sink_ready             (avalon_st_adapter_out_0_ready),                //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_1_avalonfifo_out_readdata),    //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_1_avalonfifo_out_read),        //         .read
		.avalonmm_read_slave_address     (mm_interconnect_1_avalonfifo_out_address),     //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_1_avalonfifo_out_waitrequest), //         .waitrequest
		.wrclk_control_slave_address     (),                                             //   in_csr.address
		.wrclk_control_slave_read        (),                                             //         .read
		.wrclk_control_slave_writedata   (),                                             //         .writedata
		.wrclk_control_slave_write       (),                                             //         .write
		.wrclk_control_slave_readdata    (),                                             //         .readdata
		.wrclk_control_slave_irq         ()                                              //   in_irq.irq
	);

	ReceiverTopQsys_IFFT ifft (
		.clk          (clk_clk),                                   //    clk.clk
		.reset_n      (~rst_controller_reset_out_reset),           //    rst.reset_n
		.sink_valid   (avalon_st_adapter_002_out_0_valid),         //   sink.valid
		.sink_ready   (avalon_st_adapter_002_out_0_ready),         //       .ready
		.sink_error   (avalon_st_adapter_002_out_0_error),         //       .error
		.sink_sop     (avalon_st_adapter_002_out_0_startofpacket), //       .startofpacket
		.sink_eop     (avalon_st_adapter_002_out_0_endofpacket),   //       .endofpacket
		.sink_real    (avalon_st_adapter_002_out_0_data[32:17]),   //       .data
		.sink_imag    (avalon_st_adapter_002_out_0_data[16:1]),    //       .data
		.inverse      (avalon_st_adapter_002_out_0_data[0]),       //       .data
		.source_valid (ifft_source_valid),                         // source.valid
		.source_ready (ifft_source_ready),                         //       .ready
		.source_error (ifft_source_error),                         //       .error
		.source_sop   (ifft_source_startofpacket),                 //       .startofpacket
		.source_eop   (ifft_source_endofpacket),                   //       .endofpacket
		.source_real  (ifft_source_real[15:0]),                    //       .data
		.source_imag  (ifft_source_imag[15:0]),                    //       .data
		.source_exp   (ifft_source_exp[5:0])                       //       .data
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mmbridge (
		.clk              (clk_clk),                                     //   clk.clk
		.reset            (rst_controller_reset_out_reset),              // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mmbridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mmbridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mmbridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mmbridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mmbridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mmbridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mmbridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mmbridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mmbridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mmbridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mmbridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mmbridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mmbridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mmbridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mmbridge_m0_writedata),                       //      .writedata
		.m0_address       (mmbridge_m0_address),                         //      .address
		.m0_write         (mmbridge_m0_write),                           //      .write
		.m0_read          (mmbridge_m0_read),                            //      .read
		.m0_byteenable    (mmbridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mmbridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                            // (terminated)
		.m0_response      (2'b00)                                        // (terminated)
	);

	OFDM_ADC_Control ofdmadccontrol (
		.aso_out0_data          (ofdmadccontrol_aso_out0_data),                     //       aso_out0.data
		.aso_out0_valid         (ofdmadccontrol_aso_out0_valid),                    //               .valid
		.aso_out0_endofpacket   (ofdmadccontrol_aso_out0_endofpacket),              //               .endofpacket
		.aso_out0_startofpacket (ofdmadccontrol_aso_out0_startofpacket),            //               .startofpacket
		.aso_out0_empty         (ofdmadccontrol_aso_out0_empty),                    //               .empty
		.reset_reset            (rst_controller_001_reset_out_reset),               //          reset.reset
		.sampling_clk           (pllsampleclock_outclk0_clk),                       //        clock_1.clk
		.pre_sampling           (ofdmsymbolsync_sample_control_pre_sample_control), // sample_control.pre_sample_control
		.adc_data               (ofdmadccontrol_external_adc_data)                  //   external_adc.data
	);

	OFDM_Channel_Equalization ofdmchannelequalization (
		.aso_out0_data          (ofdmchannelequalization_aso_out0_data),          // aso_out0.data
		.aso_out0_ready         (ofdmchannelequalization_aso_out0_ready),         //         .ready
		.aso_out0_valid         (ofdmchannelequalization_aso_out0_valid),         //         .valid
		.aso_out0_endofpacket   (ofdmchannelequalization_aso_out0_endofpacket),   //         .endofpacket
		.aso_out0_startofpacket (ofdmchannelequalization_aso_out0_startofpacket), //         .startofpacket
		.clock_clk              (clk_clk),                                        //    clock.clk
		.reset_reset            (rst_controller_reset_out_reset),                 //    reset.reset
		.asi_in0_data           (avalon_st_adapter_004_out_0_data),               //  asi_in0.data
		.asi_in0_ready          (avalon_st_adapter_004_out_0_ready),              //         .ready
		.asi_in0_valid          (avalon_st_adapter_004_out_0_valid),              //         .valid
		.asi_in0_endofpacket    (avalon_st_adapter_004_out_0_endofpacket),        //         .endofpacket
		.asi_in0_startofpacket  (avalon_st_adapter_004_out_0_startofpacket)       //         .startofpacket
	);

	OFDM_Prefix_Wipe ofdmprefixwipeer (
		.asi_in0_data           (ofdmsymbolsync_aso_out0_data),              //    asi_in0.data
		.asi_in0_ready          (ofdmsymbolsync_aso_out0_ready),             //           .ready
		.asi_in0_valid          (ofdmsymbolsync_aso_out0_valid),             //           .valid
		.asi_in0_endofpacket    (ofdmsymbolsync_aso_out0_endofpacket),       //           .endofpacket
		.asi_in0_startofpacket  (ofdmsymbolsync_aso_out0_startofpacket),     //           .startofpacket
		.clock_clk              (clk_clk),                                   //      clock.clk
		.reset_reset            (rst_controller_reset_out_reset),            //      reset.reset
		.aso_out0_data          (ofdmprefixwipeer_aso_out0_1_data),          // aso_out0_1.data
		.aso_out0_ready         (ofdmprefixwipeer_aso_out0_1_ready),         //           .ready
		.aso_out0_valid         (ofdmprefixwipeer_aso_out0_1_valid),         //           .valid
		.aso_out0_startofpacket (ofdmprefixwipeer_aso_out0_1_startofpacket), //           .startofpacket
		.aso_out0_endofpacket   (ofdmprefixwipeer_aso_out0_1_endofpacket)    //           .endofpacket
	);

	OFDM_Symbol_Sync ofdmsymbolsync (
		.reset_source_reset_req (ofdmsymbolsync_reset_source_reset),                //   reset_source.reset
		.clock_clk              (clk_clk),                                          //          clock.clk
		.aso_out0_data          (ofdmsymbolsync_aso_out0_data),                     //       aso_out0.data
		.aso_out0_ready         (ofdmsymbolsync_aso_out0_ready),                    //               .ready
		.aso_out0_valid         (ofdmsymbolsync_aso_out0_valid),                    //               .valid
		.aso_out0_endofpacket   (ofdmsymbolsync_aso_out0_endofpacket),              //               .endofpacket
		.aso_out0_startofpacket (ofdmsymbolsync_aso_out0_startofpacket),            //               .startofpacket
		.asi_in0_data           (avalon_st_adapter_003_out_0_data),                 //       asi_in_0.data
		.asi_in0_ready          (avalon_st_adapter_003_out_0_ready),                //               .ready
		.asi_in0_valid          (avalon_st_adapter_003_out_0_valid),                //               .valid
		.asi_in0_endofpacket    (avalon_st_adapter_003_out_0_endofpacket),          //               .endofpacket
		.asi_in0_startofpacket  (avalon_st_adapter_003_out_0_startofpacket),        //               .startofpacket
		.asi_in0_empty          (avalon_st_adapter_003_out_0_empty),                //               .empty
		.pre_sampling           (ofdmsymbolsync_sample_control_pre_sample_control)  // sample_control.pre_sample_control
	);

	ReceiverTopQsys_PLLSampleClock pllsampleclock (
		.refclk   (clk_clk),                           //  refclk.clk
		.rst      (ofdmsymbolsync_reset_source_reset), //   reset.reset
		.outclk_0 (pllsampleclock_outclk0_clk),        // outclk0.clk
		.locked   ()                                   //  locked.export
	);

	QAM_Demodulation qamdemodulation (
		.asi_in0_data           (ofdmchannelequalization_aso_out0_data),          //  asi_in0.data
		.asi_in0_ready          (ofdmchannelequalization_aso_out0_ready),         //         .ready
		.asi_in0_valid          (ofdmchannelequalization_aso_out0_valid),         //         .valid
		.asi_in0_endofpacket    (ofdmchannelequalization_aso_out0_endofpacket),   //         .endofpacket
		.asi_in0_startofpacket  (ofdmchannelequalization_aso_out0_startofpacket), //         .startofpacket
		.clock_clk              (clk_clk),                                        //    clock.clk
		.reset_reset            (rst_controller_reset_out_reset),                 //    reset.reset
		.aso_out0_data          (qamdemodulation_aso_out0_data),                  // aso_out0.data
		.aso_out0_ready         (qamdemodulation_aso_out0_ready),                 //         .ready
		.aso_out0_valid         (qamdemodulation_aso_out0_valid),                 //         .valid
		.aso_out0_endofpacket   (qamdemodulation_aso_out0_endofpacket),           //         .endofpacket
		.aso_out0_startofpacket (qamdemodulation_aso_out0_startofpacket)          //         .startofpacket
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (16),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (1),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dc_fifo_0 (
		.in_clk            (pllsampleclock_outclk0_clk),                //        in_clk.clk
		.in_reset_n        (~rst_controller_002_reset_out_reset),       //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                                   //       out_clk.clk
		.out_reset_n       (~rst_controller_reset_out_reset),           // out_clk_reset.reset_n
		.in_data           (avalon_st_adapter_001_out_0_data),          //            in.data
		.in_valid          (avalon_st_adapter_001_out_0_valid),         //              .valid
		.in_ready          (avalon_st_adapter_001_out_0_ready),         //              .ready
		.in_startofpacket  (avalon_st_adapter_001_out_0_startofpacket), //              .startofpacket
		.in_endofpacket    (avalon_st_adapter_001_out_0_endofpacket),   //              .endofpacket
		.out_data          (dc_fifo_0_out_data),                        //           out.data
		.out_valid         (dc_fifo_0_out_valid),                       //              .valid
		.out_ready         (dc_fifo_0_out_ready),                       //              .ready
		.out_startofpacket (dc_fifo_0_out_startofpacket),               //              .startofpacket
		.out_endofpacket   (dc_fifo_0_out_endofpacket),                 //              .endofpacket
		.in_csr_address    (1'b0),                                      //   (terminated)
		.in_csr_read       (1'b0),                                      //   (terminated)
		.in_csr_write      (1'b0),                                      //   (terminated)
		.in_csr_readdata   (),                                          //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),      //   (terminated)
		.out_csr_address   (1'b0),                                      //   (terminated)
		.out_csr_read      (1'b0),                                      //   (terminated)
		.out_csr_write     (1'b0),                                      //   (terminated)
		.out_csr_readdata  (),                                          //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000),      //   (terminated)
		.in_empty          (1'b0),                                      //   (terminated)
		.out_empty         (),                                          //   (terminated)
		.in_error          (1'b0),                                      //   (terminated)
		.out_error         (),                                          //   (terminated)
		.in_channel        (1'b0),                                      //   (terminated)
		.out_channel       (),                                          //   (terminated)
		.space_avail_data  ()                                           //   (terminated)
	);

	ReceiverTopQsys_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),  //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n), // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),  //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (),                                  //   f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                      //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                     //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                     //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                   //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                    //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                   //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                  //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                  //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                   //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                     //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                    //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                  //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                    //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                     //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                  //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (),                                  //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (),                                  //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (),                                  //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (),                                  //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (),                                  //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (),                                  //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (),                                  //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (),                                  //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (),                                  //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (),                                  //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (),                                  //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (),                                  //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (),                                  //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (),                                  //                    .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (),                                  //                    .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (),                                  //                    .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (),                                  //                    .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (),                                  //                    .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (),                                  //                    .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (),                                  //                    .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (),                                  //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (),                                  //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (),                                  //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (),                                  //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (),                                  //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (),                                  //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (),                                  //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (),                                  //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (),                                  //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (),                                  //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (),                                  //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (),                                  //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (),                                  //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (),                                  //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (),                                  //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (),                                  //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (),                                  //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (),                                  //                    .hps_io_usb1_inst_NXT
		.h2f_rst_n                (hps_0_h2f_reset_reset),             //           h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                           //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (),                                  //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (),                                  //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (),                                  //                    .waitrequest
		.f2h_sdram0_READDATA      (),                                  //                    .readdata
		.f2h_sdram0_READDATAVALID (),                                  //                    .readdatavalid
		.f2h_sdram0_READ          (),                                  //                    .read
		.f2h_sdram0_WRITEDATA     (),                                  //                    .writedata
		.f2h_sdram0_BYTEENABLE    (),                                  //                    .byteenable
		.f2h_sdram0_WRITE         (),                                  //                    .write
		.h2f_axi_clk              (clk_clk),                           //       h2f_axi_clock.clk
		.h2f_AWID                 (),                                  //      h2f_axi_master.awid
		.h2f_AWADDR               (),                                  //                    .awaddr
		.h2f_AWLEN                (),                                  //                    .awlen
		.h2f_AWSIZE               (),                                  //                    .awsize
		.h2f_AWBURST              (),                                  //                    .awburst
		.h2f_AWLOCK               (),                                  //                    .awlock
		.h2f_AWCACHE              (),                                  //                    .awcache
		.h2f_AWPROT               (),                                  //                    .awprot
		.h2f_AWVALID              (),                                  //                    .awvalid
		.h2f_AWREADY              (),                                  //                    .awready
		.h2f_WID                  (),                                  //                    .wid
		.h2f_WDATA                (),                                  //                    .wdata
		.h2f_WSTRB                (),                                  //                    .wstrb
		.h2f_WLAST                (),                                  //                    .wlast
		.h2f_WVALID               (),                                  //                    .wvalid
		.h2f_WREADY               (),                                  //                    .wready
		.h2f_BID                  (),                                  //                    .bid
		.h2f_BRESP                (),                                  //                    .bresp
		.h2f_BVALID               (),                                  //                    .bvalid
		.h2f_BREADY               (),                                  //                    .bready
		.h2f_ARID                 (),                                  //                    .arid
		.h2f_ARADDR               (),                                  //                    .araddr
		.h2f_ARLEN                (),                                  //                    .arlen
		.h2f_ARSIZE               (),                                  //                    .arsize
		.h2f_ARBURST              (),                                  //                    .arburst
		.h2f_ARLOCK               (),                                  //                    .arlock
		.h2f_ARCACHE              (),                                  //                    .arcache
		.h2f_ARPROT               (),                                  //                    .arprot
		.h2f_ARVALID              (),                                  //                    .arvalid
		.h2f_ARREADY              (),                                  //                    .arready
		.h2f_RID                  (),                                  //                    .rid
		.h2f_RDATA                (),                                  //                    .rdata
		.h2f_RRESP                (),                                  //                    .rresp
		.h2f_RLAST                (),                                  //                    .rlast
		.h2f_RVALID               (),                                  //                    .rvalid
		.h2f_RREADY               (),                                  //                    .rready
		.f2h_axi_clk              (clk_clk),                           //       f2h_axi_clock.clk
		.f2h_AWID                 (),                                  //       f2h_axi_slave.awid
		.f2h_AWADDR               (),                                  //                    .awaddr
		.f2h_AWLEN                (),                                  //                    .awlen
		.f2h_AWSIZE               (),                                  //                    .awsize
		.f2h_AWBURST              (),                                  //                    .awburst
		.f2h_AWLOCK               (),                                  //                    .awlock
		.f2h_AWCACHE              (),                                  //                    .awcache
		.f2h_AWPROT               (),                                  //                    .awprot
		.f2h_AWVALID              (),                                  //                    .awvalid
		.f2h_AWREADY              (),                                  //                    .awready
		.f2h_AWUSER               (),                                  //                    .awuser
		.f2h_WID                  (),                                  //                    .wid
		.f2h_WDATA                (),                                  //                    .wdata
		.f2h_WSTRB                (),                                  //                    .wstrb
		.f2h_WLAST                (),                                  //                    .wlast
		.f2h_WVALID               (),                                  //                    .wvalid
		.f2h_WREADY               (),                                  //                    .wready
		.f2h_BID                  (),                                  //                    .bid
		.f2h_BRESP                (),                                  //                    .bresp
		.f2h_BVALID               (),                                  //                    .bvalid
		.f2h_BREADY               (),                                  //                    .bready
		.f2h_ARID                 (),                                  //                    .arid
		.f2h_ARADDR               (),                                  //                    .araddr
		.f2h_ARLEN                (),                                  //                    .arlen
		.f2h_ARSIZE               (),                                  //                    .arsize
		.f2h_ARBURST              (),                                  //                    .arburst
		.f2h_ARLOCK               (),                                  //                    .arlock
		.f2h_ARCACHE              (),                                  //                    .arcache
		.f2h_ARPROT               (),                                  //                    .arprot
		.f2h_ARVALID              (),                                  //                    .arvalid
		.f2h_ARREADY              (),                                  //                    .arready
		.f2h_ARUSER               (),                                  //                    .aruser
		.f2h_RID                  (),                                  //                    .rid
		.f2h_RDATA                (),                                  //                    .rdata
		.f2h_RRESP                (),                                  //                    .rresp
		.f2h_RLAST                (),                                  //                    .rlast
		.f2h_RVALID               (),                                  //                    .rvalid
		.f2h_RREADY               (),                                  //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                           //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),      //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),    //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),     //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),    //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),   //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),    //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),   //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),    //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),   //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),   //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),       //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),     //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),     //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),     //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),    //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),    //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),       //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),     //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),    //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),    //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),      //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),    //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),     //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),    //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),   //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),    //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),   //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),    //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),   //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),   //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),       //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),     //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),     //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),     //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),    //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),    //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                 //            f2h_irq1.irq
	);

	ReceiverTopQsys_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),              //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),               //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),              //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),             //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),              //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),             //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),              //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),             //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),             //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                 //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),               //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),               //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),               //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),              //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),              //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                 //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),               //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),              //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),              //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),              //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),               //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),              //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),             //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),              //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),             //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),              //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),             //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),             //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                 //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),               //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),               //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),               //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),              //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),              //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                     //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),          // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.MMBridge_reset_reset_bridge_in_reset_reset                          (rst_controller_reset_out_reset),              //                          MMBridge_reset_reset_bridge_in_reset.reset
		.MMBridge_s0_address                                                 (mm_interconnect_0_mmbridge_s0_address),       //                                                   MMBridge_s0.address
		.MMBridge_s0_write                                                   (mm_interconnect_0_mmbridge_s0_write),         //                                                              .write
		.MMBridge_s0_read                                                    (mm_interconnect_0_mmbridge_s0_read),          //                                                              .read
		.MMBridge_s0_readdata                                                (mm_interconnect_0_mmbridge_s0_readdata),      //                                                              .readdata
		.MMBridge_s0_writedata                                               (mm_interconnect_0_mmbridge_s0_writedata),     //                                                              .writedata
		.MMBridge_s0_burstcount                                              (mm_interconnect_0_mmbridge_s0_burstcount),    //                                                              .burstcount
		.MMBridge_s0_byteenable                                              (mm_interconnect_0_mmbridge_s0_byteenable),    //                                                              .byteenable
		.MMBridge_s0_readdatavalid                                           (mm_interconnect_0_mmbridge_s0_readdatavalid), //                                                              .readdatavalid
		.MMBridge_s0_waitrequest                                             (mm_interconnect_0_mmbridge_s0_waitrequest),   //                                                              .waitrequest
		.MMBridge_s0_debugaccess                                             (mm_interconnect_0_mmbridge_s0_debugaccess)    //                                                              .debugaccess
	);

	ReceiverTopQsys_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                              (clk_clk),                                      //                            clk_0_clk.clk
		.MMBridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),               // MMBridge_reset_reset_bridge_in_reset.reset
		.MMBridge_m0_address                        (mmbridge_m0_address),                          //                          MMBridge_m0.address
		.MMBridge_m0_waitrequest                    (mmbridge_m0_waitrequest),                      //                                     .waitrequest
		.MMBridge_m0_burstcount                     (mmbridge_m0_burstcount),                       //                                     .burstcount
		.MMBridge_m0_byteenable                     (mmbridge_m0_byteenable),                       //                                     .byteenable
		.MMBridge_m0_read                           (mmbridge_m0_read),                             //                                     .read
		.MMBridge_m0_readdata                       (mmbridge_m0_readdata),                         //                                     .readdata
		.MMBridge_m0_readdatavalid                  (mmbridge_m0_readdatavalid),                    //                                     .readdatavalid
		.MMBridge_m0_write                          (mmbridge_m0_write),                            //                                     .write
		.MMBridge_m0_writedata                      (mmbridge_m0_writedata),                        //                                     .writedata
		.MMBridge_m0_debugaccess                    (mmbridge_m0_debugaccess),                      //                                     .debugaccess
		.AvalonFIFO_out_address                     (mm_interconnect_1_avalonfifo_out_address),     //                       AvalonFIFO_out.address
		.AvalonFIFO_out_read                        (mm_interconnect_1_avalonfifo_out_read),        //                                     .read
		.AvalonFIFO_out_readdata                    (mm_interconnect_1_avalonfifo_out_readdata),    //                                     .readdata
		.AvalonFIFO_out_waitrequest                 (mm_interconnect_1_avalonfifo_out_waitrequest)  //                                     .waitrequest
	);

	ReceiverTopQsys_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	ReceiverTopQsys_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	ReceiverTopQsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (8),
		.outErrorWidth   (8),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),         // in_rst_0.reset
		.in_0_data           (qamdemodulation_aso_out0_data),          //     in_0.data
		.in_0_valid          (qamdemodulation_aso_out0_valid),         //         .valid
		.in_0_ready          (qamdemodulation_aso_out0_ready),         //         .ready
		.in_0_startofpacket  (qamdemodulation_aso_out0_startofpacket), //         .startofpacket
		.in_0_endofpacket    (qamdemodulation_aso_out0_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),           //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),          //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),          //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),    //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),          //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error),          //         .error
		.out_0_channel       (avalon_st_adapter_out_0_channel)         //         .channel
	);

	ReceiverTopQsys_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (0),
		.inReadyLatency  (0),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (pllsampleclock_outclk0_clk),                // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (ofdmadccontrol_aso_out0_data),              //     in_0.data
		.in_0_valid          (ofdmadccontrol_aso_out0_valid),             //         .valid
		.in_0_startofpacket  (ofdmadccontrol_aso_out0_startofpacket),     //         .startofpacket
		.in_0_endofpacket    (ofdmadccontrol_aso_out0_endofpacket),       //         .endofpacket
		.in_0_empty          (ofdmadccontrol_aso_out0_empty),             //         .empty
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket)    //         .endofpacket
	);

	ReceiverTopQsys_avalon_st_adapter_002 #(
		.inBitsPerSymbol (33),
		.inUsePackets    (1),
		.inDataWidth     (33),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (33),
		.outChannelWidth (0),
		.outErrorWidth   (2),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_002 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ofdmprefixwipeer_aso_out0_1_data),          //     in_0.data
		.in_0_valid          (ofdmprefixwipeer_aso_out0_1_valid),         //         .valid
		.in_0_ready          (ofdmprefixwipeer_aso_out0_1_ready),         //         .ready
		.in_0_startofpacket  (ofdmprefixwipeer_aso_out0_1_startofpacket), //         .startofpacket
		.in_0_endofpacket    (ofdmprefixwipeer_aso_out0_1_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_002_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_002_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_002_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_002_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),   //         .endofpacket
		.out_0_error         (avalon_st_adapter_002_out_0_error)          //         .error
	);

	ReceiverTopQsys_avalon_st_adapter_003 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_003 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (dc_fifo_0_out_data),                        //     in_0.data
		.in_0_valid          (dc_fifo_0_out_valid),                       //         .valid
		.in_0_ready          (dc_fifo_0_out_ready),                       //         .ready
		.in_0_startofpacket  (dc_fifo_0_out_startofpacket),               //         .startofpacket
		.in_0_endofpacket    (dc_fifo_0_out_endofpacket),                 //         .endofpacket
		.out_0_data          (avalon_st_adapter_003_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_003_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_003_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_003_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_003_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_003_out_0_empty)          //         .empty
	);

	ReceiverTopQsys_avalon_st_adapter_004 #(
		.inBitsPerSymbol (38),
		.inUsePackets    (1),
		.inDataWidth     (38),
		.inChannelWidth  (0),
		.inErrorWidth    (2),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (38),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_004 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ifft_source_data),                          //     in_0.data
		.in_0_valid          (ifft_source_valid),                         //         .valid
		.in_0_ready          (ifft_source_ready),                         //         .ready
		.in_0_startofpacket  (ifft_source_startofpacket),                 //         .startofpacket
		.in_0_endofpacket    (ifft_source_endofpacket),                   //         .endofpacket
		.in_0_error          (ifft_source_error),                         //         .error
		.out_0_data          (avalon_st_adapter_004_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_004_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_004_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_004_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_004_out_0_endofpacket)    //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pllsampleclock_outclk0_clk),         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (ofdmsymbolsync_reset_source_reset),  // reset_in0.reset
		.clk            (pllsampleclock_outclk0_clk),         //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign ifft_source_data = { ifft_source_real[15:0], ifft_source_imag[15:0], ifft_source_exp[5:0] };

endmodule
