��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���5p����O+��l,�m�}xP�C�W)��Tv��ܣ%W�	�Om#�<�i�3K?E(ڟ��̔O�7�w�&ף�ߍzq�Y��q�S��#��!�|KN��텢^p�4�|@A�^�۩�3���4�
M�c��DoƦ�4cJOvKo�A�{!u�{?�Z����	ןw��4�l��y{��=��thї�8��E���؁?�	t�#���U�?Q2	��M���B4������z���A�j�eU�s�;&���4 �PV�1i3�r�ˌib�;���m���R"fg�mZ�K�,t�0k��G�|�r�΢�*{5��'�~(��6n��k�hVۗ�wՄ0-��-s6� �d�����4�_�b�v�년f���B������h��Q�L���Y��s���fP��@z@�X� NO5��d��r��v�xG�ϐ��2�B���11�.��eڭt\}�����/��o22T��%��P���1�1tϑMass�*��~� v 	q��3>\�����K>o���Y_�;�t>���!�^��:���@m����	-7��XxA7�z����m^�����O>mŒ"N1���-�!iSl������z�0�![P�y����+��&��R=�����ua0]p���}�>!)h�K����)}���h$'�8�R�	����Y���OG��J��Iz�xo�6���^���P国�|�r26w)g��J`jf�qH���>h���>�K�pY.��7OR�g�w���I��yE��cn8i����� ����w��J�mp�ɪ�7�~�::ĉ�����!��)V�b�ܞ���7�� Ô>��=�>����6+�Z��}M�9⑷5�
	ٔ/���`7����Y
k˚!�. ^;����M�A���O-�4����ݾ��|��E[3�T8hS���C�!��ʡ�*b�Ai0��J|��0CfX�Z��}���v���VMSI6�p�	ҥ%����͝�{Π�+S�����|�K���@o�������sA�A;:Q�cg9u�!�f{T�Z���X�������&ߤֆ�*t�Zب�'$~�}=��ֱ�����
�~��C;��.`��U��0�L黀M��(~�� x�/z��zo�N󀽍{�XWk�`L��&�%�h� ��y���*�WWS�6Bݙr.��ÁQ����mP-�Ms��}��D�j�st'�-�Sen��
+>�y��ɛ��EGa���,��V*׉Y�'�,PJ]���<?�2����gI\)�>Z��Ţ��`���Ӥ��u�?I�:c��[�RW��?'��jG#����T�����bii��&,��@��o�%UƓ_�a�&3�A�218���`｟���qO�O�,��!��U�Z �n�=�@Wj >ѸQ��)(��/�?ʻ~�����ˉ�/z�h�֏ }�3��W=�����9���N��>b�#J�@�[���\q��,����d��w-�.�����/���+Z%VB^��,l���y�����I����x�s����R _��sf�y�U2�̇��=����G�,|�4!l�a���,Z����
�P�[a�=��A�N_��!<�a��ul=\�Dw!�_����w�2R
�@�P���2�_i�� 0� �=�\>��j��x��*�@�^V��_o�NjD>�N�h�ִ<`}�?O��b���`L$u���C	����\��K�eU@�]��+���j9�/ϩw+q��AG������=5��{)�~��'�
�ڒ�Jޡ7~v9ج�(}��cV9~^_#�������mR�ÛD� ��:}���Iy��}8ܾ8`�w��&��8~f�y@f9���ݞB\�tk6�ћ�^�ˎ��|�O��lK�C�C6킞�Yz� �~�K4���&x����ߩ���ʜ���*E2��.Y˓���29%�NE�g�1�`K:@��_��>'uks;V/�@��[����6����N����������&TQ:E��p�J8� \aW0�:%h��-lԑ�if!���<u��!p�7+m�!?��NgT7z䪇%L5�1z�����-����[�D����n�`��5���}�]�D��S����Gm���I��2r������@�̯q_��_����l�'	z5��1��c�E�S��C/�y���uܥMߍ&>ץ��c��
`ͨ����TE��-r/�b�~�ƕ�WD2�s��e�C��Lfg����]Ğ���5�躋�:�~�
���s/�(�t����f}U�'�Q�.��K�Q�?;���i�x��_4ȏ�z�v�
�"A3U�m@sb��b�m�rB���\��©/���r�Y���mey2-���K����fx�4��=��?p��#���n��ڋ�ܠwϛ���"�y_�S��J{=���"CӀH��>!�,e���1i��j�AdN'���u��5+˫�Cc��>��!�r^\j&6vq�h�{!"��̱$����<�_�����V$.+@���1V0ߔ͑Ϲ˄�r
$�z��tM���֎��%_H	��>�P����KBK-Y���2��z�_�f2��<0o�o'�&��O�g�x����]���/���&�?�]m�;m2���&��)eh�3O��B�^7�(H /����ېD�K�."�0�8���2���c�p���ƈ<�-�fu�!Г�����\䊐�LF8��{j�6q���{���;-$C����Z{b��4�����8�� r7R�B�<���n���բv�k�'
�%�M��LB{���G_��ὧ����+Iy82�*W���}��D
Ɇ�����2�7ʑ�
�.�l�n��L�KQ�+4Hi1��gad��k�kR��H��?%|q�	�-ǅH;���j�У��� �����rVo�[��c��6H�M�YMJL^��E����3�+iɁ���j��:A� pn�N{���u\��W;��_Al hZ/���	��b}���	;^�2 �H�8��K[���G@�ԫ�&'�y3�O������N'�2�ֺ����0�T* �u6j_�8�0��{[̳������G���G�si6���`�QlGG�B��-�&d�TCVB�i������\:>�i�U/{��9%�u?4�/ϔN�2��a�B3:��A�R���b*����,��yQkp�S��u���O#��B���9K謎�}7�ZB��v�If��Ɨ$*Jz/������w�wS�m�^uEw҆u�%�zQ�=k|�}D��: e��H�Ϫ���A$�D��dь�v ��?�q2M��,ALV�?`�e$����z+S]�h)4�ފE<��_
/�F�b�S-.{�����C^.@���p �
�Ļ,)�K�@w>���6����N���4�.'8��J�����ն�p�aAC�ԻP�w�#r��S�a)�C���9�nJB'�M���!ϕNru=� ��-����@/)x���y�T��s���<5�s����E6��1} ���%��~a�m�)sGߊ�.�7�� �6��b %��M���8ˡ�-�6�;k�?�̈́ɹ��D@����09���ĸ�S�p�x7�5Mv�&6���l��=6k�6ѫ4ܟV
��Qo���X���𤮕�q{��V�B[�@w���~����cHr��8u�������;���q;y�C���e��{��G��ձ�0�RXO�nk���H� 3� ����o���=���-�-����;�ˊ�� B��iͲ��YDřSX�k�޳6(��R�z%�[�dj*Y��N���m��v�/���@��ȳ�۠UaE1'��L(�`ט6g�h��E��A�/�+X�W�a.ü^�J�9=�mV��W8�L�����a�{�s�D�u���0b4����b��B|S��$V�\�ˤM��NY���x��G�斦����&���Y=&���7��.�[{���w>e*s�~y���%�W�Ů���{�:O4z��q�rJ�:����{��5\���vL�U,�yu���)~��%o&?���L��M^�u���r�7]�=8�����t'>dX��w�
y�Y�;�.oPM�?R��$��8��h2����~,=���$rXO�D�A�C/�:)7���Q*ح.��&O�P�KOq��}���'.XO�:�s��fX풹��
���t�K��k�c
�nhD�Ugޚ]�R,��Y��Q�݇�����L�%yK�b|C�lY�셕U�?hϴ��B�/�d��a��
@N.�4�+�I7�u;^G���H)z���w::϶A���lg�U� _��x�#�	D%٣�y<�����'�\[��~J�d�'@�l5�XZ��C������Ƒ\h���$v��zA�5t�,b���{|�e�����8"g� �ɡV��l���'[�*�GR���)"����/���JQQ��\���4�t)*I��=��������[��E	�_Ƞȗ�M�@�vBZ����׭� �!�k��"�>��^�[���Zn���4����&ߛ��I�i�b��&�R�#G��15�`�=:T��_릜�hC�R�Rx�ei�֩�4�G G��x3�.^�W����=���C�"�s�H�&O�H+�1s��6���2.:N5{�ݩ�Tn#��ud����ϒ�o}KtJ���>����qwQ#�LQ�������K%�tck%���_'�N�[fq��� �Qin����c|�8�d���j�f0v�f��خxmT�Vnv�)��yja��AL�;��cB[�t�����Q��Ǹ����18�U�js2�m�q蘕�����=�3���t��5�V�\zV"~��N2^� �l͟UY'ZP��(9�^�ڰ��z��r��j�Â�7jZA�_�^�{���2��w� Ԥl�>��	�Y�v(� 5J+#ӎ��J����� ��s�tE�X[aQ�/ZT!<��Q!�7���' �0;�A�P�RdQu��������G0��x�+e�l�U(��X�����k�)i:��9����1�x.�+�>��Vr � ���eE �7��sx����)s(Ť���Si�XѨ_�[1�$�G OYkT�0�2T���]����^�Θ�4H�Z8����nX�vD��4�gu��ɀ�U��Q���#`z�劉e��'y�
���`vd�Ů#QhN-��ҵ�I(	����\��c��G����8��K����_�*̲����(T	b�87��r� �3�C��һ��`��G�!�p>�H�N���` C�NOuOK%$V��/��͞�5w�s��AY]���H�������Zm$�֦�R&M@�`!I�L�UO,Z�^�<�T���y�ͭ=b����M�Ѷ�K�c@t�Z�>++N�f;޽�qsP!W��B���}մ�o �0��"{�����E�&?,6�A���#�
�aq�c(K��t��B��>����k�A`Hl��0-�lq�#��=����I��H����KxDFm����Ds9���	�����tĲ5�|�v ��aM�?Z7��1�z�(���
��� �d�0M�e�@t�����NYN{����kd����3@��k������=�#E˭�I��t���
2n�S:�u���2Z���)����'�n�zIŕ^����i@B#M@��Sc]�����u�zR���X�i%+�v-���:�e�$�F��l,��j�ޡc���e��D��+>m��$G^R4P�O�	��4�/k�.�����\�!�{`�ԥ��-g���%��Ic��V���u��BL~�^���S@2�(��ɽ*C��w�A	{]
�{R�c�av J{��cc���$6��e�f����-�%��,m7��_�_uN$݇ӎeUo4�3W�\k�{�C{<BJ~,d\��Q�����̮Ht�T:]"<g��8�D&ᜂ�dr(�F	�6\DťO!��"�h��v5��؉h�<Ҩ��q%"�N�,r�3Rl�m~M�q:z㊔A���7G��OV��=m��Xo� ��m8�jb0e`��NB���a���˒��L5��I2���a(���?���d������Y�Ga�m�4�tZڨC�r��f��q~.&�i׹y���#Duj���ts����b��{2�IØU���X�����W	�%Ӱyc�pou,�,�[z��!^\&w9y��kk�EV�6َ���A�j%YF�% �@ӻ�����n�f*>}��*��lr�7gVْ�N��6I�#U�?09��W��x�s�'�a7�A�*�\��� c�5�~L�({�1KV�!��;"E��Ap�R�d��+��vf�y��W�?x!���qE�uwj=��:S���՗W�P]w����/��7(j�.Zo�ƕ�$����b�6���ރ-q:��l�OwT8&���7P�a�Q}[��˝_;#B���Vjx�i�175E����˓�����	e㔾�М
69�Ή�h]\"��F��
��s��p����f�Q��"��$4O��z�N�<E;�������~J1�x={�HB�J0���L��C����|��L�~�5(���,�跰��[�ʋ����X����N]��V��%la�$�a�	�:�� Fh�����e�k����K�,�M�� �G��� �)��}٤pm���:�J� ��M�.����,�Z�$�;W�����Mq�����(�bS��ʕ�Y��D����wb��8�l�Qq�M���\�ٰZ8�tnLM4�J`5�3��J.���m�~ֹ��#v��GX!��WU�-0��GSVX�E��iO�3�p,�\�7�oc��A�,p]A~n����5k��:L�c�B�&����ǚ�_��ُ2����zw�{���5��v�������J�:j��q�`m1�6*$�l���̆����WxI�l��l�����u�$pLě�L���z��$f�b�Y�y�Ŕ��C����@bQ��R*@e��W�k�\3h���*��hWoF��;tE|�+N���Y��[���u��k����+�mg�/Z\#��>N��^s<�\Y\5��]���^�s��4*3�<`�����+����޻n~�{ctHLe1vC��z#�X���wfJ�"b�~��o��R�7 �W��0l���ܒ�sYy�x��=���� E��B�5SB��J���-�v�`U�-WE�ɷ���a���Q�þ8i
bfB�0G�8'�?t�XT��u�S�T�� l!,J��>�)z��.lYoaHb��u���n�! _��ϜE�J�D�m�����?��}�o����>���?�-�aO,/5y���:���嚟���^�H]��%��/p�!V�-8?��J45�#���gaD���N'�dq%-)�​�,���o���w�{`Rm|�Dh��*��׼���n�lp$96ws�FiJy��A8���8m5ee-aq3�?@��ka��kR��&^��g��i^_�j���֙7T��Վ��}������^���><�*��+����䉛F��}n=��E��^q"��x˧W�	���]���Q�9�r�_�BN�QŐ��t},�3��oZ��S�-®ţ���uf��@���5E��9�����yh
�F��2����Nv�s�?i2���	"�c(
�U��O���mf��΃BB�Sv�΍��
�g?��eA�Mc�48��x�m	u9�U�U�y��<�r�Sb�iq`gQl��|��W��nC[eB�:��y���d0Lي�rO�.�;�p�N��QLҋ(�`�������� �d�h���!���Q�����0_OY���j�&�>��ر-g����eQCn9п��#���A ��":�}�I�L�J�����a���\x3�Gt^���i�kG�-�G&����U�Sv��e�P&C[g�ǗQ#��U����`X��EA_+�'Fe�%�i����$������wנ?��m���g�[*\NS��%�������E��@�f���H\/�p�!�R�o�۰	;o�A��5\��ܡ��Ӫ��dmҔ�����
�\���Q,�?��7�)�I�@�w�