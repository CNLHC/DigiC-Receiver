��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�@��x��QZH!/h�0��i'�M*bH�	��#��V:�b�dR�\YŢHq�ث�gHgG��N�6��&Tz �J�t�����13��T�>P�w��b ������o��γ�y�;�����;�A��ćV˴��1�"�8��u�K^���V>��
N\��Xy\5��=N�{Ώ[r(73F:���+��G�>�cFt�t{�
詢:�>��u>!:��k�e��w�@���&�(�^�i����'�-q�v[�,���تxr�}�+�T����G���k�d��;+6a�^��t���j0u�Ŋ@��qc� Ȧk�Ƴ��><!�\�Җ�����Y �`UmA�D�3�Ȍ������;�jeW�,�8�i��//�T�}�)?���W?Dd5y���i��7y�����H-N��Ű�/�4.�¾�V��®��,4�0ťU*�;������V�#���[�S�aJ�aǙ(l�nT*],�AihF�~����^Z��Jk��1#.i�#ܵ�;��o~�o�vҽpss����8qu�)m>I)���$���-���t7�_�qK�ݵח��1��<|i������@�����V�0_��*��m����b�IvS�C��=Ll�}i��֪T��G�=���A�!�#��^�C�*���0p>Ť5|�e�ԐQ��;��N2�Fk&jG�K���7Q��B���D��chV`[�z9�W���[�y�i�6.j,�`"�Ǌp.N�j�|�����|K�O,�=nT�8἖�O45}�E��3<�����/��Kj�M>9�O ����KW
Pn�#٦�΍�21�5�ɾB�c|�7�+�!��z�=�'�#�jT��6�^E�.GS�F��.R4�Ô�ibW���.C���ɦ�������>3 ��ǎh^�9���E��$n%����=��*L <}M�[���J�$q3�k<��%o���n��?���ev���	
P�z�����l�ࡵ&�^�t���M���'�kS��!�C�c�hp�.
��S��q+�)�I�I���%omR������E�a�"�����b��+Ĳɇ2�A��(��5B�ʶ��[}�(�� ���ɚ����w��Q�I��)R��_7���r_�ټ%�d�_�w���G�x�B���="��+�E�,��<4���(
�@�E��=��L�{��f�1�����s��@�������k�z�e�rA�����Qԛd)� ���.qX7h.��7Z�-9u�'��ot�w�i�*(;}�׼�L'�����9��8s�u%�f����9���ѝ��r{�G�/	fsW� �g�*zi��\�������3F��{g#AFE��H.����_��*p��R�$!.�X���l��@�UQd=Y�v`�q1J��cMD��|�g�m���T�_]���&�ǋ@!�ͳY=<c�!Q���=-W�K��T_`�>W��[!G��H�d�4g\��7t\�'�U�*���Z���o?Ԁ�o��Qa�����8�c�Ơ��J�'i���u�ؑ�����B���A@4C�e�DZ�PXD��M�B�t�e�M��|L��\ ��@��h.q���D�ʹ)��iw�� B���wu}�Nja�����o���
;x��.��Q�"�k}� 5>X��L����m��R*7�����~y[�6�?W)nυ��0�W�r]F����3v�����ʛ�U,˻{�D�1�/m�L���&�ů}E��bUQ��$���8� GЁ�<���ҽ�����a�5(��4f|�Kx�c���:��@���aG��kW���n�y3 G�ӮwK�o�[WX�D�-6��� ����I�5z��c?�*p_�Q�9����Fe�
�y�L�|R�· ��R�ʓ��]U�9�d��Gp�I�!x�)�R`���w��ѓY�����!ew7i6�<ۧO!�:�=[��JR�u��z�'Xu�l-N}j2�W�����g�_��V�#,�ʫឺ��oG�8��`����� �9�C�P�h?��|2���h�t5��
ܸ&��i>����<�����/�O&n0��E�����M�������3����mh�Wf8���N}ua��٧[{y�Zu��%3cp�(	)}�ca#־x?���㘇֜��菥����Њ#�6/4%td	,��B��c�?�oZ��|I{�h%���m��=����@z�6�5�&�����rP��kf `d���,'�֫�&v�1�<��Fj!oY�U�p����Ir�������iA?GsH�p+�3�����/oz[���*))szr:|�-�|�r���Od�dEpZ��՟�k�Q�����<`+��w@c��U�@Mi�+O.����n#��w�@Z
�^��s+�6F`��<��i(-�Y��9��he��43�M��U̔��E����Y����;�O�M����Ǟ��4;������~o��*��q� 
��`�W�����֤ef==��Ms�zC���}]���TR��`���:�~�P؄�}�݈V���Cay H8b��*oS|��Ư�i�0��j�X�������G<'��н��x9�����m�Gs�=��DUvA�b0�ĵ�����Y�M�J0g�,s3���=�҅{��7��z��XdD�����Y�@M �M�	헲�6�^��R�%�j�t �|)v:d�D����nӱ�� >�*�M���(� v�tM�+��WNπC�PA8T�%c4ϢWt�/2�\�tK t(ނ
�6�
�yi(l~Z�|uF�K@=Tv �۰!2�� 5���%K]�W�c��&�GKs�j��S�~f�RL��ғE J��br8YE�H��\�&���=e�P�5����D�w�G��$����>1JU��Z�o����i��v��R򹕟�>P78KVtYg�T4s@���T����g���� ��8s����O� ���.$z�.�U��xMF������ܴ�5;Q9׀�n�/j�{@R�P���%L��'l��J��Y��&�y9C���
�A����ǌ�� ,U�(�v[Y���ݷ��,��X����Be�FU�Q$�S��\m�+ό�2�v^�Α{[UL�T
`l~�.��jtB�UAB�|a@��g>��h�'2�Fs)
��n�x)�H�����5���d�/?>�G^r|��v��=6*5�,,��=����
X������_�����J޴bu:�L|}����P����M0U
E�"��w��|�� 3�Q)k���fj���k9���F�O�j5'�qI ���`Q��+�z����\�tn��U������8����X�b��Jj?���vf�0:h,��eX`{�F|�<���T�6;T1�8���r�����!���K+tb�"����ǝ�sC�AZ��XTU8(iU)'K\�j��$2?'N�yMA�0�� v�����O���CDa���V�@@�� ���K�YWY��Wh���/E\L���Ǯ�n� ���'��ab���S���'����*�%�.�"����=N�T�
�P���P�#�DU|�]���C� 2|�urmRit��Q�I�K�����I.��o��/x�����^��X_X;ߜ��cg!V�9����C�Py�>���+/�m*fy�ĳ�w�_{CS�k�B������f�ā���ǘ��v
k[�ݔ��Bh}�m�L!���dm%�辪<�ޝ�h�h�@��%o��Ϫ����ZW>�� �
:�OV��R��o#��`��A��g�,��yNub?r��2;㷩�F�&&rE�#�<�=Ա�?\xێ�`N�P_�Ld�C]�5G`�?_�]#�.Ё#f[h�c��U��zZ����P~D���co�)�4�c1���8�|w"��$l��RS�)�E��߷�m�E�hV.�"'l/v����pd2���7q�D��9j"a	\u`��wp���s:�C��H[)Ă���A�.I�\;E�G��@I Cx�MU�<u��0,a�^�Y�/ŋ��6$F�-��� Hfz`I�7��\8d���5���(�꠮�R*]�0����=�؎�Jѕ����C��~�bDi�� '�BT�� H���8����ϪU��O9j~=� 3
�h�9o4��r�å$�D;+��T��K�cڈ�U:��!
H�d�$�J�L۠�&�dl�'��|G��&�&ʓ0��'���I��O���SG��_�h2�3�  �>	�˔O�?{x$��K7IC��UR2&Ȃ�+���#�ǣ�v0c��M/�3u�M�5�b��r��h)�^]�I��N�J*���w��[�\m��Q�o�o�.Z֑�^ըR����x^]�ڛ7��`��#�rK1��d�[f*�1~�e&�C{��Su�v���QM�}���j�G�a9�$����j10Dq���˲PPA:������풵_�l$�έ�-e��jI��GD���j�I���ܒ��t�d�~���:o�r4O)�ϩs�|�5�}{�p���YE3��H��jޔ��}7,x2�p'Rx��f9���Ow�}!����<��L,��_}e ~'�/\�f�$�i�0iX�Or����}-���������E��]0&5=FK]r�;qw~ ��T�H?��ؐ��s�Ŕ�bb?x�����VP�Ā���F�'=��hD���|�ٴZI�cwȂ�f���܇7�O���	�i�Sc���AM�ً0-���Eʃeb�L
4�`�K
)Y��)u_·�I����;�3ޒ��[/<«-�>;T���`:C c$�������g/pK�i���m���o�D���̐k����S�fy
u���s��vP�磲�X��I���!����g.,��4
3�\7�Y�0��W_~���"��*�n�Ҳh̓����=86ZĜ��X�s{�'�.'�G�v^�pJv��VH��7���"c�	Y���C,6N�G�`~F��`5m�NA4�j^�p�R�(�uS 3�ڙy��ݖ��!����ZM��б� MÝ��,�v�/*���աgp/��H��T��vQ�h?A;������{�L�V��Jl�(��S?� ��I�أ+�&P��{�0� �����ű�m�������ݦR�G�4m��;�V���\m?�\]!Jqx�~`\Q"�2,*%�Q�1�AI� e�����6 M�s��Yp�%.��y�����h��[?>K�`(�w��ؘ-.���U�R���f���E�O����H���dR�l�p��`?�)����4���,�G��jry�3���L7k�=M�r�����@ةwD^�0��m���1��"ى5����+Yg����eV�s�d��b�HA���_�c��'�w���L
�ѵ��_��5M%��8x�,
�O	/��Y��u�|'��/n� ��ᨸh( 	`� _�͋��LQ
�	.�0��O;�,FIŒ��E�a��3�e�* �q�Lg�&{g�}�ǽT��Ʉu����wi���Nv���_��������9Ez���h��\͘���K�����p��:1̃TYome�[�hn�;�l}�(����;"� ��lbjT�!�J��H��Ȩ���)#P���*{��Q�	6��+��t(cTv��<�7|F�A�B�x��R�3H�I·V�����z�1yU�Hkʠ"�BЊ[�U����L�h.8�4
i[�m���J�ύ0�#yn���Fua��n
��30�3RC��G7��{r(��b��y. ��:<�5�;�O��!N��v*J�*A����м�P`E��^�m�]�g��yD�X�i��%��&7I@�>+o]�*����Ys.	UC��)<��kP4	�#�	���8;�ݭ�o�;0�!����ݞ���5HU�m�_�2f\����BQ�<�k��7�z�oq�x��I�-�+ PeЇ��	��fr$��9Y�r+̸X;}eiq<�ӸW�}7Br�g5H�=��L����BcI�eTⷍE5�z�]�-�����
��O�A����� \��
��뫓�{�`�*��dFD���M�h���ݏ�(���H(e���#��r/;��D䊩#+qi�V\��ƭ���
�����i$bŤ?`,~��$T�\�5�e`ԛx��v�.������|g�G�Q�^.=��Q^�qOI��ݣ;"��k��hč��d��'kp�� 9S�?�-�QE��#][QG�����	��CJ�K^�к���((���5L�,����.���6;)�Rm`k��b�X��1`�^�����W��� 8:���譑��Z��c�^:������f��.XnAP�6
�"�Y/ �w7�U�jJJ��J�˂����M�^��Z0�߆����6�=r�\O�`����t����9|Q`�1q��5:ش��x)TI��W�{��@��P�5�~`����HP8�t�WǼ%cH�R]���lq��6b�DJ$�|ь	"�/�[S�+�j@�y���I���>
�Z����#KĆ$� � x�w^�������	pv�N6�����΂ۏ_d�G-�Eᔂe�5��r�s�0��6f}��k�f���'��!����Kt\�f��!���Դ�7��vI���ķ���q�h$�@��H�?�(;[��bs���G�M	ٹ��U!&e�aʃU��B���$yu� u����짤��ܒ�L�(�(��?����@a����lf�&�Б����nnA��FZ2�ƫ���-����_��D���:Ǖ��T;&��⾸nĦ�"�N��H��5HH��]��
��A|�n�T�/���u�z��x���lE2q6sM�b���cI:���s{SJ&���� }��c t��6�_�eO���p��g�z��^�9���I��% � �8C�1��0j9k �6�\$���=�`��RlƼ�U#OX�m�_l<k�9
�}6̩#��wԟ��툿�7$dU��ig��mYK$L��}�{y/�W����W�Q��v�Dл�+��><��Sw~��-N�cD9��@��%�v��\0sWV�A��j���c���.;���ǌPMy��N]֔�ibSKt���@��QaLT�٫;EM��{�[� ��ƕ�Z�)]�}>3�1T(w��	*�9�/"XDB��+�����F�y� �!y}��0�b��T!�e}��N��_�_�2!pf�P�/��k{�t��۸�nÜ�MP���ҟxdl�+X�c*a�UC�Ե����ey}�點F_0����Z�X
���z['�:���;' ��R���[��Hx�ϛ�6*H�=SZn���7�<zt`���i�z���y���g#��F��N�O#�&CR��YӤ�{�L�����i=h����&����n h�G�և�!M�4`�%�6n�Ѓ���oԍ��ɚ�$@�����ޙY>p`0���.���=.Aݎ�?%p�Z��{��x	���(Bv��s`��+���i�8�K:k�\O���:B�L�����}����c~)w�Z�YU�`��J�Q������z鎑�a�mr�.)�y1)�6P��ߡ��F1��g��D��J8m���.��!����ءs�O��;�[��HpFk�46�����pr6���[�$�ڋ9u�.�&�e� �Ag�8C�b扭##�Z�����8�ۄ{j�����/HE	��R��?���#�a�I�%�Q�'u��Ôĳ�Wu=� ����������ޕc�a�T������{P���(:�7A��m��O�;X��w�� �p'4~�D)U,�������s	�[�C}����}�NS��tN��|p�;wa<\T{M����8��x���.� �хU1r�҂�jVq��|,�Oߦ�5���U�%������ղ���C�L��������T�:�أtQ_=��ݿ�!��.mLV��p�T�^��y�;�D�wز�ﻮ��ڌ�������4�a��Q��,�!�.����J�xY�����[��Ƶ�01&��'3CPu ^#�*��sV��E�u�::�1Ѯ�)|r'e���6�\����1C�'r`�0O	�$À�x�[�ڟ�Od�����Q,\����j-�u�0�W���n�d��%��jr�-�9,��3.��⌮�^��-Tu��.�S�cN& x1�#h�S�w��yO��q��Jܫq֨W���덤��-�U�I���}.lX����O1��Z�x�찄�O���Z�b��@���#���l��4�?�lmM��]�Fb�h�1�8 ���7M:7!�A)hM�h��ŏj,T��$<a,l�O9�H=u��ˌ$8��r� �$_%[�8J3Jt� {�h�V=�P<z�m�|!���&�O�e���f��i+��|*M�����b#��P�0���V�k��z�32f�g	Ix���[�*����A��'5�ף��/i����U&�Q�P�԰��cDfx]廷c�Q��z̘�y:,�c�D�E�~�j|e�!����=���ީ��ȅ���mrtޫɢ	�#�hޤ�)>Q�
3Z�}1�[�5�J/�3rK`��3�/��/=T�ms\�)oYIsO w�0��MPo��vK��SZ�X��K�g%lg����?R�P`����i$�����;0.^[XSA���N�CS���05�2X:���u>���%�0�~�xo��pX���c�C�rKw����&�p/��)rL��D���pw�[Te]ޡ��:sB�0û9��a�����nw�oJ���x�coDxn�N��t.X~Zr=mA�0�����#~ؙ�9�$�=��~8^&���r��H�\�t�l�����,1��>ͮ�7��GX�:uz���u�+�n�5q\�Ct�E�Y�J��p}W���:���~ �ha�"F|ye˨d�t,��z�(.�&`L��O-M�)���%�^V�S���%�G�Oә�.�Z{qp�fX�C�KTs|�6�L�<�
q�ULm5�i
���k���T�d�ِ�@3�u� n���eЮ4�e��xS$P�m�^��ۿ��$�ٷ�Ok���*�!�*�EK��G�vA������<H\�Py�?k��q��P���At�N�Uv:��Ӆ3Ч�]n �O`S�B�ޡ'2	��!�K�xQg�nˤ�Ҏ���Pj�/��أ�L������"P(�
Ѩ=�86�4�7x���TB����}�Ύ7�Rp0��"
q�fư��>ڴI���j���!:N��\�Lrj��(j�1����^lѼA�/��!�I�Ud��^Od��*�y(�@�9��]U%`�.��`fL�"(MG�[<�4wRK�wW��:��:�2�%7�����x�!���z��?�D>R
���}���3�A��[�VJ�Jƅ,`�\�Ԁ3����j��U৆5�O`��¸.\�s��?��y�c�ѕ�����ۘJ��΋$8���*��/
���Aߦ�pk'�W�YP0�u�D|~���uJg���L-�ť7j�A�h�6���F�n7Qc�E�>Y�3����<%�\B��2У5��Ͽ���`2Z	{A͟�x��x��+Z��}�\E��@BVX8	 ,�`�����E�.?�
���x��u�Q�,�L%������|Ra��EJ�ŰU�&rł^�wN��������ogO���Ԍ�5oq��񔺳������h�yz�*�㍵v?}|��[������/u�q|����P3S�*���R�����]�3�>m���=<(1M-�����aV�DRu7�q+�g��T�u?�} ���;���Y@�^�a�_]�!Hk��ƌt����5ƽGnv��r�/�6��������"2��O����'=bW��j�y�YϠ_0�*�Y?.�K�b����1B�����þ=ͷ���\�Fm[�
L��Z����<��Rhl��Җ����	"˽���F�V��bIF�
!�wdE��"P��VS���j@NgO�1��Ի�s+�_�02��a�U�-Wk�@N��q��2uμ�2 XG0߂)Ґ�}�di� ��֒���$
� ?3$x�cS"j��W\p�9��c<,9�k��M��6=��p�RS�Nj󃭍��ݲv4�c�3'bٮ�?�/0���*�gY�^��ή�Wof�gW ���GΊ.�[��������s�iZ waS͊��zbγ��%�|	���/���S^�P�|��<������1�\�#Qx?�RM�o5�0��B{ƿ�x[�/�i���1�G"�����a��?��4�~р8��xչ,�@�r���@UX���m�`�Nv���%��]��ޠ��^�~]��(<s˖��n������M���kw���r��fg�@���)�%��Ǒ#b� �=��;�:���C��w�˴8v�τʙw�U��m
����(�:������\��VDܿ�^��w��9 #��Ρ��wsP�C��u��UԷ�(��	�5JWl�A�sF�d�^�k]���u��Tg�;O�é]��0*��`��9��!���kXo�XQ	��r��G92�w9�h����K�
m���'��O�	�<&��A�������-g�ƽ̊Ƙ8{��u(�a�C/�
dy�lt���qŶ1�BP!h���mIG��Y8fU��,�"0�u}�^�X@�\`������>�k�2t[�L����/����Ǝsf6	5e^x@Mt��"y�zJk帻�R�0�-<�=���m�4����_�3�q4B5�ꗣj�8��ч�E��n�&E�t��c�Ԏ�o����+����c��6M�X��r�� TϵN�w�kmo�Q`�]���J^�`X-�l����6�2
�����Y��mO%kN����K9�Ѳx{��>�~�3˩��%�g*x�=�Cy׮��ý����������N�T���Ւ�Po��L�V������\���_��ѕi��(��&���!!�k��P��hx�Oz7���o5p��I��-lS��� �:����f/��3�C��^���l�i���P�wD�-�� d�'3k@Sȇ��K'efϧ߹����B̄���)�+��EZ���ʭ�{ԲR󻇦�>�I`��u������4X�tbVͭ��`,r��$q-}!�d=,ET�V#�����a׾#���B�B}�D�>�֦0x��W�s�\W��/�5OP`���z�{F1��y�{#�.�-�\�Q��v������7�$N#�R��2�2�6埔,b�Е|E��2�)��k�ӷ*�q��2��{m����aY��E����w�������yk1�RsH��㖊�`$dV��+�)"}{AV�b?����;�e�L	��G�;S�j��N��5��񶏵�uj�XcD�S�L��%ң^�d �T��o�������3f�%�^�
�7p�T���,�$��IZH�V��E�.)��zI������vc���c�y1$���4�5�	���_�R5��8�a����=�0E�yp��GP�t��$0���9�0.������i%e�	����5�\C�����CQ��2]�8�����"92�9	��7L/����H�y� r�_J x���jv��v����&�~�����s͑�X��I6�����`����g0T�(X��Pq3�-�[R�%xYm	O7c9�ky��Rf�f %6�t�e����X� 9��|�c[=����.��Zz�r��p�X��
.���4�N��bh�rYC�MH{�|`2�H		p�Ҳi��< |(���%��3����-c
+�y5��QDfH�8ů1��Q#���8��a�g�W���϶�K�ɷ��܎-4��zy|���<|,���!��~�:uK2m�蘣��f�a��(T��������3���DǊԃ�綵N��6k�J�������X=��0 le�s	�;�4�躒q,.G�Y�� |q0��Wl�R? ��D�!��^V5�@ηd��~�6;�; �7��R=X��Q"Y�g�^6�p��=�aԹMET}Op���[�J��f���DCQݓ���<�����>:\'�a�J��2��2t�)�e�_���Ss�[5�ս��y��'����~T�+{��~��P=�0�kq+�}��Ff
ʲj�`�2��~o���r]�������2�-X�H��`�G���/�$DL���zny����lX�D!��Wy�/�t�9���k�^� AZ�{�c�(��v�vm��0V��jdѻ���!��u��ɞ�N�[�t�$�^��_��b���*��K-�|^�JG�x�y����k���N$���u��>%?�O�Uo�;�eoi���h��	��4�10^.'F1k5�8���<��I �=��mC�V�lp�>�1Kx~�Uh+������ŀ�@�,�I|����U�����PnC�����9�� z�:_� �"��δ
�$+�N�Gt%���H�d[x�]�����F�X��ru�E�<p�SV�� k��&˹(�/x��:2w2�����Q|�Ò�f�(-(��F���~>���4�!!�ňy�L��;���@]/�䤜i�)��������{��U�������՛�r޲��vb���ɺ�Kg�s*�%'N,�	�#�o;]]H��:�^�M;r�������)��Y��k���w�E���ӑ>c�B��X^����2�Hxvf����.����"�6�M����:r#]�����p�m�rt�PP}�5���ڦ�������M!��(֟gA7��&$ۆ�$3j�L���+������/���X�¡@@Kvۀ�lf)���l�gNr�VUýW�'�$�^-$��6�u��I	�l�����a�=NkX^�%��i!S��-LFM�B��]*��`v�I0��9ظc���Q��yM��ߏm+�lr��ep]֩UHq$h�:���m�W�s�e�Ӽ�-h�b#�t��Pj�I� ��T2�,�oOک�h�����yϽ]�!ywSHB(άڄ�l��j�\0����{��z�ݜq����ڦ#^n��:\� z�>��5�
��<,'!�̆��9DD���ذ�G4��e��Y�f�N!&��j�[Q��=�	����ͬޒ"��c���.������{[��L�����P�<	��a�ܷ��'�u@-��wq�{��r\�E�����!<��9�Ŏ�ɵE�Nٍo��6��X�n�+ ��߀E@Z���rh�P׽�� yJ�����&1��)�7�h +#���b�m�]�fSIUe��b�x5O*�~C�l4G��-�/�D?��O�L����@���Vv@�Z�������\X.Ε��4;��RM��e3uqL�<���n�)lrRRI߸m�Ӈ�U�Pi��s���Xz}]�%06�m�:v'O1r!ݟ	s�Q�ü_^)E$�n+CZ��E闱^�\�5@�:S�?�Z۠5���*�;f�E���wň+�O*w*H�=Z?��Q�G����٭Z�;��O I��G�:��Y�����D@9��};��@�f����ld�f� �ȁxE�z�W�90��@�1C�oS�R�����W�r;5O�;�Qp{�G>p!T܂��Y�j�*
Y:˘���"��!�Gi�7"]����X�Asu����z���c��1��!a^g�W�q>�v��G�
�k]��J?q�ǖ��F�F�<A��{��G�!�����``�J�\=Et�����3������$KiJ�C����jm����`���.sϩy��:U�B���f:�R�ϬQ !�Ɲ#�v�0�M��e�a"��)�G�L8+pgB���Z�8j���֨{��#���0ȴ�xIr^�`�毘�;1��m
���F�7i=9ϡڑ�̏�O�_k���5ȡ�6`�t�ԋ6���C�[�Wɠ��!U�J�,��d�
���Lo�{w��:����:1�x�ӭ����1�aH����csP�o>��a�%��?%M�[���򓟇&�*	�Id�'�hpVC`�|�*4�T�|���G��S=x����k�%�r��㹄���׆^͙l��� 'j���*_.�]�Hg0�uӕ��
V���y����H��?���/�[Ec�R�aF��{8~1�'�F]�E*�R���#�b3�x�4��]�
��5o���bd<�om����)ݝ#gl�Ǆ�<�P�ga�P��Ў:,IM.N*;	j��I�i� /y���f�nC��NY���1���7��W�v��up�t�x�Y��uy��z�����]���f}Hɬ^�������+��&Y�3�e��������'����� >=�#&�ǝU��!��~R~����-�q�<_��2���˹	
�)����=�\���79wؿ2��!��H�}`�Xpz�r��'.IlT��$H�ȋ1��=u�<�����պE��p�C`�A�	di���us�&���]��K��sw�BG��{y&�EXB.�U���*���ѡI �z��iW���Sy�6��l��Q�@iz�v����	:��z3�j���������<g�=y��$r���w0"a�W5@�[ύ�$�_$G��Ë��th�\���ڍ���/k<�y��If��w�Eg�m��z��u�p�-'3_�n�yݣ*����@,~�K�S>���
�����9@Q2���}T��TX6�èG)�P������@��P���Y��i����R@N3V)��z��^�����&�Rh7����E`{,vk���d����@l��)�sT�E�#!RMj�S��j{f�;(PFLׅ7�NVE�ŌX�a4�d�������@�F�k�4�(jUI��W�v��&�Q)�[�+�>?�]P`g���D�؝�AA��)��04"�E��=�|�ܞ���a���=<��l6�9�x��M�;p�7qHDE��[������X��l[4Y�kQ���S����.���":��o"AZ�~�c�~H��SUS��M�RHi�9���k���ST�vuj�~�`����H�NUG{�+K�<���ܴ{���z�~[�����\U��E�Ჱ��'e=�1���}���j��VY��7��X���p��K[��g�v z"+�_�CW��p�g1�T�b>~
�S�K�p��<LoZ�%����y~&�}N�)�痞�i���ox�؃��r`�#��u�a6I{c���7�0��"�K��'�JF�o�h�5e->�Hs��C�ʜ��}kOW�4*�G���r�B���	��M9;��ZC�"?��/��@�|į �|H�yA$�� GuؑB{V�M���?������p�X�Z��6�i/VX���J����2�%u7%N�Z]}�U��%y��C��H;>���2c[��`��A[�r5���"�{-�[���WiI�qD�	�>s�d��*���s���\@�} ��k���1�Y�C~c�J֪׼M�h��2����u��F�hL�G��l�� ������ #+�؏Is�%�g�HkOM�{d�����K6PO ��Ǔ�Q#8/ߍ��/�"��em����vD�j��-����h�"�XdL��!l&(�uy����B-����xK�ǆ�4~�ʊ�gK�Q�'QH�_�%�:1`�H���/z��2,
��H� 2�����ѩ�ArL{Y�l8��������)�V{4��b,踫!�]��A.�P��"JL &�D���るLy,�U?I�̺jߪ���A�Y{\�Zm�u	B�Ҳ��6b-�WdF��pϗ���D��S�o�c"�""ɃO�*��~{Xp�����SܚJG�2����q��Kq��U�Ha$M��Va$W~�!��%>��]�ss����(�6�-,;+�`s��ŀx�K��NL��C�N/�~��@�i}
B��&�j8L�)6�� v?�y����Tt�{g�a_ʵ�/���V�g�|��$�(�I������q��'�vױ������5-���7�=�r��+X"�)"���<½i�qJ���n)e�ǒb�)�!]�ʎ��e)g���)�픚��T��Ɵr��B�~<��.dX���YȰ����g�s�_Ͽ�"��U�P5�מI�Ay�_��oCF�{�'X�aٖFU@��y�~�p�~��+��14JP�X���R �,��q�\��n*=ZkL4YlF�iĴ����ܯ�ڍ��DM��H7��U��1ByA�����q�L�L=V���nX��AI���]Ҡ��v�D�}�.#ς�Ӹ��& �0ԑt��,0�"02�n���g���)+8��?��2B�<Oy! �l6�
*�v����τa�ah�\f-u��c3Ff��/�#�x,G��_��w�_ܝ�Q�'�*n8��]`��ʩc%�DFq��i&�	���4-��&xϟ璔�4ͥ��}ĹF$�[ZS,l�9�/|G���k����#ۡ�m^��&&�!Z:���tewQs�'t�
� �GXHZ�eI��05��m�xy�F�9�J	���
�V�R�Th!��톚��:3	�m�\��t�Cb�!�Me��&v,Ke�đR�+|�_?�\�7����~�
�Lg^�&�2v[u�fN�tQE�Xn���8��j�V$�k��7��S�|��Uу�=���u3�z8z��-���k�Y|����Q��}K��u�H�P�Ť��̱�/P,�^��9���ϊ�,������(v�HJ�W�*Z�w���~�������Ey����2����������^����$Ո�d�er�����3>�U���=G܎��9:"��5i���	��˪���@��O�Т ��V򗙮R]�E������GM��O�C���0_G��z��`B [���f˙���F�V�5��)9×�s*�����L\ڪ�#��dxɤ��$���&\2:�Jr�� ո^��s�K��T�i'
NW_z�^hW�E��ھPHk>���ɲ*Ư8�6Q�n�3��Z몽ȼ��א�th���T��(J�V��-ދ�-̐�����P��Z��F��Ʀo̾�WC*�#�/D�m��>����O&߂O����兹�����.�RL-W�$d]6b)������ϕ�$J�f�q݉V�4B��.UI~x~7[A�8ty)�G�)XF7µم�6�~�0򧴋:	�� ��u�l%���T�?�؈��cMM'�1~.�&jB��DQ���̡,K!��"$%5��&E\B�
�Mx��6L/��eH�.G�Fi�a �<왧U����aj<<�<L��L�ސkCg�I2=<:���*�d��V����E����z�[��A=�n��hf����<�ūq{ig�d��P��'���_��p1_@������X1";m��l��(���w����C�
��'�`ę����lk��%IG�Y��5�t �QH�j���!��b�cFB�'��r#�����s�2_�*���5����(8�8�7����sWiar�Ȇ*��9�Y� ��:̨���7�����_!��\�w}:�J��o�k}�H�C�N��7��~,r'�NR��Rd�.��F�`�,��"� �k�TS���k
+%������d�;�6����5���H8�f�������YJc�3IF9|���@+��E>�rZ�.>-"�s����f����J�m.����E������Z��'��R������#��>��B����0�p�O �b������qF+�2���W��؛<1��z���I-Aadjx ����[O��������%L5����2�YT3f��x���ъV,�#��3+���L��������G#��WkxP�ll�f�u?�pƓ���2����&�CB3���A����ɛ���'��|P��((�.)F�q�6�(	[���Zv�.�pv�6-.��\�~#��M%h���XZ#"��)1�F6�\'��24}ye��χ3]��#�$���0u,11���_u�KY�����Ǵ���]D�?Q�IP�7�8���B�iK��2
���p�媇*�xQN%���l�q02�2kx�qj)���
���\��1�6-M���)�fz"Ȱ����> ���Nq�&]3u�d��Ѵ���r"�_�����P�aO��	T~V�'`&�vBd��r�(���%^�.=2@��q.߾O��pC���+��C�f��8��@�o�ŀ{�#4!x�@Ҹ����콲�Y���<M��pb�S��W~y���۞�`K���v�ۋY�P��	�CzU�����R�I/��/B�!'�	L�~�H�?�M��'A��K��3ҩ5�Շ\��즺�E�a��]�Q�;��pRO�/�t�|�"�6�ķPQX�|*�,e��(-�Gm?��z�i�x�Zh��M���V����x�+!i��)T��D=ɘ��2���52����+}7�>���c�Gܨw��m��p�"�4jEb�h���<����?�z<�~��j��(� 5Ջ]2�����=��R�KhrJ��^����(� ��3�>A"�0<Z��*?�V�l��,��LU�����Fd�'�2r��M�;�0�������X�����U��[C|/�q��pw� a��"�L�Ze�5�������4�Ys�=���ZFG����gc$�ěrT�]�_SK{c�v�BB��|�=vM��ُ�8h�vB���R�b�3�%9|?�������� ���do�K�j�<�f������6��m#C~L,�69Bhu�����0f|[��N�}��%��eZ͚��(C? :92����t�~�ήOΕ�BoOg�L��wb��#����L3��C��O��w�a���||���r3���3`�?݀���-�0Ȟ��(焧�#��<(o��`�B^h{�lk���sc�Y��Bh�A尓�C|l���F��b'؟:DkD�L������^L��*�QWp7O����N"��57�$>֐f6�T�>qFwӪ�����rU���4_ZV��Y-)���t{�+B��%,���$��Or����`6��T�8�C���a7�
,�$��pU��1�r)��IPd�P�<��Q�q*���A�/ӣ��G�@��&x^	�p��
:{D�xY;3�劘{�=8�@eQ����������K���Rh�4��.��l���ڔ��D�gr�ܾ	�u��F��
�����NF�"J�n�n�ȴc9~��>�M�H���6gұ� ���T�0��qk�G(�~$TG̪�¡!�F%K��Y(���#�fk�x�&�Y�ֳ%c���~7P2v�K�a�c��00���V{��j��)H�����~���>�eSW�������h _������&C3E<��j�����$�V���_�yrFl� �N�)$Ĳ�`OK�%��G�^"(Q)?J�p�i�wȀ��F��2Sk�Xيb�ױ�������H����2c�S:�g��65����[�	���C���23�R���3��ۂ�6L:�����W���S6�iZ3��c�B�yC�ъl7@�a�+ؾ��ua�z�D�:]�o���J��?��C��R��Z�?���ɤ��c0p�$���-�	�z�B���@0��b�&�[�/[��I+C=Me���o9���|�f�qtH�>��6҈�?��E^��h�
�#dt|�a���J�mq�L�&��P�S\�^�|����q�r��3�&. ���c�&���m9�ۄ[�"�LE�<݅�Qb�L6+�yk`��*B@��oM�?���Ȱ���sr��8��O�q8��2VYO��R�R�O�?a��Jf��Nn��X~R}?��8wV��]q���9���)�:;�#��iA���6o��+c6�DǄ�r�S�iK
��gd�e �G~Jg��\l� ���@�'��W�1Z]I3NpBa���̚9������|��
���!c���xav�9�s�,��R��H�L�zo
Zc#���u��<�.K��=���`�D�oR(k���R��n�V�W2/!�g�4�vM�G9�KW�47�*��?��Q���:�����ge�p��!��,�����ϓx|�B�EQ�k�t�ڞ�ǜQ*���6�f��眝r����S�G���U�|x�f���0�ٽV=O@��}j��B�t�����'�N�e �k�j�n}�ol��OT0��u���-V!�����3��-=@��:ധ���œ�X���7�:�l��م�5f@I�����J�w
���^*Q���
;�9�Q^�>��*�Lj�#��6i�{������.��p�� ޘ	����E:i?;�R�\y%���Gƃ�Z��\.O�(�<��Q7�G��G���ޠ~�]wA'��Q�̷OL%��<�.m�<Rr��`����h�j'#B��k�3�C�����v������16��ur=S:�S��w)#��d#�Hv�kIY�sF�-4p�?f��.��Ƹ���i9�[�~c��b�rO���Z�1)hg1"DR}P� Z��0��I��P�b���u(�f[!]���'�^8<��ꖋ-�C��Z
[{H)[*���F�r�Q�ZM!׉��h;�32
ú�U��Y^]����|{X;�q���mQ7�]"-T�{W��?���ccOD�e�b��@̠f�?�V��r�g��7%��Px2�������BA��Kyw
�L<���+�(L��Qk�z!�ǂ�iB7�t}z��Rey��K������b���.$ Z,ԾS�!.[b�L��� |AV�:ޑ�ؓB�ufݘ�`�Ʌ�-T焎9v݉���ķ�o��KVt��.5.��n�`Y�`>�"�*�Cލ����S\�w��G��j�aM���������i����yM��Zj�Q�^j}X ��"0T�0?h��:���[9��)�c��}������b���OR�d���O��!��������\613͋��W�=�o*�e�I�k#����]��~�����~y���MC���\Y`�8IiKi7���c�]��c� a��9������ԯ�>�g�|�n�aj�F[$j��pް�fJ�?.n�Ȓ�+��gW�mSFe-���g��b���U��'���P5e�ef�%�y�u͵�֖�r)��9�4��n�����]btM�G{w�����;��R������/��b�K4?���r	A�(D�%�[{�v�~���x��>��Ҷ��_&�^�i��s�윞�I���`�P���F���(=�y�aAU��(�h�,t�qt��m6O~NBr�Ȫ]x��{��球C� G�kG�g�gg~ou���P��'Ÿ���N�$%H���a[g��o�)��L�b����[���{��y�����R����3���h�t@���ʡU�U!=�?�����j�@��rN�D��d��NE�ӵӴ��vb0oW3Iu�����m��: x�#PsίY�ژ�|�ӲS���7
����_Kq�]DSX��f6>Ҍ���� �!@~�-2�b�疙6���\�tu������:C:���ìϵ�A6E�SK�@u�'�x�`�V���"�6��gW�S�i"����i�
�0�D��l�\�.��h6�%�[�o+�$����K@�^N�����$��!�͇��u5S�3��@ڡv]!2q�)��l5��/�.~�$Ģ|�z{���e:�dp�����bq�|+r��]8
������l�9{a/Ei����6�G%~����#�~��pV%B�m]+O�i�L�KFs�nPT���F*�B�'%]�\c�l�Y�.��u�
0�62���: 
��V�lTS��'�U����wl!���(��S�Pi^B��S�{���m8��1[�5���2`�u�Oe�%��4*�`B#R�ƆU>^�=������2���?��|�C�m}�t��
4j�󓎨�]S��ٴ�3���j�Ɔ���|툫!����]�'#pJ��Q�@!<�SK�x��g�y�8�U&���k�俆�7�0?R8�+a���3���o�0����X���6�_�lc�]�w")^�x���o�~u��y�(��`���ǹ� ��ܵ!o/�w�R��"Fcz��'�r�� �]��e�ԅ�����&���Bπ?m��/	�g}�P���X���C�q�\PV6+�-��W�L��p�='l9t�jL���T�M�|2�@"�W������o� ڽ�&��r|��˸��ψ���AL�F��P�g�(Bw�p���j�Oh���Ux��:U٭��W����� <[ɦ���o��km�ʋfp���-hDX_�i�#ώW�o9�uRq��s���K�J�>J�\$-��:%�$v�� rD+�b�-�R�u��a��)V��\=�U������M��:	�XM��ajJ|�MF�ݥ��/{I���(��#�g�V�i�f���/�����#Hs{&��#q�_D[�՘�eܕ�_��V���aݡ-��U��j�d��om�d����T&�z���O�P�6{���rY��	�թ9��/���0�E��[%��?֒.�=�Sx5�-�C��CL��b\WC�7��'�`�r��sBĐ 4���t��؀�5O^{F�%�:�y�_��Ѡ�x������`8��(����fy����ݶM��v��~�'s���ߙh���a���{t}\�6�"L7ԩ�����0kLh��K���܎#�bj3pB���0�CMu���P�N���b>����d� ���̰��)5���&��sr6�0�r�эy�M���n�N�eo@'��"kKp4z��dڝ9ql��&�g��{Ǵ9�k?_n��+�����Ӌ�����Myz=$H3����r�CO�̭S㒏��o4i��A�H?��W�3���O�;gV�_����'S���I��U۬��L����>��K��h���`�]���e��n!�DܐX���ͬ|��7�c
�ŧ*�M�tCIFw.$�!S�XH*ƣ$�/Gx ж��l�����}�y�&y���� u�琈�?�+	 ��L�ն��G*�����6�#�2�M1��ȸw�9���/�S������eG�-�i���&:_�`��0�ml�.�v/0}PIH���ﺂ�Y�%&΀���@����R�YG���(�����6��O$_b��t�-FѼ�ůZ��.���G�g�*d)���u��;c�Y[����x�����j �?�� �R�V$K����V���ͧ���7"^87�]AV�$���y���:��]��[٫�4,�[-%XRk��0�l�1Z?M,W��юʧ�ߊ_����/n���.8��u<	��D�C��#��g$����E����H��V<��~?#��a�B��P(���#��{fR1�'��1�jH4�7��<~3��M�XHI�8�܉Zk�� ��-l0�յ����p�z���'LW+�0�p[vM��/-�ʢLaXU��l{[��Ul4A�b�˄������CXO}N����a

$�!����Z�l��*�]�#v,���>;]$]���9��������׀���0)����W)	���<��;�m����H�$C�V;|C<�z���� ��D��H[���$�X\1�'������D=Yu�d ��K�/�N�.����@������IBFɟeT��0�� F�S����J�TB�~)�fA�p���]19���Y�eNE!a
�%9��D��=�`q�����bA��֬�!���eF�O�^+�����N��,�ƑI<��Q%������"%��� ���|��{ �(�X��Z��&}m@w�!��*�1v����0��o�/7�:&����ᢤ�k���\�D��:�6zɏ�&�N�4��]ViR8��άs?ìe��u=Н~�Fp�8����%n ��1��PX��e��k��)1��(�`s4��	���,�Pd|�N*f'6<��1W]�B(6�T��J!&�Vh^����~�r3C��F�)'J�����,b��S*�":	���~E��->SZA��B䙝QD�^ŏ���������I$@��a-���d mX;]]��	zIOkFO�D�3$�<-��캤ˍ�����#`��Y�*y��:"�>"^��n_�%��SϪ����#��������&&�M%��>���Z��B{2�̼��v3؅�d��m������ɚƽ�_�,�L5k�5�U���x]�D�%B�L󓚭p�6}7Jn= ���;�ߙ������گq�"=(�k����ԁ��kq��\�Y��=���3�4#�	(J�4�sMp���ޮ�b�p�H�Eᝫ��#��]#�r!���bT���0lS�.l�f���VgD|`��t������VwUBe%�q�-�����V�����.*Ƶ�-a��{g��ӽ�	�yQ�R졙�t65�h�{-���z������X���Kg��fh�d]k?�d�<��|�,]^��+x�%��A�̘�ؖF��{DX�����<1���N[^_�K�1�|{����력��j�����g��qU��I��z�?K{�9'��f7��_)A¤#;q��N����F� ���k�_ƨ�-#A �z���1�.{p���R�&/a����i^�C.}���l��ݙ���샢�����d���X/�h6
R����t�nA/����;�f�@ Uj{�%.\2M"Aw����7�����Q�k���Z0�Wn;q��������t�-/�=�I�J:5�l������v��/��b��7���_�@��e.9 'U�ܯ�"(Ԅ��E_�����x#t�VU�F�W�!�I�\gV�%�SS(x�a�WL9�N?Җ�-یs���"����ܲ�u���K��h���Z�3O菴�+;����1��lu���V=��FW�)P�`x��zֶ�����홠+p��h��Du,�QB�6a9�U�þ�?�.��gߛ$��a�#���|�V[�#5�`���J���p{�[�Y��!z&��P�C��3!�xDQ/dmz.f�h�MM�_�cŌӇS�P�d�W���w/͕IL$��fO��E,d�6��۱J��s�6�p�V�#ː^p�� �L,���]�y`�Yw�%�����5D��!S�2��(���s�/�^1V}�ƿ��������L�#"��q�wH$�A��UH�G�H��dbZ����t�Q]p"�]jl�e���f���T�ۤ����h�c%�1�[�IF�=��!Ck�N; �%K�ʀ�&
�#�(΄�����:=�f���w���{�mcp7\|�����bw��
v���7�C��U5�G��� G�'�'c1$HO��î<��(�"I�oi@�S����-0�-�bJ��ƾޝ�F:�Y��-���]�5�F�]k��^h�Upp�����=��1�_k���B?���~C�mϻ��1�����Ѻ�(jb���k��`5R�ȷ�w���9���~�f'�.9	�^I@�
U�\'3v�����+K8X��g$G��N�xNC�0Qd�^Ώ!Y��ۮ���$v=��ewc�8��Iq�b���2�wV׻d`6a.�#�2�*c�/��N���%�����������5'�xH���Uk�K\���5��v����X_<w�VE�XVmwdtq��]���lΥ���5��ѽ��]ǭ��M���b���)f+�Ti��8R���q[�y�>kF2F��.pԲ��C�)��5��U��=��V���[Y�m�۶9�8���(9l�D��SZ)��P��nZ#����NV)b�P�MM����Qw���"��\R������8\#��'+^�&���;A��W�"�3�TKc~�n���+����LKK�A���8�O�և���>�B%��w(��x9�(��[���(�ǒѶE�����{F4q@�21ot��J�C#1D1P�\:� ����Y#�b*�G��)C����\)�i&��M9�7�.�J�΃��;k�gQ��|�:�K%�(jpVF�%���^r�R)"��ƪ@��KͥRaS�ղ)��U�H���p�f���x��u��C��r���L�S���tӍ���BX^�*�;��H�3�J;Tf�N!`v3w���{"���D�Y��21X�ȝ9�ݕ|~�}��:gK�<���9%���f�Y���5?�DΜ?O�m�c(��^t����~~���Ms���w�֙\�=ߓb�c��W�BC�mD:W�����|Q��m֎����PQ�O�JN\�PkW�~��e(���[��mksnZ��L���Gt����51B	DXU8 2�����!A~	(�D�͒[i6#�_�c�ex�Bq[���v�B	���e	`�LՃ�A�����7_����ۈ�S5���R���V<)���_��'����%����:}L{�� �IqF3���)�����e�ϙ�?P=�ˀy�I��"&[�"�H������(���`��kfղ��}���e#vI��՛�#��i��^�����toN���!�̀;�M�>Yʚ%���'�it�r����,�ώ:/U�-s�ĿY�o\��{bW��Gt̗lU�*�lV�=j,�ָ��dvʙ�ێQqMw��v��g���`�I����O�~��E"��RQ]��M�u��o�V�`|<���J���A Hյ���}���M�S�_�'�Ǽ1��(�T~{�c��k�~�L���}t�6�h�'�%���;����|�L���(o��g��j�ƿ��QG��	pOzIs𻚀� rDC���8�\�T��ҎC�,-�Jv�ϣ��
9F��
�5=&=�]͏ύ�|X�c�q�(�K��6��W7��2@j�̤(��z��ꐌ^H�IZ�E�k��/#n�6��K����f�	6��������y�|�>M��E�VG�T%FnwIȫ���fV64�xZ�Di)k9�AVUQs5�@�X�v|vꎵM_�������l��*4�<�fU�~�๶u�Ҁ��wU:ļ.G�^�d�W����)r�\����H=;n��@�>�Z��0�2E�� �f� �Y���}Zw&���~�d�ɯ�"h��{�D���6^���5-���GF�Hg�n���4�[qb�Q�y`y�.��u��h�bȳ\#�*�jc����;�yh{�E t�l=|p0� ���aS��S&����B&�s�p��1��W�5�����a�����m>��	�Z�
R�[*�㠶P���:�3˓��}��aT��;Ѹ�p>�W'�	�ҷ"H#K;��������M3���<$>�U  Y�}2����y�џni���4��7��e�|�uɄi*Bz��,���ˀ�1y괤����,�>�dnOi�[�\<�,y0u���7���?*����5RZ���c����]a3���e���BO�ڕ}i/�J��h����x�<�ao<�L P�@�9D��v����o0?��������&����kEl�*UZ��G/]m_�D��*� �[DW��9���@���IPF��j�DЋc�Z(�Ѵ!s
�3��4\E�T_T��y����`��ֿN�g�92Qݼa�n�c {���ԨI��
�w���B*��zx\���r�1K�,�y���\�>^�{�^���-�$��L�N������Shk	6��x_��eWM��d��!��|�V^�nf?]&�]d�JR-���O�7{�,z7�.6��$r-����QB�j���Y%w���?@ŏ�y.^o#K1Uc�f7u���I�}��S�K���Z�Ie�o��	��˵�"��yn�fsI����q װ���P����2c�b=���r���G,
��T�<�k����?�<]D��M-*ހ�n��L�^���v?��e��n,����-8��O'�'�m�ANQ�'��q�k�cu���g�����X��@�P���y�dNJ�ҭĭA�M�3���z����]_�K�L;�h4��,��ۛ��f�C�!��6��xpcvV'h��O�1�(��,s2��t�h�V��xI$�g������A��&�v�v;/�W��0M�
~9�&s��37��N�c�o� 7�e�� ��}	�������
��jY`��Tʴ�q��x5��fU���'�W�~Y���	�TO�i� �u���U��'1��[_䓘���[�'�C��r����lX����
�60E�ƒ��"B8�N"餏���g<db��0����%V#]/�=Z	'�.�!��]���,TBlO�(��.^�'��V��b֘�#����7�����f9�)��F���P�q 3�{<Ԭ�[�!2b�H��Z�7L����*ob�mys�ܐ�'�c��Djܹ4h#�V������[�8�xeؚ�9^�3�dߍPta�W��_�8���a�(?�z�K��*o�$!8~���b�A�f��8��k����o��hXޞ�)	:���6*�Z��t�@�e採eG25(��������I����;�$�����@��3=F��BYP��zތ�_B`w��7�7VU�p��N^��PE��)q���D;�&}�������C��n�"�S�!A᭑ty�8��ڻ���N>í,��g��]�)n�I�����Ւ��NA���Z�y)��+i�A�]�hs�yZ�q8�������MX\����h3���_� ���E��V>_�K(O #ڍ�m6|i�]��\������+��Q�^.r�Us�#u5����p��MV�� ���K8�)1��?ZQu� �ԙ�����\��\��|�(�41<�L�J�a�<�=~�����d�~; ���o��Mk��z�o|s�5:oŗi�0��_�|��5������<篊�q�Xh�9�WɤR!��=��c�G��yϝI�658<�A<9��J�C:V�x��+��~��Jc���v����=$9��$��x�5)]�v|�ia�4�k3�K�D*�<�VG擂�(�l�	���ϣ}����;Ƃ��/9/�-�Q,�p�Xt��[�0#�-�ux��,�UB��̯0l6#�]#��.s�vt������9�$����k,��j���~4-\��i[f�f�F��qD�Ҹ+\#��Hn�|�Ƶ����uV�.h$�mȝZ�}���?�U]X8)�槟Z��,�{��7�[��{w�@pd���`��@���A���Z�Ji���!%mG��7�����c�hڋf�][�ZX����-�U⃞�3��r����W�ԢQ�"%[�
c��E��@B�;-g9��?$s��	�"��p�7;����a|0�qc�<7�ez
���*��< (w�*;6��<3x�����JXь���_�|�E���-�邁��i����s������~��9E�6�H*�Gs�i�Ve�ۣ] �a�\�?�»	.ٴ��C]r|�Zyź	vݹ�= .$�����<m�ˌ�j�Q�8��Fh	�q�E�'�:֐�z���3�͌F�4"D��T�DT)sVE�:��u��_�ѕ�{y���<7))'�̹�~F�Kּr��&h���<�5�v4�)����	���X��W���m1�DGsKCg1L(��0��ߐ#�<��V�A��*R�@�Xum䌏�1���:�U\W�����|�o�4+����sH!����ZL�����(!(��Z����|��-�x�.��I�����ﲥ�l���)�a︃K𶿙ƈq��A� �U��oc���:�%��hX��5��]�3*!-9��@H;�F���ā>^�o�� �;��<�_ސ� ���ȣ���<�7�͸�W���K7.�c'Zń3�3G�FD�W������ :���ޠo� PG���s�o��ḯ[�Ŕ��C����`�H�djBՏ	V�,����.�q���˞�~� ��ұl����3Ns���-�������#DR��Q�v��6�Nry���Ӟ��Y|�>�?�������91�o~A��H�"22d
�����P.kn�0��Qm�ڐ�U ?�����E���~���F�?�̣\/�.TNªT4�⽧��J�T+3��d$��B���Z+![���`C�e�xg��4�Q��x�F�J�c=��I����1Q�vO/��Q@�2�9J4ȭ�F��?y�l��O��RD�× ��+��D�"8Z�m=����uµ�2���T��]�  �b������H����H`�9�\+���C���q� ���&Tь�l��:�@^v���~�/�ܭ.�Ҧy���b��S\FT��=�����M���� {���8��5�KV찖k�X�k�~g�.����[���^1�fJ��z��C7 ��5�]�:daU6������~k���"�U���Q�����_^Ja2�80�@��8NX������N*;�`0�{���Y$���6��g<+�y\���&��;2���Q�`c�e�G�O
v�*~..0� �G�}v���F(���1t�dD�^���]��8��OU�)IoלCc�v
��{����
���Ɲ_�~�xMV]y��B�oH��AN* Y%��I$M��6rl�y��!=0�D�u��H�پ�s�\�nuRD+�'�_����?���L�&
��l��fq���R��U�U�&bgғ����ZE�w<��{�ң�����n4�R��k���V6�RV�]Tp�i�*��_(�TYv;s�F��[�r��Ws�텅lh�_xj�[����G�%��^"���2��~��de)�n��1�*L��_������;\�YXNLe}��n��[��פ
�j)�;0��}���@Έ-�?I�1��x���?8|�S��u�[��%��V�+�*�e|��S��٦֛����+��+�;A���T�����~ސ{�	��/E"�˞�M�f�������k�)@���Y�����CQ�>Nruo"�9E��}�>�s�R�3/�x`����xEo0��jH<X���[6��S��}U��6pó���Q}�(��0��r�!c-�����^���Uaj�zv&ɀ���+!��	¦ȕG��!�,`C��f˅�[�RWq:ӥ�G��x�?�2a���D=��R�dV���	�V��UU`�o��[�iMϒ�����*��Y(���j
y��P�	@U8�۪�t���Ps�Wz ��<�ǀ6>�k��AT��pf�7��V �x*�#v�@u��}FB��I;��&{�0-dN`$�I�g����i>�δP����?�EAx9���=��$Y� s)T-wL=.V��W�NawF��>"��/�X1O������p�k�f0���dd�|���"�k�k��<T�;Noh��`��c2;vv��9>�r�����w�XO8����b��dU|���P��c7���Y챛�zb_Te>[c-)Ш����j�}r��KpJ��1a��5���sS�N_?q.���-�k
n�!�۟�����M����Y���4���1�?��[m�I�.�o}�ꂏ�I!�~B�Y���(���iP�����o�W��%��/�/)�l`Z�+�?q��EY�]���F�>�ۍ���E�!1�e���U�Ui�5�|�q7�(��	�N4�:")�7�m�{w@�[R^	)��BY�>j�<ki����:3zY��f�����YGP�9���lA�FA��,%ہ����r�|�t/�v,��c9����xs��m�s��;j�Nʤ�+I��ld��'��J`[�6V�
5�Ձ�\&5�,q�
��5cE��q+A��C�cz��ty	��u(�f���A��ˏ��bAVq�l1H0�Qv�G�wCG�mȺ(I_JkMN]��$д���t���qM'�u�N$�_�2�w�/�>:Y|���7}`�����a=�}E	QQ.3��W3l�"�
r�B�+����*��ix)��	_��o�Q��`�$�9RjXB��jJ��6j׸F(`�y�!7]�`$��� ^�F� ��Z��(ɶ�pm�f����7�nTd�!	om�T�4+	�N��Ojxa�{�`�q��P��M\Qٕ�gC/=�5%c:�n͒ے���3aj��ۤ}�N��}Ɉ� 1�Fk��1�&/Y,<P�w.��7�U'5I�TZ��f	���>�_��+�nJ�ĸ��N��?.ޒ
 u}���x&%�0>�-�Y
Gd"�J���Ba��sD�2� RSS?��d�o�Nb�CaV�(-�,��L jc�8����o�5���ɣ}�wɷu�q��r���$���X�_�M�2�������q��y�6�ɧn��W���?ڂ9����4y��-qu���@�O���Цx�6͓æ�m1�8]_c�r;��R�V �I*4X'>�F�xa�ɶQQ����R�gQv�������	�W�0o��\Q�?�s�]X���38J
JJV�G�9��0�^��}3������I#����w���}�����'v�6�F҅�8�o��b�l�Ul��Υ�<��},�T(�p�ԁՀ�\rk3Vf�-"��7O�$���{W������WL�h 1����Pfv�s�VL_���9+i&�Ñv�������|6zr��m9���}k ���40`��.�DifC xe��x"� .Ɨ���l������kI��lS��W`X������@y�Wv�q��Olf�Wg�#��y�7����%��۳A34�ax8~w;ْA4�ڏ��.��A��}�I�{P�~Y�E��&�v�V����3�
��,0�~ZQd[iH�G>�d�z�`h��3f�����0�X��&�4AK3)�����p'��$b���ߖ��a���`I����uMt0�x}�Ea5��}��K,�<np&^��`Ӆ|��.eƪ�QuF�D��GF���d��	�0�̗��b�r�Ia���j{�َ���I�����f�c��'9��b�!�����8���"^u��Vq3�Q
��X#�Jj� ����u,��@�/�C�a4���3{�Y��>�3N��
"��+��Q�T�w�p[ѽso����Zp���P{nf��F�i�}��x�8�Y�n�El�M��+��+C�3l�g�������S,!6@������8X��y {�/Z���O�:+�׻�>ª4[*P��6b�B�b��CԴEW)9[��S,�Ѵ��.�0H�O�@���1�ˠG��o�(�;Jz����?bT�f����%H�no�#-�]#~G��-L���/�������qn�M�^�qM��uu$:�Wn�8����藞�C�>���s�B�A����j��u^�: �*��N�}��kezaΨ��%b/��,ı��f+�<�<���}�#��=[t�g��.7#��Q�p|��#W���ͱ:+"�!�ɷ��3��;�ǔ�mm~rFlI�]�c#�3�B�8Z�w��5��\>�hA0��>�^��@RV����f_�R��*�To0��>�Q6�w��b��r͓�9$�$Z���[(�A�i�T +�D����y$��D�t����ؗ����s"f���o:�m+/�X(������A9e������mz�R!��r{�A�"��)�l��Z�C(�cx��̐���e�Zso��%G)Ķ��-ŏ���^d]���cL��Z}-�Y1��Dy�|FF���՝�T�y�!�ɤ;E�/8�)�W�%Cd7�N?�
����i�Ͽf���:��$�<�3�,�B��[���URɶpw4�?�z&Z�1F���5��	�G��e��r�(��7���^¸���o���hmB�^�I�=�+�MQ?�!P��,�PV�>����E�,��Q����D*�3b�����V���{PKlSê�u��\�K�������BL���p�uۏӎ��n �
/�ͷ�]Tf�J��x�]V�*Ub���#7��z�}�е��x����w�".�����I �P|h;��P�ơ�'�q�-GV����է�B8߻�
 \�����L:1sx��	>eN���X�j#rH�~&D%�L��<ZJ(<������߁~�J� j���hl(���ޱ .X@n�*���C�HaR�H��J��Ga�#���u��,�H�����)��4�
�;	j3��ad`<����K��3Ps/(V*���<�ˤ�V¯�d��$Ul�#<�	�DoA!� _-}��&���v<4�e$#��fϤ�m�� �Qh}q��Ѕ{T5H_��`9��4	sE���L݆*�a|Ibɵqع�Xl
j�{��xӍ0�"��MJIO���D&��Q�����B�R���?�@Ɔm':�Y|d��1�״6R����۱	h~R��b���	�`��Kd�F�4����m��T,��|�:/��D"�� ��VVQע���)�[��$�Yɴ���a��թ���[��s�&k�f`���<�������v��i=y�f��&�'�ɪ�g'�x�.��z�@1P���.����mT*Ek�䤼�Y�A=q��V-<W�'f��Z��7��y��m�8��N��W�e�/�2�+�r� ���={�X�=�����1�|�V�@��E�nt��G���d�t�R�O��"-����ܨ=��܊��ժ�_]p��6��Gk׵�]�c�� h�t�7X��E�[;���^�b����q�W֘ȝv�����>w�X���wz.`��W$��
Y�I�D�k:4`�^z���ټP~�|vv�����}�����=�u8�ړ�KA�����\���W݄NA���O�ٔ��'H���4s���f���yF�'>.R��4q��6;9)��Y���nbE��f;>b�;l��d�&4Z7C�Β;K&���z��`����:zq�Z���Ӈ`�1�s��f����͋�r���J��\ ��(��f
��%d��R}~��^��x�]�{��H�`�=G ��NGG��-�Uɲ���9l���	��Ul�ʛ2̤��
�4w�{��%R��<&B3�E���1(P�[	�}��>�RTid���tIm��Μ?�p���!�rE���=d���9�{<�w�|+�Z�Y�XH鸎mS&�5��ߺ<��~c��`�:�t�"h**H�x<�(IR��"��4e�-���f��B��,�w4ꚠ�,�%Z�	��-d���h�Yf�߻�;]}�}6K<�]�Q2�D������`4�e$�]�CT��+���ƽ$�w.���3����R��}(|\��XM���<c�c*�^��p�k�LB�?�3pC�M�>��Ӷ�9�}�
@A�G̳���p����"8�z�ڑ�F�B�h�+I�$��_���q'��c�(���:ܼ��-T:����^0��QL�^*b{a{��;|�+�r&QD9�o��0�c͘^�D��q�~y�-1d��Ѡ!7Qn�j��6��<w�v�W�	g�)-�d	ޖAd�	^w)�f�����O�1g(����f�t��+�!.��c���aiѱ�u�������OK2�Ѵ?2��m�u�;j�C����N��GzW�PA�a�rw�'���[��3���V���&߰��#���w�I�K��� %��(�H����h������������R��H������7rl�ѷ�]�&�F���N�lI����Oh��d�L=�����ls5;�,R�I�5���7����Ñ�ZD��[��(��-�](B�`4����ħ��W�n��x���D�j��nۈ�5!�ۼ%�S�g���W60�w��&u��k�=.*�-�ی uH��m�\�k����I�L����cX�0B{},�M��o6� ���sr��yAY�[0�'�����	��N#U�r���<T�����t������v��K��޷�k�8�)����pR���Q�y){���n9�lej�ε+0�D�i����`
T�0FV�9�;�WR�.ζw�a.����}�#���m�޻��/0ۑ�LS2i$�l&F��~Z�)�@��o 0Yb9�>�_��E�ʦ�Ʃ;䉲�Y�ok�,�����L5��:��{� )�i�#Tt2xxa9ڊUP�v�Ơ�|lO�o�M������I:�y�t,�C"�<��|��o�؀���f�l��X��<�j�8�UCo0[M0([���e͞�^��8��t߀\S�䏳�~�ؗq�=GA���{z��\C��4g,eb#�1rI(�ʥB�W5o��ٍ_���S6��<G�;��t��������[�n���zZ�����||��^lM�{���H����g=�Gw2 �P~?��U
Ǹߐۮ�-&|�����9��*q�6&��&` �!�UX5�5ApU$���KP���д���� �?q �.�
D^_2�_?���D\Bl�V�L������
�(�"�}����`�.)�h/'���o��q�0���IO5L����t�����{��#�ߣ����⽂���u�c�O觹k�l�S�%���;p����������\\��V ��F�l5���U2�0l���͍b������2��{�&�`Y�\�BY,��#��,~���t�����r�C�$ʅ�BN6��n1cq�3�Q���S��e;��v�̽����t��t��,����a�H�-St���)�g_�4}��M7�SJk������c��OcM-B���X4q\~YtQ�d�F���}�Q�m�4��\.Z��#��Hb���E���5��f����q�$�ɻ)��4��}p�]kMX��M#����-�Яkh׊�,�Qlm��fg9%1~ �6c�	Q�a�+ ��5)���q�9�5Y�ᦱ�M�� k�����
����0�5� ��7�U���r+��#f��펉��6��j�Q�Ѻ��!!E^��M���i(��~�g��u�5D�.�ɧ��^�<.;Y��<�=�e���L��'$�l���G�Gࢴ3���@gS��k�a�v6ڣ`g$��
���\%�odo?����X��V~�I���Fv��$�E�{)�K��w={���3Vz>"~��}(���GY�9l����++�63O��X�OA��T|��J�P�?�rٍk::]���c�͏�2qK	i��t2���W�!���H�*�5���G�=��Pvy���1+�u>�sL��6w�V/h������@��Q���aL�7U���������0��$v��վ7
l� ���;m��4� ����6aZ8���T,���ںRZ�֥Dp����DƓr/��Ғ��IvH���T�,����ms��iP����s
�فLU�@��}B�V8���J�����C��O�����-�3�HV�UQ�}a���<T�Ff=����~���[h�/K�䧄{��9���+�)ѭ�`��ؘl�3�% L&"��o����\��ހ��'�!ˀ�֬���1|L|1��ĥ[��%>L����S������	�5"G��1��}ie�7����a���|
�ڪ��T�o�L��ی��H��X"˽ġ��1��oX;�s�P�z�D�ΔW�6;�1�R0��֠���l.��9[3Y^��5�5��S%Q6��wv�K[�S���1d&�lx�V�|�{�hސ���:z��X��ϩ¤�X����CZ6��I�_6(56V��.E*�~sI�B�/����.�.��_&�էܞ��Ig��>�Ӡ��!�\da@ �@��.�X��%�T��6�W'4��(��9ܨn%��J����1U�E��n�l��=�@�9H(�kx��
��A��>���Ů]�w+��8V����Go�aob���V'����8���+0�����ų�P6����QŊh	X1�zW@h�'�]o�=��\�ӏ�3}2_����È��G��P��G~M��%S���AB������v��5fP!��>�g�dI�s�D�b_%�d���A��[U]~�^��MjlⰣ��j�Y�7���6�伱bd<�G�L��GH�.�r�����[j�,~-�$��a�`������x˰�ݫ�io�R��A���Sc�x����D���5d�o��!�m*��>{}mn
ҫi+w�0�������V�6�ݎM��N��l�=jF��M9��y�Imϵ��*��T������i_7�h��2��*=�#[�E8�����C��;�*e�kH*_>R\5֪�7B�bh�K�X��01�E�����OԲ�X�������A��m[t�#�0XĲ))�1moYF���)��*�=yu?r�FN�ј�W���s��	��u�����d_ȗ~h|�G@�ӸW.�2�`"Lms}�.��F�)����m�n]@ǹ���Z��1�g���mNC�:����'9=�qfQ���
�+/��k���.�6��ε8'	�����\^\o�]r������<�{�̶��h��F;��X��ST�����#OC�����e�^� њ�w����Oce��p�J"P�e�e/}��/�(,(}ҹ�$sJz�R4�[��Qon�A9�����o�>%��r�1һ���)��ȑ��*��r{�W[��z+�3x�*�l��2w��g�Q�}1���D[28���F.J{���As�0HhqAJ�qW�貎�+�0��Q*�6��hp^��F��hK�z2�ID�q	��b��y؝�c��%a�tgd�c&�%(�1�f���X��n���	-S��$v���cO��(+��J���G���в{�ݖ���M�upADظ�-���Kf�hzXF��<ץ43*�p�Y�a�Pvb_/���Qʗ����%��H�qHi�9[���ڵl���;�Bm�K 's�c���򰺛����W���=���-
�*���-B�JG�9-v��LJ���:#�Q?V'hn�� *���s�/��-�_\�t�5��V �EK�
y��s��V��!s�,�">�?�m:��L"��2�u��t�1����2�/���O
��1��yN6*��ȥG�1�:&(��G`��E}�r�5йKA��> {C�S��H�H`C�(�fbY�D��� ���^o�]y[N�&ZҹK���a����٩���\A�8H���M��N���%����@���UHt�gP.B%�.�X�䚌4P������2�-A�`�߽��0Lю�1�v?`�AP%��程 B�e����ß��xZ��4�y�[:�Z��+Ư�,&�F���xe���F�DD���d��Z+&�SӼ��T6�����l��r�\໸|������K<��K�wO��m�z�'�cQ�B ��$[z�мM>�M��ʝ��x!����s�~̑�$#M�]+���ܢA��#��'�C!{{U#���:�<O���@6T�)���+��ÕO�)�g�Q�iM��c�@��ӫt`J��Lh�w�+�(�+a~�7Z��U�J�l8��tKkV���peu�i�u%ԗ�H�Pא\Ok�lh�������z���;�3قip�b�(�|��`�n�7v�E]w/�s�5T�.*͈ܙ�rW�)�vX���)��z �⫼M�L��F����uqK��w3�[)�\�f�]��7�N�?���'��r�����@H�_/�Lߚ�W2̋Gq{���_�6t�f��O�,�gEɧ�p�8�X��E���I�n��L�5�9����R�$s���Z̪�̾Nˑ��Ԑ!Q}���m(p�h"��;Nfq�`啐��K�a�qO��EyήO2CW���eՒ���`�g�5��C޾����$�Ѩ}Gݣ��\�+L�9��OF�nSCV�ؽ(���	�g�q���y�G�,T2҄Y��hh����1_��Ncs&%�>e�Պ��Efm���x���f��ߜ���5�l1<$���r�JXx;�O_��d��?�&%?7��B2�1>�ߖ=�"�g�[�qޟ�`C���p�U��,Xi �/��+V\
@b��@�}�E�����+zL��	6s~�g��}�,i�YS>��'4ӒW�$���+;���f�����?��uAa��K��ab�g]�n�a��=���J�i� �	�UW+r�|����N��ϳL��ȖjB1j���-�S��D��z��G��~u�3Z��A����[k0���.�[���
FfY�kF�0����3�4M3{����1��jW!�K�4O>�ԧ��J�)'O��V,���R���1�ŜH��c��Ec�����k�2��;]G��]"X[���P���	��'2#]���pX0�>ʵ
+O�g��e�#)5P��m�N�i;�D��V�Ӫ��r��������#W��Eӕ�'[w�O{�P�q��y��lRbW��#�TyP9;_�F��O>m�s��:�y�N�[Xj���I%�풯b���KrI���=� ���"��I�[�88cC`�(!h����t˗q��g�	T�y�lr�*��`��1��A��S�./H�&c6P�]W1�pY�0&�[�˅U�4	֏�9X��Ɩ�����  �%�L�`�Wp�҄P��ĝ�(N��yr�
��=����Ӳ��g5Vtx�=C���%��R��ݙ�\h�=
N���ѯ� '��O����ْ>�&����,��*�}[�</s����a�B��o�
����x�r ��<T5���f���us*)F�D� �`_�����O����hrjf �p;cMp��MH<����l�os�
�u��W�����LI/���B�|�wsmQC�A ���]���D]�8htu����uR�w[��� ��ۺ�Ϩ��H��S�N���A�ʋ��^ܾu�L��l�+�~ =2ZXƨ���Jw1�z�?>}]j��P�7'��P1MȔ^=�+ҟ���x��޾�/��?`�������w���LChek��ꉞ���� �m�����}���{Dn<߫�1c�2*��f�D֗{����t�&�YLE�:mq�k�Ns|�|�n""c|;;���_A5�F�;�E��ƫ�:�`N��R��.��/�E�o��f��cPF�G�y'u�T���5�ޤ���/^��Gr�\�dSO��}���&3jx�i�X�� ���$(�hEHUH��p�Rʃ���1~�Q�b��xu��4ٓG�>�J#�6o���^�&�-�Iu�[#F���Vî�1>%�)�O[�<��q5��G��D�湸@�L�~���y^��T�l��8���n��4�!�x[��O!�k�N��l^U90�`9���D�� D��E�h�(�ܣ�+���ikn�Z���"ˬq���ҩ"5�'X�7j�'��f
�����]*�y���\�����-xSJ�����mצ�)t���J�o����!5����*g�knk~\)��rE�$�z�(�Sy��v�m2��k�:3�N�f����T�Y8PKA�ѣ �Zѣ�ڕʁY���Ӓ���[�T����:�zn&m帲��0Nf�
��v4s.�>�:���m�:ڮkԦ�_:�!�8V�2��p*�1�F�X���$��-i��,aO�����6�h���x��d���"7/���O(_th's�ȏ�\�D�68�$u�G口��H�¦��_z���'����d?�%4�_I�p1�AQ��k<E*C���2�~��*]�u��9;��R�QbB0P�F�%�W����M{��4{����jP�_�͡��׈L��8�fD�I~(���x<GwV�e'_�1�r#�'��� �֫���u�tw6�ɉ3�	��������c-�Y�0G��"�q$n�a���Zȶ�)U`yL����Y8�9\}��6!@5��z`��%P\P (I�*�L��Ϫ�3ՍGn���05~�/��2eϏse+ [�5���iw�dEp��%0S�n&�5�t��͖?lbXe�G[#��s�Ź�g��a�s-������/����ƣ�6��0���q�e����86�+�҂+�8���_p1�8�J����P�ʱ�y�f�W�gVn��慪�TDߛT�k��U(~����>�u�bh��J����U'��l˄�3A)/ԘI�7��c�VV+�Fy��`ǯ1�l�y�8M=��eGsWb]!aɏ�w|g�o�9�A}�ޜf����γ��kr%�?�5��м�l5�$%PH/�4Ր�����Xj��I�3�����ͦ��D���/M�9�g�bN�">�|�wM^��t+O���pcc+f��D6o��tF��p�iL�g�v$6�Q��ȃ�sM-�b �gFflXw��l����u���9b�\I��%�>�gmB�{��-�4��O�]g�7ӌ$Ed���)��Zk�.���cY��2��$Y�TX�nj����s�Ԟc�mB�|-�մ7�V�B�q�,#"U�p��l�9��l4�b����=����؞���R9���7-�`�eWE,�K>�v�@{R�S]w���:{Q�#� !n���$�	\��wW�C��ޢ}�ͷ+��O7��m��ٮ��F@0�6��u�ʀ?��$;�-�����߃uI�\$�-ɪ�0����}@�]�>�u��4�yM����w�]��������W0Q�\�}~�&q8�§�.|_X墂��o�>�2�=щIs�G��+��`����ƒ�T��F��q�Ki*l�m�:������5��u4V����,��j q���|�U(��N)�c���3>�����(�K�W,G�|���l]@H��竵
�Ěx���(�P��)�)� :�.�s7&���ԟ���y��X���MV��Ɖ��)0/А�o>-��?���~�a�t�q��ӗ�I!�q�hh�?�9��P�u��h�(�Y˱rO]q�|�"&��%J���]�hQm+��i3�1j�� ��Ys��m�4�Ξ��n��'Qv�cw�..'�ax��J���W�Ye��R���V��ج�+$9;�nFW,��6���8��؍N��5��y��P�ا|AY�e�����e)��+��������my��&=�w��-�MZ}�N�8}�=��\��`B�K���f���r,������(�m7�:����G^��L�*��ĵк2@N[	L&�Ӵ�3��a�e#nx�PQ�E��Z���*3ؒ�3fa�&I�pwX�v|J6?�ؐ�� ������qp�ҩ�LC�pϕ�_�Z�l �n��I�z�G3�&��ĉ��=3�5�M��Y�T�7R�����#L/�CM8k%���c�%`���-ɋNQ�0>�>����R�2_oZe=�Zh����fM�G�	�e�iP����m��6���؋.��45����Q���x�5%GX��b���#��������$��e�n�m"~	���7'Z�㭉�;H��UT	H)�e3�Y��g��zn���|z�k��������{N���j7�e`�f��j}8������Ğ�s��Y��	N?�)7�G��K��.��L��ۭ�q���$w��80���������󀳱�ƊӢN#�(x����P�?�����2�,��ʚKY�fi9�A��?��_�N6`4�x����Tu�����:Un�:-[����SdX�۠L����x�1�+��X����|��Rm��7^��&���O�9x0�;1��*����_��"��:MɄc��AMK- v�^��>8';�II��m�Â#+<>����W��?(��P|�_�������9v�)V��p���锄��e�H[d=e�$Ҥ�>
BX�q��R�7I��J�$�$=�\3���#XV���ƚ������#3jJY
��S��w哮_�z�R^��<ӹ�bst��ۡ\�����N�P�n�E^�t�6���]�ء��tW��T�4��3絛��y<#*滽}#*~<��(~��^���uù5((��H�!�r�iR�g��8��I�"�%�;K�vߗ�̡��MM`�a�-U�:�/����0�b��g�{�y�9��8����={R-G�vn�,a��P��0z��'`�)9�3�ß��f�Pw��/T�6����ϫ6.������%�i5�׉�a��iB{���*���g��S�)���i�z2�ދ�C$�l��c3�,&��"��E>��9.�8/Dz�
���oS_�ߊ�I�����7-�	��5yaZ��K�N��j��t
��p���z�@*��k1^�@.��[;��ᙈ�Kݔw�`�Z5Ot�9p�2��r�$HFgИ�6;|�CK,���X�����f���٫f�Cg���P�-�4#lR)<'I��(c���H��&2�����l�42�����d�`��H�C?�A�H^��N.S��f�SoIo
��ۓ��W�j�\,�!w��Ir_`]�ɳ?LG�&�S��x�>���,1g���.U�ބEr��V>�iz��6p�� �N��=�fW{���_mu���f�bS��Wx7�C�z�C�w��uw�R�S��qaI�؂ݶx��5�\g3��"|DfȭA�H@�s@N�_S�"��APgO�ȈF�
�݃��Æ����������}_�h�Jo%������6�NU���/B��1����[u��l�v̈���G��hc~���s7��"���`j7�]մE|��1�u��?��hAUel�u���\԰0K+W�v��#�̆
�� TA�C@�����:+���`��� �dx�����}SeI,I<�\.��3JlX���� �SU{��	����(l+"��}M	>*[�P-�V��d'i��K�Uf��ܺ��%߅eu}��1�<�7����8������و�+�`��n�)���2��^�-�-�-ja�J�m��	��F�9�[���Oі�h������$������qQ<h�}���^�1�ȏ�1u<~Gd�� ��f'zZ�%�<!-5.�8�G�_k��䥆�I��a}tI�D���2�ck�B0�����$�2/���.7�E���Mm�A:m�QA��=x�8�^ S�;��<����+d9�g�0����Dw]�yU�x�?h���a^�?1u�mn��+�]�O���c9&�����m��z�M^��z���Į%�r���z�� ����I 6<Z�2@�c��qEº]����LW��uH�øk�ǁox4�����=T3�S���T���N��?Ϲ34^ �\wA_����jɉUPj6��i�nY����Q+b���aR��k7ʉ�O���V?D�����C��>WҼ�}a;Ɇ5Y�H�·Tc�|t>Y�N��o{���0D��$�<��r�û��	�wiW z\U5]Du�B"B����x�t])^�/��Fk�V��6����*ܠt[bA�����dkx���y]�O��Y�}�L��������wmLT�k������V<n���&� �"l���m+]X��_~��ke*e���f��tui��5P	@z���4��N�'֘�㮿�eQ�Y�@,�r.�HSv�/�=Q�]�@��"���L/�A����l4��O��)�=�7�fރ�+٭ƦC� C�	���&7�����c��"���}c8��1�.�"=)4j��s�d���	@�{��R�0�lY���]���S�
T�-�:G�<� +YKx �BED홄�`��-�vEހ��N�&]�%���=���Fb�)@+��S��[S�����鯯��x�M釢�oa����콈����t���պ�]����f���<��� ������h@Ο��}K�P�hO�-�Y�����$�����j�{	�UW��&���ɥ�!�M毫�Ql��r���y/ԕ,�#CUi(�&6�E�j��ug��1R
�~�m�x�����<�>�����x��y{=>��Z�C�� L"5꒜�Ёe�+GI�29F�=�����	����)�r)�_	 ��0~�e��ƥ��؜9�j+9#���ݛ-���}ŋ�lC�������z|�u��.�[�gٗ!�i}��H�p��mD^;�:ΥQr@پl�L�9l]+�t�]�F��Ll$��r <���D�>��&� [�mO}i�>Cb���4�:6,���A��x	U�U��խ�h̏ә�&��_.oN�f���D�\�)Zn3�h(8@V"'r�����r�Ҝ棴I���ɤzghR,5R�dR '��2��W�,��Sh�tJ{�H��R@��(�k
.w���l��F�6���KT�q�$��T!�(p�^�o�J����x�|��jHj����SG�-m}�?췃G�$R!���T�^���P�6�F@��D��s����ܝۆY���S%�}�5:��|?@�y��x|��0Ƃ9ӽ�i�rd�;�g�,s�n<e+�F�������&Q���c|��f������Fy?*�˶4�Y9TݛQ��d�h��s����^=({U�O�2w�k|�v���^dS�Ob�6��9��ii�Tb�	e3�L���X�TUE�FA?fB��4������r|a��=AY�y�CľA1]P(��m����<<>>�'! ��ﵴGE��sE��u+`[)4��)��E����H[VV�L��&�d�-z�~���;+x�9��@����$�X� ��'_,��V�D��t]ה|�X�m{|��:/cش���+�uJ��B��e�4��8�Jt-Ոeڂ�Y�	��"����k
V� �ʎ�.P�@^��x�;2keȞZ�:Q��~{|Ė4KnO����Kp���r�_��籇5�_!�Ge��! �)p���,�w�*�P�����;����<7F��u�~8Gt�y3�!���L���8��,�?�I�z�\��Jy��qA��~�2M�fB}��ɶs"� ��!��a/�d�'��Gs8z���)���Y)�f�%>{'��G��rf�vL=�`D�nT|����h=S~�Ո�\�	ֽ��K���GS�IE�B�x-AG-�U`IP&T�7��,�Z���p�t��3���4�����M�r�x�}V�Gۿx��Mj�q��)W���4į�' v��V��=�QŊ]��N|X�x�����"�SGwi(~�&��R�����tw�?���]�c�kbuI��wa��1�԰6� ��ڕNq�d������o�v�@B/7{�	�>pA�aÏ�������D����Q���	���Y��/�`�A�ef����s\YT�	k���xΕb��|��0BK�y���>�y��4�#��������T8߮��o��I��%{��y�B-�<��"���TrV�j��g@��͇�{.�Cږ&�tÊ�H�%�Zѭ�P֗�ӟ�_��ZV���P�Hǡi�g��T+橏�[�1<��b��1b���7'�u�
���@r��a3��xhFz�,|��:c� �\P�~�@�E�ߐ�DˇS�/6{����R��Jx-�JF9�;yr��(�g;	s�x�e\ kB����f;{[j7�a��B�3g{`������ـxGP�)��e�>�^�@�� �IcŎ U���/��Ҥ�4Ou����|�w� �ij�L�윘m6/�1я�sv��nGc�-�J]9�OD�s���`��_#���u�eu�a�`z�mV�b�o4�ʙ���,nV�XXz�� 6t�5X��F��F��|`���4�5��<-GC9�?�hF���B5�F�����c�cv�.[rLAٚ-�E�Sƪk6�wɈ2�ur�L��o}�oi�(�TD����N�p.�@K��G�֏��H�L�5ewU��:4��1=h�;a\�b��2(1�1]0���74Q@�aY�����@��u-
��ߎ5����nJ}ښ�����U����"(.�A$��8����is=��]dߕ~��I��a�$B"}�cN���������q���T�[�*S��s������%�����V/g]D��1����Q�o�R攧TGġ�HЧ�HL���"����q��5��q���!E_|EW/a֐��a"�W ����6�w��� ��<�p�ֲ������5�n�\����ڕ������o�C=0fc~� �A{��2!O�Q{��Z�8 �77�dsB��zv�A�2�NGg���d�Oae��q�����2�����i���>�zGNSA��Sd_�a~���QG��6y�2�ͻa�`kօ�(��{(v�Q6?9G���Ȅ���ʻ�l������ #�4_�$�}�ü�Y͑�nKq�q�
�֩�)pʐ�+���!����.Z&���%�'��3Z�|�Ɩ�X}}����'�ײ�N��5���4#��A�S��j�93܆�[g��i�e���+��l����M��x6�'� T묤�"s��G-��L?����3X�an(�!-JV�2�Ӎ2><Q��S��f�e��uT
dг���(Ïts�c���g��_�-QR׵$*K�?c7�e�x�"�1�y�Z��ȝ<�������ħ��2��.��1S���:�EA��ӳ�6�s$=5,@KA*y�b`�U�����I� �,탾]����EN_74gsh�N-����݀C��D�D1�W��gE2Oz�����s$�3�2%��@$���b.�1T�b�h�� p�;��xr*�מ�dG;������T�~��+���*g���
e�i�In?���yf�q����O�;�x@���є�z�te���S�t4p�l�������'�Sy�wJ��mPF$��O��qbv���隨˦���p�������?C����n���к^z�����A��,�����mݴ����RV[�T��,I���~����\_[����q[͆���ɗWE�|�����4�����CV��*���$��ܛ��3&^`�Ff6�u�aj59�M����}��H9�"�$��A����CJ���xH�Iݭ�rq~���c�݆�p��2T��xx���/?�|oWU����i�2^nm*��-f�a'l�9{s�Ize��h�|5=�U��˂k��U�dս 5���"�BEz*��n?�}&(Owޞ�*0.����"6�� a�j��i)8�c�MϧZ崩��yB�B���?uT�c}��P�:�ϺS��f/;cew�ԽU��U��-�Ў���4G�e{��(T�8�g隉�Dp`}^]��kj-�����xL��0�!́�KOT�o:�)��0�_��ڬ"�{&����l3�I�GS5�o[XӞ��nK�bv8�	����O��{jCu����W�ᭀ{l��z2�6~1Q�nJ"޽sD~���kp�9���r[!C�0��}ˆd�`ª5V�l�.���H���DdiO.Q)��Ks�6v�І#�CEAu�����J�?�J���NSB"L�^a8�:�ܽ�4�[��LS� ��6i;���{�b.�l~��[���F: ߾�w*_����k�@.L[ ���Ơ��5�c��͆�܈�`U�(:#ȏ�L�>���B��m�߃�Ak�
to�NR����C}�4x @{��YJ�e�\�Swh�*�N���f�1	ǭ>��$�z6L2�!4�t�6%5q����m`�:#��S����s��Xľ�	�܍�:�V�	��z?lUj#���Œ`��� )P�b,����p���κ��)l�Wؖ"��u�6���^V��L֗��Qw0a��m������.�t��E��|T@��Ֆ��@,pWϷ)9�O�C���F��\��Q�C��2R~�����/�tI�߉���9��Mm���+GAc��rA�m'��v<dzj��� ��f}���A��X��qgR��́�NTS��*��P	 �HD��Б��+ۤ��P�P&�!�Kg�I68�q�@y�jj�^m
9�53�!v�b�!ˋ�s`0�N���p?bY�o9�YT;�Cz��ai���	����97�E�7vR�N����0wd�O�T}G��D>���A=��hhqF�4������ND���_�v�!�"�Z]vS
�l���1����-n�ad������WU��kPvsux��$���-Ȃ��t���~�_ԗ"�@-UX�)D�����ي�ܿ�Ɗ:4���4|�"�C���0��	{4�
�"]p���%�qk�j����~� ���e���n�UJjb��Μ]�E���ȱ�jl�[��/�O1��~���W��(��]�C�6Ld�ʓ��&�Z�yM~�����<�dل�ji�Lx?2a�n4�R�:�
�a�V��=>��3Y:H�'S$	e0_��.�����&��+����4��pҲ�} \�+=ߛ�0X�)�֬��˪�y�N/��B*UŮ����n,�M9@�'R4��>�N:+p��Dz�Q,���%����H�Zm�B����mo�h�f?]���������r_�w?�ig�^��!�b璗gȳpZ�������3.ǃZ�U�~�����lH:��H1E���m�?������	��7m;r�%M�8���ckj�H�W��?���kW���!?��
Tt���{̩�{9��^:����]}