��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���P<�%���>�8��nW�_1����)^�[rCs�`��?�mD'/�E�NB��ѯtg���U	��L�goiY��(:�j����<g������8��U}�Z�u�'�Ϳ��D�1���;7�h{ҦP] ���'��I�Zօ�O�����5D��$礁ª����x��P[A�H�]�&�;;:X;H�V� �y���쪘É�o��t��G4�i쵸��P�縃O�<�&��ɭ|:�Y�PuN"*�d�J3�q���,����>���;:�,ܦr�-i���iEL},>�J�!Q��>�e�.Bp��Ԫ�Ʌ{}}���3�j����P�F���6��i�U�K�x���һ�� �
Y�m�b��B��������al2X�Sڋ V�0�W39:I��/��ַir��y�?r��Ɗ���y�lwx��a4läY�Jz���AF��t�&\���# ����JQ�p�'�#=ؐ����}*�K�j��'8I�v����vb��˓6��{�T�s�{噋��Z2#��VJ&�Os��wNa���O6�s�d���M���KxX.ǫBVlJ�`�����q,.hj���?f�0`+�-����F�+�ɋthS!�lRJ����ީ����]��|F����e/r:a�C��U�Dc!�r�`����+�0�{���&���K�4���'��Qly�����*ESy����p?��:�2���:�?�6��}�u^����$K�&Bu
8��~eY��q's��j�_K+� g���
�԰N2�HmPB5��M��+�1�ᢋ�1�XS��_��$�0��֡��&�n���eK~�da{`ZV��\�X۾�+X9�$L��%��21SþF�V��|��&|�=3���s3]Ɣ�p��u*yEŧ�t�Pܳ�j��%�d�C�<�x�3�
*Yo"if6K�r�ڵ�6A�
�G&�-z�9]��\_ !�*�*�&�y��̙��D�<��/@�������6�r�o�,7F�6���S}�K�3���t\j���r8�^�w���Y��֝�Y0B��!x�:�kZf:/i7��|qPKaR9&�r���0�� �G?�1����A�+�o:�؎�JG`jcJ��M�|c��.�7�J�=��c(R�!ę|J�	~�_6�y�Zc�ed�l��vkDC*��ߎѦ�j�z���8�*�>�@���6��t���̊�-ޟ�V��QXZ�(����A��`W���m�����9����s��T�[�}ٲ���S�Wx֙���U#�"=/�D��s�C�wc��}2�Bmq�&_��,�]��V]S�r\���w�uX���YRBmj�.6S��x��c�F9���趬�!qYjwQ�I��O:u��.i�XW��vج��53RM�ϯt��?�@�/�M~x}H׾���3h���'U:�+6"e����+@2��9%¥tcMl���{Z��=�T��ol#��uQ6�U��_Z czGLh�rb&r�T{y��'j�;�Y� V�_��!R��7�ٚ�s+��Z�M�k�a	�K���e,��ڱi��@�q7���fa<'�6��\&NתQ�D���A��0���+j��b� .��F葄��N���W���Y�i��&oc��m���¼���# �`�y�-Y���FJ���h<�<`��	;�����f���Hj���B�'_���M����{A��ƙ���DW
JӮ��#`	�a-�v�pP�v8q� �e�jb
���d1�V$���׀��#���p�3f�p�86��2y����?�Zl
�j����2�l�CK�9+�F?��6��-ٞ�&FA������Wxz�������2����a�!Ad���=�W����{�^L�L� 2ݫ	�Ƚ��O�]Ç>�#��9 �ք>�3�i3�M�����h5������>-���F���g#Ԏl�dHm�׾Y� o{��m��0��]�R�B3w��	������~�TX��t1_cϷ��}��X��*�W�zd"���}�}4��2��7�Z�lS_�P
wY��0 ��<)"����
̤kmQ�^��܆��!��q���?��Komþ�I�h<M���
G��$&��^�@j#:��[]�S�㤍�V��7ۙe� �������
��xA����GU�x�2^A�íq�N�ሞ$1hn
H�[s��j�I�ڶ�j~d��柅��LF��?�$��$�t�3��O(T%����}4k�,��u�X��N{��㞛۵���1�J���e߸aث�tU���`��U�3�x랒8��x���_��l�2��60}]�S^ ��iH='�&���i4�����	E�,�=�q��F�v�����"/��5�ۆ�}(y��S|lԡS`�Ҋ	��%���`%�/�OKР���p܁@��@�$I�A��;S��=<�R�b�7�`�4:��s�n�c�&q�B�3=��J~�<L��D~i���'�MYxџq�ht�"��*ՒN���(�.��i)еfAcۨǠ���XK����Ď��9�T�~���$�Q�
?�9��'U3�����x�;��<�#2��v"��kU�K2�ʠ��	���s���T���3�1�!�ق���t�Jy�6����]#P1s�h�,�g'˚tE`�����xV���}��TU� ���L�W�W�r#ueK��U���(~�'6�;�!�'�!q�F�UIC��p�kg�����L��a�៲F5��b�-��������]+���+�[n�@�Ϥ��,��E��י]���v����U]�Tv�KT��f�C���2�:���\r��2�l�ݘg�^�a)H9k���wޥ���1+5+5b�ꄠ�Iӧ$��2�W�Z&�үA�b�u�=_�Y��!(Zb��;T�\W���W�&6p���L�΅X@���M-{B�� [���g��qQ���7T܁jg����
���8��/"�p�i
/���e�z��R`�'A�����pN{��cu��֤�#X����*�Q���d:�G�����#�@BK�mc�ݜMfc����<�(a��������`�ڗ:�V�$H8�_��(�^��o�X��$��Jn��Ec='��c��R������@W�9b���ok���j��ɠx������9J�ZEꃼ�\K
�!�@�*�Q�'G1�ͷRGU챠#��F���
G$��܏<�l�P��fNBƯ��W���)�p*\\���Hd�|��&+@���H���-G]����M&?�� ���mQ���y�*<<4�&��c��
T�P� *HF��O"ճ#�i3Y�0�,��\��"/�?j~��_Ĵ��_�V����j!a�V��:�G��I`��H�>ݵ��y���t;����<r���_Mrٽ;v�S��6�SI�"P�i�ZJ�`�v����)B�/������&}q\�(f_m%�O����t�-K��*1`�9/O����⸔l*����[6#��(�������	K�Tg�N�GKn��� ä�����H�%��g��@I����	�5C���>'���۪"�n�����$��4"g}Ⱥ�}P��F�����/���I�ǣO���E����8g�B>�{��BY{.z�T���W5 Q�C x���5N�A<�-Ov
�*	}ߏ��6���a�A��đ�C���u��J�-߀��ŀES����^w�NxS<_��5g�Io���1[;ɗ�������u�Z�r'\a!J�'�^�?m�R�t"Li@dHJO�-���屟1�7H���D�.k���j%��zd�Шb�`���\@p$fvAg���8�����d�Lح�_����w׵p��۷� <�q��vXO�2�d��w�v�w���o�#g��n'Y �8C��M���,-R1xt	'|'2̒��c�T�Vɨg4.H��tJZe����0��E��\�����ˋ�+�j����ګ�Rp��oF�X�ckr��!߆�Nl�!�'ޠ����gb�W2F�ZC|�p8���u�c���Ȋ���ie�W�t�I@�"��U(يm������QV��y�ˈ�s���, ���5u{&d�r�{��/l��k����d�f��<��t.q��V�dS��:��F���D?"miO� ڼ���Q�X"��;�H��`_Hz!
E)z�1<Wh���[G�\������A$NL��5B%Yu��$%�}�O���Gǐ�F�x�j��32ɔ�G�¼�*T"GD!�1���S����+�~^	*�w�l�5��"_'�P�'�)�\z|D���lHE��/޽�5�L���T�j�)�2�ڱ�j'���&��ux.{���eVi�m��e�^�_�$}3�9Û'���Sv��G2&����#�A{C2�����?�oV������PM�A��&_�q�!���0k��L�L��<��S�w]?m��|�H�⩻���<~��0#_�W* Y����j�Az���N��� y�#���6�㖰=`�k�@�(�)���:f6G��N���[�}�l�s4�� a��R7'�c���{���q���%�1uqBSg,U5�|~��ˠ��s0Uӈ҂Y*�F`�r�xL`���5i��$?�8��2��>�-�+[-3�:��3�A�ߕ$��|��Z��AK�r��h����ͫ���C���`�����3��7�,��z1e��PB>�z\t�̹mJl��Pȸr�nP:���)����*7�Ú�ͅ�ȉ�k�x�-r�A�� ����j��a�z��]�+h;>=N�nݪ}��A��>�B����cCA/9Nfyl!���D|+���7Ac~ ���ň�z�͟���)��C��TTF�4�)�S��|�d� �r&AUӛy�D
�e W]��+� ��w��	�Tϛ�s��x�|_���\':�*3t;ե$��R^<���*�YK	25��_*ڛ��&�Ur�q+�X�mc~�5+Y)GA�͔>iի�D��e��EF�+3����qC��4c26��w�z�4߉y���H�0}ϓ��������Z��T��g���j�&���~;5��e��B�w��"��L����V��|�]�L��ڵ����y
�9�l0�c����+kL�(�>/4�W�x�PH,�@�_������k-���ϔ >xe��P��1�X(�@)Y�2��Cԏ���0�[E!�Yh� ��9���\;=���8!����+�����IMօV�h���E���Z{�hfE���Z8³K��;��k>yq���A��VbK2f5tt:�W~</F��~�|�,�B�
�F�LЧ��2ӷ# �W�೗����!-���e~�xl��>�2C�n����_� ��U��u;�"��/�=��0��)�W����4ꗶ��h�Qlq\�G՘���/V�C�{�xBɤ��tj[�a�XR���UÄ��S؉Zln���>����[��E�#�[{V%1̂}M���P�QkB��� ښ�����7ݑ�G���v�{��4�Z�������`L֭����3ߛLP��J�Q����x�����e�R�qtns��֦��dS^�<�7���|(�&�VĀ�%�a�*5H�G1@+\gc�÷��@~0�EPN	h0�m�W����	���'2�m?��'vW�z�q��V�C�<���H�"\��o�5��n�I�O�����G��\��q5����t4[�����A������vr�c��"O��p���(*���#�u�([����w8:���\N5N#.����N\'ɶ�}ݚ��Xt�v?\���۪��Hv��ieM�A=��3&����PU�1�=B ��T��A7�0�車֙��,u�>���s)ҀZ�rt��7"Y�Z�ۏ{N�f
�E�ޅBsti|C�=��W�-��[AM��R��#}"6�����ٓw�����He�^���Ք��cw������o�	�A'�Bj1�;�ϟj��@T��U��W�4��� o�O��W4P�g�_���&̚�97ץnWˆ_/�,��ch{d���qJu���L���qF/JؕN�Q����'UOn�g�[$�k�:��Kӥ�6��dLC)����#E�% �G{����c�Յ_�4��� ���d����.F$$���X�ڶ�k?��C�?(/�
�"�A�����i�8p��ߌ�I��{͐��7!�m����RS�7�w%U�w�Ғ��m�;Z'�d�Ϫ�2��]Kۑ�Pq�.��v�f�tgp=�{G�5N)|�����f$�N���U���y咬0e��TOG���Ė����!3z��!���*�N���t"!�\�u�Q}�Ԫ��E��CՊ����
�,�l�4����@֮�l����uԭNT~���,�*N2aъE0arD�t�[�����������#[��T"�g�����9���y�|RFN�merf^GEYC�umjqB����^�$3�,;m#VE�[�oF�.E�j8�j��'� s��h܏C���5{�:U�2˃�� ��@ �Z' �,(�p#ė�^c��9Q��Yv��AEX���e��W7�U	]\{�K�4جΏ�$���b���0��9��\��b��֐2O��{3�� �7|�%��BD��q����%�7�Z�pq���c/�2k�ŧS+��l�9DS-�1I�r3��f�b3� �*V��*�a��+��D��ǰ鐱E_�"���ȁ#���&�'�aesj���:������s;��'|t��D����G[Q�]���̈́$�+��\��3�׬��U������,|�`v��^H��M͝ɝ?�]��`�`�g#��P��˴]6��&��$R��{���K����>}wi+D�V��5�^�:(�~~~�`�\�T/�n��_dᖜ �4n.����g�g�{�?B�a�F���,]`	/_�\Z�<S�HN�9W<7���z�u,�Mu�H}�v�A��T��C�c��N����1檁��-�?P���l"�K;�8@4$�g�i����q�/�kLҊ��s��\b����'�U��a���$B�P�ǘ�kq��.��6��������VgoIyhc�ꟘU'9#8��]��y.��`1_n��<��?c��������6��}�v�j�-���`($�p�m��6�ɱv֡k�vT�;�z�P}���u~2��֡��s��shޫl����o1cJ����r��q���;����Ͷ�ݵm͝��`�j�՘�� ��e/`e�*�>�F:}wI6��N�_�֩i�{�D�m���~�gO;�bA�:�?Y�%Ϙ,V5����Իھ���,ٵ >姺��"o�k�RIN&'w�+�Y���2|���J����W\͙?�I���0�=�ݱ�T�Oa�OݤX<�����s��T�ה�
1we�)�S�ptl#��g��2C���No���%����nI�S�pT.��O���m6=q��0H{��e%P�J�=��%�!�(��%m��eƵ�L�d����w@nV�%7�O�������P�F�ZW���]�o
Z�oH�S 3N��K�U,wbڊ�!�0B*�d���U$A^ +�D�nԫ|���uÞr/�J�_�!']f�lzD�,IA��W��8.���^h/�������|�n�H�B�@�ZB�WQM74K���Av�}Uݡ?Q�0f3��9d���O	KI	����V�����5�p4�%��x�漑h�᜻f^����DR�?n�o��&Ǩ�:&mGtN��x�!j��� �"�$���sHԩȠ���d0�2q�e9Ý!85fxS�4vܟn�m�$;;���U�����Y-�����nO���*�o�ɓ�m��i�ܠm�FU�]�
�o����xa����NMi������ӽ\��b�0���0��K��e��!�t���w�b>pJ�/U5�)s��#�M�ƥ$[�L�f��=8��E�>��d�S� �ISa.���_�ݴ6A����Dt��yV�@�t�y|:o��>n��ѩ�N�6Ԟ8��<J�s� �R���y����a`���I�{��������|��"˾�/Ж��mu3s�x��Iw�P�ߙ�E=٪ڀ2B\���A���JCDm���m}f�xC��tE�	�ꊹ6h��JS�ɃL6��s�5losO��yW�2	%�ql� �?�r��&�T8O�������!Ѭ�G��r ��L �3��]�C�|`3zA�e�T쳩��Ky:}eQ�gn�W3HΝ�?��v�Wt������/n�N��u{���.4�,��M�0��"�:�`��Q-�;�[fK�%"���A-M�"*B�fd8Q\�� ��K �}{	9�HcLzs��_� zJ�]W6���T�ͦ��a)��z�.���\�*��e�-�S��5��|���(;m� T�A=��d�i�x�[IV���;N�w��TsM�_w�����77��|;+�����>O��>�vW�9�U��=���T 򞙱�d6m��7��j�>*��&YҺ�R�h�p9j��9&�62�v���Y�dL���2R��\<��!�����0|yA�Dg=?�2��v#��Ufd�}����`��h�E�]�̂�����S�#7~3�"��%Bf�2�Ԫ�8�
��5s�Lљ�ָ�������N�|��C�@a'�b�հ> ��&J]��c��hƫ�u�x��|�����I������P>� �O�'T�<t�4��q-�L�S797�'��cQ�diY_y;y�����[�}/��ø����A�����	>��J^h���U���G8�R��*����KHLqw�`EJ����lY|��ID�T�$LcH�9�SG��c��C�wku��Sۍb�>YF/~��w�:��A��o�֯G����y&?_N��u�)��Z��I<���Ƒ�3:��pea�����K���\iM�9�9���ةbꬓ�M`����Y6l��X�M_	(����r�v�����#�|�g����u����l�c�x�3
uT,�:p�z"�����^��$�"�L�I!�l�g!�C���cX��3_I�Cd�-��rO�7 ��|�WN�I<y( յ���
.����w�Z�-Q*=��-�đ8�c����{*s&1Q�����v�L3C6��4V��jmZ�#J�Z�a7+��/�P@�	�m�D#@)�Ǐ��|2C�b�Y�N�ʥ����;��'�\�Aï�1������*fIdB��w��KV������ٕ�*ͦ4n^ˎ��<�+B��R"���%x$ l��MJ�O�t9�B�pn\���]��%���e`�u7�K���?�X#��7ݲ�4��!�7��� Oȶ��<{/�mMߊE�Rn�/֠�V���eZ�=�ѿ�2g5Q���꺍��	3Lp���l��rUf/,H��9,�.�6��HЌ~��|d�a>ږjQ�Tgv�jAK�_b6���#y�� ��U�������C�Ko�uD����/��������#0�"���S�������EqdS-��lo���%���r�W�J����q�j����m��|(ư�$�/>�z��q����_�GV��NʤQhP~���'6���'*��cEAسUwS{�Nޯ�.��I!{<��0�е�qRC��һq�("�Ezy=q_Mi|S�ʶ#��g�ɹN��}�E~���y~�7�:Ŗ���{ڎ;�3]|˗m��݄:�����g��&�|D�0�DJ% ӏ�����e<r�dr��z�J�� .w���m�;?�w�#~՘l�_7t�cv�踝X��i�U��E�ek���'�7�&I�����W�11��e�f�}�S0��8����A��z����3*�_D��L���iƵ�z.Ł�S�)�8yۭ$���@Lb����Z%��T�!R��/\�r�#��}/�v\pQG�o���v2V�2�2����v���6���kGc������ܦ%��˷� "L�n�A6c�g�Zq /���4���-R��K��n�Q�Z�X�X�nw`f0�{6��� p��Q��O�_̛�)
���q���9�*��(�fjrJ}PQ����j�Y{>����p7�]�%��H�e<ÒpR�&��MYj�V��R�:v�"1��[y�|�Ez��COԞZ���ա8to���"Z2��˻��6F��͡	��6Ƭ�aX?E����Hs�O����4iC8�t�-��(u�"��v�-�)�\� s�t*Q04_���Ok����_�@I�h�t�iTP���G))v]���;�;C�9%QL��յ���g�[6�ka?��P��j ������ٌS����Z��pg��7����p��.ˍ�2��p��6�g��Ѕq�M^b��N>P_Gno�Ku"����A�|�_�����)�m��%��a��g��e��D�n���I%��Ҿ��4��o�(�ڶ�J^و�8�NF��������3�K��3#IW$��ϑ��2�$�p�+N@U���^�&�u�#^������j��7q�t�S^�f����-^�IҡQ��k!��򹷾g}T�C)�J��CF�<AAK~}���hM�_61n>WZBT��dr�����%�-���D՜3T�`�҉�X_���QY�)�ƷA�ƻ�&<qoȁ2�Зw��!b]�� ���c#��g�m���7�^"�cX�Y_n��qځ~���an=�?6�'�	���3�^_�"�;s q�{���WeG��s����K!����~��8� :�Xނ��)�V B�����:M_�E�C�\Dsmi�|Z�ǝe�{�Px���x�3x��TK�N���F�1s�l�`Ӽ��|�5.���ڡ_�3������%K��`m�f���˴��L���従��S�-R ��w��=�~����7$�a�{?=49ߖ�6�I2:�(�Q�����3��~�7*H�j�����!Ჲ�d���ܥ/d���`(c��1��oV��2n^$��ߦ��z1}{���V��b�T}y#WbT&��&����k֦y�]J���}����-g�Ւ�s�@l�p�I�lpn=�fh�@b�r1���`����
�:|:*Wћ#����u�k�"�5I�4����ErG���}��@�Ǔ��\dp��J���s�j~ʷ�F��ʭlo�M����0�m�_�@L���`�Y�B�3�&�f	�б,=�UT��x� �`��%m����ĀQ�t��5�,tѴ�OE��\���������Rϸ�Ay��ݿ�1��Y
L��n���wq�y���A�$�X�����\k�aX��R"՘���0�������XR��P얿i���;��sL���*4RY�x��Hr�b�>XВ�:�e�����'�pqv^e��=��ˡ��1��N��l4�x��K�Mَ �z���ӎ��{U*��$�66\3CX�j�z���o������y�'�]��R<�x�S<"'ͣ:5�i�������#�	�V[iL���}:���R����E�Kƺ�ڏj�i�n�,+�N�9���}������.`�4{E��z��ٓA$�ϧ��zch3���� 1�f	�Pٜ붸m��4��ۑ�k�� �V�#�y������$�*�d�
���_K��Ő���� ��BV�U�4�!wX Da{ ���E����YH�H�!#a��%�v��)[|�|��b&���8IdR�
�=�����WՀ�|��3>N&�e=`�QL���_�a���u�5�����̄Ң_붟w2�*2�6�����ීc�R��x�I ejMI��n��I��16m5����N6�E���R47����+.���#�dW��5�mԆwz���	k���]$�D��nT���荣IU-��;��h>�?��7��q��[�(�_l#d9h�VT$>4��?���9	�o/��<�3oqGX|y�g9ݎ�`w�.��ѹСYd(Ic:�l���>(0�Y�+����u�3��=�Ar[{������yES���:����*b��ɮ�`��䋥�o��!̄ �V�d�A�����j�AF2�6EV[o%!j?�0p�{�p[%$�}�j9�H룜~v�7*��|%\ע��[Zlٯ��8��A{���(�$� WW�r?�u_V�u������X.�k���4(�[��v�d�RSo5������\�!���<�aX�kI�{��.�F� �_�H�����Vc�9�bp�{[/�9��.A|H�*)cL������N��݁;u�谓�1}�I֞AEh�z%łIb�����W	#�'�[����`�Q���N������E2KJ����FO�9��}��'��'�K>G��<�/�̘�#��<��{�K`��jڻxÝ�;U�zmj�El�s{�����)⸻�V�fs0zPI�ʰ��wpR<���j��cm:q�Z��)y֘SBJrc�[Z�t��UČ ��v��p�x�˿�"�H��J).�C�d���x�֚.CQ�t�����A+R����FB�u�sT��!0�1��)]Y:��
~[���4��Y�~��l�M�0=P��9�I	�:�ر��� �Fy]�BCpHFP����` �3x�����;i�z �'���Z�e�ʨ��#��#,�����Tݕ�6�~RYnwޒ!��~ݸ!sރ�~����}T�ig�}ZP� 
"a��������r�ʾ�����pHȀ8�ꔛ�B20�K�s52Z�5�ǡ����$�2�`���f��kKF5b�V2A��Z\��w�X��-d7T�l�ck�P+�b�Qվ'����)N4ՕLZ+�]�A�{�BA���ao˱�i����GM��8�C�n��,뗍C�� ���x?6%x}B��ma�d���B+����X���I�H��j.�T>p�|��E��;Y*�;�W�~������@ygF'��YⲞ��WȻr/���տ��q�ܹӴ~F�=xβj[�X���Ur��`?w�cIg�۪�%r��k��o�1�_�L.�,J;�z�����	�h.$��EO���;S���j=W����S������=��P �ۣ97${^�����j�o^�,z���ж���������R�+�m���?d|�-��!`|�����p�W<�@^~���q�a����ĪšL�u�lU����6%Y�"^�S]Ec8
�L;˥��ϲ�$�D����?���'b��䋲�"'4}�/@�ֽ�4�Ϩ�����q>��*���|���_��RCm��zy�UťJ"iq��͙�/t�T�|x�R#�����/{�X���&���!�b����4���2y��$�V�pMw��ùT��)ڪy��� ��ZR�ІE^�39v���~�rs�h	0(Vp�� MR��e#�|�Q��$:�n!���^��W�F��u�d%�/�N����ֽkmmO2���z�#�����>5u���r��IU5�h}��c���xs�8���+������Y�!�<�0�iM����8Od�w��@	K�&�3��������IڤHT��^�y;Fж�˭g�������P$|�_�2��,�]��i|�� e����!m�&( D��G?,*9ހ�I�7+��!�a���Y�1����(2@{�H���q��p��?{�z�Oq<0Wr���O����F��2��a)!$\�z<�%,�:T����/⏎���7��51G#���&<�F�1Ƽ�R4���l�L�w+,L3 d�
���D��<Pc�8��C���h�Y6�" ð�];F��ʿ}�/�D%�U������J�>pAz��ɼώͥ$�0���������ɸ� ��T�R���[�$����`�Р��O�t���o���|!���/f��mN3�.�'z���C ��m���
�U����\�U'뗷DӖ U�!��u����<I�I��4]+�@�+G;�3^�4�ķ!�?2�˖e���������慄�.C�l[B�J;M���Zm������B�*K{�R���ѣ:X���Z��\�5ꌒi#Db	gY���ը�ĻA�(c�A-����~�L�����q����H~����
ܑuU4��H;�q�v{-K��CV�`j~��ni`U-��Se>3��=�=�i¾�91⡀*�Zy"�$�ϥyM�l�S�|gh�*�R���ڸ�����qZA;��t�Z�6h�yv���v��/���;�[����ᚻ��T' �^�7�?�1�^�!wDp�8M��%צ�	��l}��!��R� ̌�'��^�]=���kZ%���7���T���j���ľ�H�j^���d�@��l�X����jPi���"�w�P���>QJ��[#���V�E0�3'>|@L��)�����td������u�؍�򶾭����MW���<I��ٟ���o���U�+yI�P�L)l.��n�2ᑓx.OH��m���[���9\�7G?�/]4��xhZ�M*kW{�g	Q�&����_�3{z�짦��y�z^,&�Ȓ�K����=h�>�ho��721
��A�� ˗L��e$���s�w�VUq$�rE�G{BW]\)R���N��E�ԛ��5܄z/�鹯�Ue"�;����6la,��w���ŤOz�W�k�v]���Dj~BV!���v����e�x�Vs�Nж,�F����<`h��o�k����.Y����+��%ZAa��n��?��oU�����H.�V����t�1}�E<��J��)t��N~�{��'(o�`�z:	<I2mN6�t�c��������]�8��X<�.�a��(�W��N�M�(����ui�.���jӽYK�xUܤ?W���U'9nR��288��E�O�́�������˂��|?���W������vՠD�W���E�~\=��-���	9}�u/�{}��IE��x~/}dq%B��
��ge삛��~��qLț'3 ������ϣ��A�ۼX!�Π�`�/�g#ʗUVM!�� �3wQ���S2g��|��C���u&�dS;UF��d�l#F�w���yU�MTf���y+������B/�&&�<n֦u܎1���7M�ef��KQ�t���ۡ;4�D�QC�g�o��`z�T�w�*�@k{�
O��V&�����|c�
�F0��٠�e��xA��+M1��Rߋ,x�wgg2L6��R/��;�GK�����x��&��;=���g�&iQ��c4��Ə(��"f6�)��`�����Q�[Q��}s.��G��CX�m��K�u��+�$]X������H�����e�����= @�ѵb	]��{��@�
��_7SL~H�^&�D�����9�qe����|c��aN�}\��G�V	M4;��`����8�+>k�}���u�W2������UR8�xbހ_��َ�-�QS�������Aw[8@��k;]� ^�[77�d�B��'<z�<�h_L�ª揮(�kxB���X�[�'㾬gi����"$wLA/.����Og��&5*ͳ�mD�����e	�u���<�M��勍����]]N4>�LY�K}��4Us2�j�Q���C�Z̺ļo��Vk�:l�fa�đ8P�\���޻f4���I��V�q �@�<'���49L���8�-;�X��u:��ǅ� ���s��[F�r�Q˂��lL��Z\Y$O&�y|g�q�j�Y���Yt�$d�%���D:xC$>.+��=�,���/��:��	�nz8����1S��i��X��������Ќ��"��[�r$BL�[������Fz�c��caG�M-]�B$��3��˙J�Z�w��(͌��(�%|+A��Ax���WFC�,�V;�V�6�KQ���y=	�`�
�� �)	h/�˼!�=J.p����5C��f}�o9�p�����-����dJm�+��o����%Gj2�p!�w��-۰�*��$�P5I����l�;>���),���D=߀H6uۍ�����U���_re��4������&���e�����	 �W��e���=�D���0#`�	��U�ҡԓ�H�M<�/4�ʭUhM�$j�����*�Y�/�%��� �ѦaGp3;���
g���r4	�7�$�=F������ı=�U�m�<������-:���X�JwB.�N�u��������V%T3�auO���C�F}qb,��柒���2H�����E�M�}����F���F�xF��NډS�=�B�ͯ��_a9V�&��P�ܲ�"7�%e� �ďͧdXvU���~���pRY��";��Ug	쭁�AOx� r4L�S��D�;��ӳm��|���Z�˧'��Ŝ!R�������;�r���� 1������@g-�圪Z�,<o��l��T�T��A�}c;:�<�]��p�ڧ�O[���d2vF5�os#�Y5`�0)��т�'$�W�UM�EQ�%ޒj�ՠ�f��$�^#�0���ASnG��G���g�(�BNd�R_h�V�������"��A�]��?q�<�~���8�Ĳz�U �_���xNy5���!�����"���+9=*\D�ug7qG���v������M,o�'��q_��'qe*i0A���
��~
�$h�Ɍ���%��W���Ф<���6(��+��Y����XPq�"ټX���T��
�_�$C�^�<��5J֮�~Lz���#��	�V���K���e^O�7������Ӽ��iܻ�p�DEXs!��G��ҟ>�2y�/+g��sy�Fѥ \��3�t�g���W V ����:Z��g�f�nz^
ƃT��7�ڹ7����nU���I�_����[������T�1*�T��c8{��|Co@2a>a����e&؆�����0_��4�N���$��w�)��<mh�7|	{�e���v�H���(&TxޢY�E1���O}N���A�q���mcs��XI A� ��kz)J�#������Ml�s��N=t�C�ӓ,&k)(U��`y��F��O�G��L�/t-�|c��ҩ�``�kU��=�f8��r+�P~VU�tR��\C������U�ފ7�	�d!��B�N�:'!���֜==�\�)���Qa�����[�B�6W�y��,'�㺰R�c����Ohti�p`� "�/�*��σ���Fڎ������Y�=��!�~�xU�>��E����z��`�r>�h�ʗ�<�V�����|���� � �����r��k�xp|�Ԯw �IV@�i��*],�]��4l�Bwr���{u�iiː&gSk����z�E�����44T:����5uS�Z"SLY*=�Kc�����(�����ja�Q�82O�FO��]���J�5����4)���i2*�BK�nډ�p���טv�v�i���S��%��d��MO�(O�M�ɆQX�s�E��� ;�Z��� ���ZÛJc`"�"�����v���r���)c>�zY���d+�>�����P���9 �#��Ӄ�Ɨ�̚+L�W����F���>o�A�������ϣ��#�ye۶m3L�Y�B�`i�ۮ1��w:�M^�*<k{LKX �i�(�Db��Z�~U��֓MQ�@g�����F�z���˧(Dw�>7Ѡ �8	l�t�S��n�N��K�shjP�9�'�j\�X�]�
_0
sma5�B��vL�Y�_]*�JX6<Z�7�!�7**or��`]�9���D�|����ބ#Y��x۹9*�����T"��k�j����H�f�J�D�%���뤍8�z����y�B-`�:��5KV�[�DYG\E�>U#�p,����~	p�y��|��
��εXy��T"ʱEy.����,�2�:���=�X&\P}�����t�i�=��ԀH��+�[���vo�S��Y�o6�wX��?]�lⅎ���1��Y�&�*����%Ѭ���V��珁JT�x�[R����E��(%n7hZ�i$L��.�Olr�D_�s�����==�f�U��W���,�m�o(�Cþ�K���s=xc���#�{�1;Wd�]�!���#���zQ�4���/�5	�B���bb�;�֭:,NGC@V���� 1�գ��@en�Jg�&O�+E����4��a����&���Ǩ�bc���]�_^0"!���(��p�|#y~�l)s��(����G!SfS2]F���\a�����|v�0*�s��؟�DT9��
E���DȠ	R~�����o�f%���5"�f�z=�og�{���2=}�ԃ�)����rB�g��3~J7�g`��)r�U"m�j�?�3��a�V9�-T�]vX���DZԒY_�O3Y����P�sјK��IS����z��q��YEƛ�K��ϫ̷�����`�4f��e�ŧ��hm:��&|kW�(^��1�
�Z&�D�4�^�[m�M�(��.�,2J�������U�U�U"{{騥m�s>�/qP�6���w?�_�l[���C��D���#��=���C����=�3�+C,ZC�4�CM�#Ey�Ǖ����cd\?Y�r�Х$��3$c�K	��	���i��	�@���N�N��<��&F��G
Î~G�9Ĥ��L�
����~3�A�׻Mf\�fH�.ci��t6���&���d��ꖤa|��c��5K���bN
�����q;Y����1��lFj�"%����hUtv�(ɉ�$H��eMp����El���hٱ�o�j琑KC�!Q�&πڊ�q�B���A4�͘`���`��OH5����ȿpT�1�0A�������iP����^M�I�N�	D\�6�J���R��-(���X+Z/w��hC�����-=�{M9-�C'�;L�%��c�+�U���(~)��.�L#/!�5f��g���B9-@j��r�E��~�)�hS��߆�&�����Z0�&�"��b�S��J�J8�Z�yhW���/��6a�6��Wlm*]ց�=�J�+t�0[+�\']�T��:2iK��Ϙ��6����dh���,?Z��|:/�E�O�T�Q��ܱ���}쓑�6ޘ sE��y�Q����p:�V���U��/E��Iӹ��*hTL�;e�}����,[A)��A�Bj���X?�X\�5��P�gk����x�-+�pϘ|���=�26�~�5l�&�+����,��9MfO�"s�l$Ɗno�����5�h��$���qT�Oa��u��-)�4$R"{M�3���HȡZWu�h�Zr[�Fh��_�y4�%���0�zooO_���a%/a[�.z�%�T��,�e@�n�2�|���\�@%��� W5<?2�Q
�t6(��k�N�>UHu�}o�?yq�}�%�J���t"�$��R�����e'e[P�/�� �+�d��@Ӝ����r&�s~�xD���xO���Y&��6�U:�2.�0�G������tvK=��%��F��8�V���m_U��15�ߊ�1Z��Qs��>�g��oп��E��Ӆg�X~WZK���yg@{���-ާ0�+V�]!IĴKo�`�{���k���[� �0�6OQHmc���}7��0P�W$"xD�Ȕ�DN�L�l�[1���SGn�䨊�8N�;���_pE7�⒞ٸRC��H>�]I��,R.�>��n�+�Ő�5��%P�y�J\�:����~���U�Q����x�6I��j�-�;�����7v�Ć:dmm���f+-����-�%e�{�<�j���)��6��U�!���
��Z�=��r�i'�oCj� �{���#sߵI*ysӉ���كohۄ�[�{�O�e:Q���˯aj��`2ѝbOi$��HN��+�H�;D)�� �8S80�P��O^&�r���ReU����lg���d���h?�N� ���he����y�-�ddM!�d�M8�<��_�:�H~�M�P���%ت(��
`�`vQ�O+v[M�&�#��&NX_�O�Β�R�D�	�v%:�"	߿P2�N��������%�\ƌų��L����I����-9���2�VG�x��H�^�=(L����l���sY�]e�m�M�>�y�P�]p#�фA�k�Wo[�=))1�2<�f���j]C'���ߨL�|aݏ���T���S���^}k�tW���.��R*�u���5�b��?���͆Q�����8`�%�cP���4���/v���@F��빲�NN�O�����Q���	�QwK�nM�4hR�ӻ��<�t�/�[�����f�%m���m*s	DA�{���>sZz�
�+)�T���E�Bpc�V��V���?���3	� S;q�A�ҳ����hC!�n��:����U�%l� �j|�pƜ�=4����:n���5��lN.���)�� ?c�U����TW�"c1�`�M�!ʭ_h��Q�C�t%�sȌ��'#1�a� ����pV�p7�}�4�4|�ۜ�H�;�v,�����F)J�Me2�U#�E ����J���#�.�<�kVA;�Ư�+<ֳg	n��)�<a��AM8��	%s�]��,�O:�3p�C6��(�ym��D��AnV8����o�Y�w*.S�W�^9mӞ:��-:�X�Y�@Ye�	�X��}fh�"�l��щ|8�N�@�M�k�\��rR����+�C9�^ت�l�^�&Dr)��c��l��`5<�\�쨇�ww�.�f��aD�ao5|	�}ֆ��������d]���gق���:�nR�/1o�&�!+^\b��Vݥl�����*�D�~g�Wh8���X�)B�b�ݍ�CA:�H���z��P���1��6��gi��^	��̶m@�EVؿ�VX�,A�T�ZӷnǱ��:��2�������/1�V����2]��!H�ʉ��M���O�6V�����Z��d�!��W�X, ��'urH��*f��H��wŊs��^%ۺ0�m�i����m�w���>��x��^�:!�8�&�u�X���zV�܉��`�o��k�j������:%ч�s�:�z���2e�ϓ-���Z�"�j	H@y~.i��ُ�.b�2�0�$��àt�t=.��$8@�ްGt�d�ȿ�p#8
��%��]�Z�}џi��M��N.������U���G���<r�Zޠ�q�,]�R�{k�@��O�|K�L���)�\^���[��e/���t&Y���V��ƪ˃Tm[��{�Ӌ^9ri����8:| �k7�g]E�k������_�3k�v~�&jb$jIYBO�0�Q�����\(�Y��s�c�eCE�(�_�6�	�\�ݰck0'*T[팰����HR?�B��̢I�,�R�����}��jO'i�S���C���I/�7�:*u/���z)7&?�$�E����Ӿ���Y�t'������X�G��l���E�b����Ӳ���93��k�lu@�SӇ
0��>2���S׃�ԥ*�D-�d�<ҋl,zL�\����f�s��0�K��Wy�zЌ�l��~3Ԉ�fZ�*y�I�ⴴP|D����l�^Up��b�C{��xF�V����n�$��� K���vI�^�K�Ft��Z71,Cxj?�������z�7W�[I�Z`x�%J���QL����Po�Ʃ
|,y�LZ@�AM0�l̺�d�Gi@:֜$&�p6��G�Bd]}Z�lb3q�� |��%Ӭ�@��W�7��1�� hV�9^A��1� ���z��R���ߣ����6�g2���ê�7:�r�p=��)�f9/��0--�K���y��6��=�K��-w��@�ȁ���8|���0Ѳ�hEM��45�����C-��n�1�JV[~��J���y�~ŉ�xU-������$>A�E�Z9�����H�=d�����}[0���)^R����+!+y��!�-{�j�I����z_u���2���MHa`����oМ�I`����k(X��( ׫T����XtW�/*�俳F����϶�$<�W�%���9�H���3'� ?�w�wZ{��O������W�w���}ˆ�T�pj\��@@w
�����_CA�k�Qp�#����KSa�~[�{���7����>p���1M���4�D�㕱��y���qKQ0{0�88��\p�k[pMs9��ZC'�Bۂk��H�hӂ�y�p00��4ŉ��ms_�����i�[�8�q�Ѩ�,�v�oV�i���/Vm�pakQcӒ'� ��F y�0��~v�׈����D��=�i�㊿=��tI�9�v��q���֋����Q�^�Y͗_c���Yd`,Ͼ|C�6��G
	?��+� 1a%�Q��s�-ɾ OO��y����!��	a0�=g�;2���&���MS>�{��I̒����o-kd�!�@�*�Ǆ��^O��)���\�n��H��rG��a-l�S����:��QW���$��H��><�h>��x/K�5���97�@�~��Dx,���BF��R�Im�b� ��ID��$����}sW~ֹF�.x���7��@��sb5
�k�J�+�H2��"y�aa��آ���E��iR�KZ�w.��n�#NݞYZ!��˪��q����ANp��C�>��⠾E!�� �زn�v��7D�NNp�����h���r���3�(�J����u��H'���!��1]74�C�WE>��0�'��`ˢ�9�o���b`m��Z's�� .<������ކfٮ�e�9�3�kˀ~A�\i��{�8�_��"���n����/w��ѯb�NrgY�)�0(�ȷ݁F�����K/#
���g���,�y�@�ڍ�YD�!޲n,P����i��!1�eo�r{���$?��ڎ�� ����m�P�
���߱+I���b�Eb�\��6���Vu�4��<+-w�hV����S9j�!SٱA�V<�`:p�
wY!j���̖�n\�и[ZI��vZ�l���2�T���&C����}�xE������z�D�� �Eڒ��N�$�?��Z�yU�������{��@���a1�7+���d��`�`SÞ.<�_��ך���uc��]�U$�D9��W�����j����3��E
��1
��E�=cj+{_&��	�bZ��\Ih�_꩜�B���i�H�_^%!���`�;�'dHK�k�~L[�1�U%誳^8s�DW4�́��g��v�����js��}v7w<���f�G�z�6I�k�q3�����OMc��ϰn��"�}+$O��[e�����[:�G�U�4��f#�=A~N�0��!B��ͬ��8m�w,����7T/7��T'���d��ĂE�F*"q�$C�>h�l������{�F%|� �e�֑�� Twr���J����%2>}�P�����?�}	�:��|��0]����ἤz�ڈO�(
5͇��)�v>��[�"�`��8'P��)F�=�ƽf��ա7�ڪ���\�� ��W�97ː �y�Jh�#dR�����z[P��4]cF7veFI
�5��	Pn���d����KP�F!Y��\�PvN58%w�Ir��e�\A��G6�����z���e<�����X���鼐�ܧ1ʹ�����T�dߞkI�a��F5��D�������)DOG��ny@���E�b�7r��m>b ���R�S�rO�-��@�J<�˫��! M����%Ť�v���W.�}�Ek2%�V����>�L����۝]1����k6�ݜ":�hz�=(�K�#�.J+�?���Y�k󝡷��Oq�氖�	B�N�Z�d���z<���������lZŚ�<��Q��e&.y}�@��"2l�~�����('@�\V;�As��/1����1d�����h��0����Ǯxf�A��y"}9Bɜ���~[�l�� \��� Es����x�`$RZ�C|$��g���m!|�Im�&��%d�#:�����_#%�6Q>���s��c�ܬ�¦S+j 	�'=����d��~<�j�x�x����m\fwL�C�����E��2Q�`Gm��b���t^��-�-W,ϗo:K ��G��Ⴅ���go���{8��4�s�"�S�n-DOL������Za�K��i�-@@;��Շ#�>�� j3�x!�
�/?Ju��d���=�� - a�pF3�a��9��!�06gј��|e`���/6L�_$�a0,�!��@�Z�@bN<����J8����,F	�Y�$C"x߰d�U/���D��A-����; ;�(2,i��mOI�/>�CeY���D�#�p�&� ����)9J�p�Ԯ�1�������>���J�4m��R��)����Y�N�],�j*��>�����7xm���v�I�T��C!a��{h��	3����a4+�qD �V$�V�ڧ�̝�.�{.�u��C����ٯ�v��A&���Tn� ����a��)~����H�8K%�p�b����EC�Ϲ�1)Lҵ#��k���Z}�J�W�x���9�_���b��? ��y$���ac̺�#$����AÜ��� ��1�ؼ����.?m���/� �}���b������5ǒ�te���[z�8*�X��T~3u��.�����������V�@��1�l]X����������������rz�� �-A(��)�B���W����G��ns�3��Z�}F��l��&��ȟ D�	I2� ɖo4j2<B�/��3hf�d�+_E3��Z]B��j ��<���0�������90�vh%��(SӀ*|#,H.V
X?�jl�x?��`��'10n��ծ��P���W����@50w�4�Crώ�݄�4��z��7a�ޢp�x�qU-��VӬ�柍7�	b��/�z�$_�K�pZz�}YF��,�4���L?����H`����	Xm�Q �7��}�K��GH"(�7��Z>������t����tws�:tJzIXLQS��G7�� �t��^�)s��|�go�ڬm�fO�����`��O5�Ԛ�.�i�x<��%ka򴌄��lz�D�ِ�Z�z��=�![�₮����Z�UG5�3�qfLG�t�!�8���	H��.�y�~lW{ŵ�?f񺛭cO%5S��#Y`н��l�z3����ilE�T>��Ҧ��T���A\ �(Vr�R�����NgW�n!��mWA�s�>�w��v!Lȵ#�3���!����6��D&w:)pN�G�a���Ώ�Y��t��?�� ���?W�GMҵJ���[ʭA���R�P-i�5�w��ᡑd�����Γ���Ӈfye�}ŤG��T��&#�el!�lX�|"槟�٘�/�����s�]}�Ol��1VlMn��Ә8��˻��M��ÑJ��P�]�%}3\BUa�o.���;�f�,u�Ċ�3Sٺ�֦D�wQ�Wz�T�+Ľ;,k#^�+�� i���LUU1����.�)yɷH# ���3��8�gp�Iع��`QU'{�g�l2������+�_�������?��8#Uh����������D=ct�`ѭ�������j��m<�M� �+h-}6��{���tk��.;���rw7�p͊���K��d����e�c�Vh�#ҿ�${ٔƯE��޾�7�����Z��`��X�96�y
yr��:no ��H�kψ�c�dA9ه����-�<ʵ���mJ�湘�ԝ�[���D���}������g|2�{	��>"�E��6^&����о��ꨯQ�X�>}����
��;�2�k>}��%I{9hy�"����ꛈ�l.��Ӻ�%�q~?����'� w|
>���x����.���;�/��v�,Ae�\� `�-SBK���6E].N���/܏xƎbfq����1�f��P��DόyK��-��}:��Gy��֣�SJ,�6V�eX��u� =%����OkM�
�A�2�#LKoP���5�'�����
F����tfA�[[3?��[�x�����Ƚ~o��j�X�`a��-�>=_��W��ؙW$qE��D��i�8�Sqv��S�}��>s�Mm@���5��S���:�?ϧ���Z%�O� ��ىf�Gy ��g���\gΝ��3_��k6�������.:��7Q����v�E��q�A���N5�78~s�^��y�ͺ�G���_��[�}?����Q5݃�N�בQ����31�)�����;�iAD��&"Bam�Ek���{�l����O�b�7j�.G�8cs5:���M#k�$D<]D�D�!eS%o��{O5$@
�H��|S���gU]����!��'������}�1f��W%= jЃ�aE�����X%w�'�P�NU&M%�n���,��.��쩗��WB�m����-~�z���lZD$������K���{�'��=z�_�O�L��&�d
t�F"���I�y�����%ko[:I��&w��O�:�g,�G�]�(�Y �R�Hi*��.��Ӝz�aچ�)!�M���n]������hV�(�$)#,ECL�	#c۱�N�C��|��Yeԡ��R�,FQ3>NԤÃ��X�ײ�v >H�ل��yw k�s���o�,��V0�Ʋw"yA�����	
VGM<�˺VT@!<�%&�R�U����*ww�����W�3ː�F�o��m#h2w�=�/�l�k����_�C�n��=�Ձ�	e�f�켃^|�·�򜧁��?�X�	:)�T*j�b \��x���"&���c��!/1}R鼖�58����sV�懻[����e�
���6�OU���i�e�ξ����܇�=M��~�dgۨW<N����,��o���K���o�k�1 �x��kn���0�d�j��FC��	�wK��Ì�	�QV~ E<W��G(�m��ka<�+wcK]��ˀ48�N3��E�ró �"�5�ZY|�?�>�8��7Z�|�����T$~��4��.mBm��F"��-��&LX����[c��cm[��<H'�<Ĩԥ�ϋk�m�PV�@���`���:���k�ֲ���Z�^Di�Cڿ�|+��L:�{6��Z���8a�q������9�S��\8_@��[�#we_����93���υz1�S�G�!�:��'D��C󌏨bQ
,گf]�^���*����)/��_���4ہL��OG�a8��@�����񯤔`�X����=���]ˉ����ն��G�T��^�A�6Rp��VHT�5�p�$
�s�Y�B�����!J#�@������"bhu>$Wc@l�%a������u�G�^������[����cL���{��T��F��ȫ_	�����?{�z<I-�7?��m��t��B~~��沐`��HB7e\����_jY\�1�oQ�O�;���dV���P���2�N�i;�SS�'iD��P�~�ǉz���q3��1��.�Z�<�+�O�Y�n���nB��i��xTTz��G�������Ԉ!�9�Hh���F�d �k�?$�,�\��Ǆ� J
v��񠿏2�i��~ ��yu�_��H
8�e�?>�I%�X	b�Y�ddĉcak/�zD��YQ5��U�_0'����Ĳ4m5���fB��R�&dS�YL	��"^>��SUl�W�&S�Uv	�q��R�C̷<��-�uZF麐Gsp�WX�|< �>	���M���h��ة�m9:j�@��*O��>�l�f �q��t-5���]�����#N��V����a���a�8b@�~��/f�����$Ħ� v���t�6I��' ������e���^뼦���h�jbҐƵ���������Z����WR)�9E`�q���^��νO����yꌇF�?!1���1��[P:LFd��I�v��Ww���&	�0'�� [a� ���YŘ�p�s��;^�e�gh��P*C�ki���O�d����Ef��<uI���`m��8DD��$�lO�������J�y[je��"ͮμH&�weH���b��R�i�M�x�o�#�\:k=�<���띞��T��7�@hrƟ+QZ����t5|{ښ#�`���q���u�U����߸��O�N	��V��TS�,)μ�;�g�NM�a���
��^-��i}��ޮ�	�)՘=[�-��� u��h�+��#o�3]ZP2��u���Kq�83>;�	���Ի@շ��0�+͑P�-�8�,���i3�u����y]�X�O�Y��8�Ľ����V_Z,0��
�O)6v)�ѕ-n�G�VQ`
]���(�epg�����F�jP{�C�ȑ�zN���5�1��3�A����7\헞`�n��+���z���/�����_9��4��"l@5)�ne�(�Q盢|i�H'b�
^�ڴۨ�%�G�����W���ь��c���/���]���tGgI�����ٱ��hUҡ����ح$�[WEǏy��;o8��Ϯ�v:�N����������!�H���h�W)܀�U[2�t·��՗����rĤϢ~oc�-:{È�B� �'q�e�4��(�rh�^��K#�3c�T���W�v/v��Ȱ��X�����p�����+V`��)b�0��Vq�ag��x�1���rq�:��9�u��<,��Cg8�M���]b<\Ŷ�\@�[�~:$�V:I�㱄��y8�%���Ҋ�i���ӄ&B���W�Y�J��1��-W�ŏY�/�0Y���&4{�2����J� ��.��;{>X�� �5�UA%hF��)ǂ���2�'o��-�Nx��_bו/�(�p)�l��%y�c���OfS��6>o���v�F}��FW
x�
;�w�Kzt�W%pC����� ���;��}�B��1���qi��mް9�u�H��c�<ލ>�kVLy*�]h��x�ҬHp{{�goo�pI���r�����BTl���;3L]���{lf�"�=��KK������0m�	�Q;Cȼs����l�)�Dg_�V��; rB:^8v�wc��.kݴ��7�v��e� $V���F�$��z+ʦSym�Ƴ�'��L1
L�4jS ��zC,��[��E4!����rh��������P�;^Ki����?�7t�xq�F ]�7w�6����h>���08���`��<* ���(�N�b�S�ԁy�Q�*E� �W�9b@x��좞)�F_��b �'Z���
��0�׫{B�a[;4m;W3v��E||�2��ef9_�m,,��D?�Kjr�V&�9�*0d ��ĕ';���X/�=�^�^sEXe�\\��cZ��@�|�~�k�6pEN�&~0&Y��48�-Б|�;;��� rl�C��u�D�I�i�Hɫ���������� $�ZϒVx���Ėz���	`#�1�h-���6t�A:"��$ݓ��mڕ񒬬�y�M�=�[���!2�+ƽ��x+�����l��X.ӑR0�0��9�͑K�Z��i��s�n�v��᱑�TC�7jRwRԝ0E[׏��6^�%�_QzI�h�$�v-vm:�� QM���}:;|��ϟ������=P���0ǀ(BxAwnM�ݖ��syiO-�h&���"d��'�+�N�ӊ&�����(kѷ<}&��go�с��L�M{0�P��D�r���S8G-���	2�� �֬�9扃���ѧ�Ӽ�^�s��C�t\�9���S8�Q�D����A�R�-�[t��@�y�����#�r�(���ʒ��TkPj�	�aJN�o?IHH2n�J� �ؠ���wǎQ]�
+�aXG�=5�s��Oz#"�M���>8��0t��>���O�k�%+҈��<���V�E�7\�Ag�\�@�ۅ[c�p"�L��Rħ�+�yg�!vH,�9�������C����䢂;��X��B�8Zŵ���އ8� ���3%��� mR��< Œ�@O��2��nmUW<6����}\�W�Qڳ�s1��!�j�d~]O$�^�`�i��d�}I���Ɔ8^!k��a�)�b/@���̱�'�#O�Ұ�V���a6��2cU(�{��bD��m��z�x��ӗJ��9q��i�-UeF���@�e�ƁP�8��ߐdV��@���Ƅ}U���k�htyh��y��m��uwsu�Z��<�=*|�qG�k������Y�S%U��(�j�$FFg%D�1�Г�����!KX�p���c�޷��HA����ĕ���7
ip�E&<��."�@��/��d����T�~�������A�~�`����D�4{��UPK�F+A݈���*"BTX�Xغ�4��8�lN���٘���>>��d���X=+�`@��V-��֓�w�4�5c1*���k�,�gf�����D��kC�#��U����-��ȜS�c��z	ߵUw�gQ��ڰ<$������UAU^F�4_v����#ǡ�O Ȳ�R�
~�ɽLl����	C�x}S��	�^��1t"�O�� �4�о:�EE
�4Ʃ�A����z�q��8�|�qB�����0*��PP-�RI"��%��b(W�{��u���P���BT�2���j�g�2a# �5pF�����*������ĳI�n�Zg���H*��\\^�nV=�f�^�aa�s���Q���2���u7otR#n֩�I�sn���ې3���|;�8�G�'�^�}��W�3����޴C����~���R����cHp������ڀ�h����+ۜu�o�+}Y"���~_#�:@/�����G�OG5�~
�L	�5wsFb"P%fA�½{�Ad��������=�|���U 3�ux���$�l����wp=�Vm��f�ywz��Ri%������u�-����f�2��=�<�n�+$�ɧ7���>������:�e��ċ�=��)f����6~��ʟ�d�������;3�6$A�(�v����Q�l���l��2<�j/Ӡ��@p���Q��J�
(U�zl��ɻJf�M��R�%��I�g����$���'f|�ㆍ�Y�k�
3����X�3`�	qșV{�h|�J��Y=�s����P4���I��`߅k=�ޫАWԄ�2_um����-uUy�U��+6)xD�~�j+�,K�p�&���U%�DyVB�d�%����S6�$!X�:duKm�١q&�r����M�^s�A6[�pV��&�jL"/_�E���X�����,C@�_�Ř�<6���^|L��������-q���2����^�^	����U��W��	�^~*[_оe�����\����0���ך �i�7m�g�z#��LP!� 3f:����:ڦ0�<V��%g�RYc)� |�����r�%���!4%U���1��o@�G%�^qN�t��_�?{��)�K	2�'֋����H�N��h� ��������0���R�֠� Z��^cA��E4#�X$f�5�;�h�e����"N|�qZe��:�b��oM��Ƃ��
�ٌ��kwt,ǫ�H��e��E����f�H-���k�����OO\h�S3{��S�9�PQ���i̔m\�(��D�������GiTԗ��MYꗽ��*,�uJ�������l�3��܎�1���!1��H�X��oW�������(��ZE�M|PC��{ܶQ����h�>g+��B�4_�f��e�j��	?��a�N��������]H+�r�%��-$���L�ɨ�A��5�[�P�=i�Q�����{t`�����k��M�=�/;�r�Zx��W��OƆ;{�mqu��+�)�[�˻����[�OO�s5
�[���*	��&�UH��3=z2�Do�@�}�o��QB��3�I������bG�Cick������d�s���R����Y��j�s��zG{�j�OV����`���8j�~g�^�Ӑm J��H���]=Q�E$�׼�:��V&��n͘��Q�j�.m�c�	�m�Pْ�}�3�£����k�R	i�=�06 yj�|�w6-}�>�󃆎�%u}�@���AN�ˈg�%�V�F]G{xF�;n�d"xs΂R�Z	�E&%ɇ�AMl2tA�#�;��\�YT�&��腣�A��h2Bb�A<��*�>�ߙ��Ȇ��6�Er?C��@77�77���߇X�L�ΕgsI\A�S�T�)o�r�)l��u�K£jJ�t�r�|]�I��h�7ә]����d��RIy5�� mX��C��!�G����8���9���!����|Խ�xQH'b"��|o�4,m��5H�DR�H�)��n�.�w�"��ƸE�<(��m�0�~t�� .$I(��r�/vI�����������KQ�xig���V����z�<���q?�o�5[S)�{�o�g�}<��8zK���㽢8`~�v�Ƌ@���uՀ0h�zj���l�l|�aj�&�ȟ��V���Y��3�{�PD���z��U�f�MB��9��Y����SK?/���$	Z����@k�n�D-��\=s��O���P�^[�`���A��J�jwk�Sq��d
dv��`l(6
�&�7�dѾ|d�9���ms�7nէ�Z�7�s�8���i[u8u�s� z�ĦǏ���R'�E�����~�6#�J�FTy1h���*qy(�h���Ta5}�R����y��0`D�B��fV��S��!�:ҡ'�*����i�I�_t�d>ZR��2 �D���>������(tBJX�z�_�9�웸>�V	epxWI=/:�Mo��;�ɩ�X���E
�C��vJ�)n��\��G��j��3ӳ
+�O�pEJ`�#�z����B�D��|!��u:T�13�-�|;��n	������������+�i��Zk�
}�'z�C�d���m*]%U��R��]���/l�.�-i�f���B��ZuK�|˓���T;�u;;���PkM~_�>���nO��w�83�2��̖���.z��٢
"������J�gY.��)B>�i�� ���2t�7(R�6�m���}�r�}�:EjB|;�w��
�̋d$c��)E	&ޖ�(`�"}���$�('�T��L�N J�y�Yf�
ZHF��+)i��:���c�s�q-�d�I��`b1֤�ȱ���V�)�A�I���<�X<�x���V��m2�eO�ǧ#���:������Z���t�I7geVץ�=�� L۫�ٶ�l i��80#䳃)g�^�0hF��j}�B�?������ �,��*�4�L_C*�[�LiP�LA]A�����]_��(Z��:{/r_dj1��I�3�h=�74x��d~"x*e�	6�JT ,z����S�mo@��,�)��!��vS.ӷ0�׺
�
��6�H��`q�?c^~����}P�I�-��ޚ[軝TtH� �4q4�q�3�A� ����]��w��­�BK$o�#il�4& Y�s�����߆ I�!�\�4?XB-Jv�?���'�5��\�>gY����j��ѧ�Q�.�wdYMM��9i�����vd��x�=�x-6��!���O��2��c������>��3{_X�@�'�
#S�l��D	S����A+�9[�4��lK�S~��{��\cU����.��0�ǁA�j��Q��7���GQ6�P;&��~�H4����H� Z�3�X�rż��AQ���&���!�*�/�&��ʄIZ�ű��foi:��U#ܝJTaU�����RC�l���j��������P�V<3��6Ua��E`���a������/�b��6�<,�y;U�=�U�P��X`o�_���|�@z֭�^����G�NJz$�1�<�
���� v�_��ݽ���������}����� j�5N�Η�ԔL�C�Kcj�L���/��'o*;!��! �3ym{^M-[2��_N��I΂b��ٵ7����v�
��l�ҏ���A�޹�^E��x{c����;3œ�JTH����}�j��?�����t�>�M4>�
*e�ee5��</������l�B8���r�7�`�WXfS�PN� W��Q��������Ā6|���d���ǆ������I��C��� T	&���ί�E#��{H�Cr�T�Ĝк0�����7:b���U�e��c��N�	է�0�������KH�ck��+h����vBbƎ��Y��d�"��3�s�AІ۴.O�?��l7����R�J���q�!���,t� �d�TT�E��$K�x��uh�(��N�W���b���g�m��bm^�e����N�6dU�O�?RY�m2[�_���A��,�w��a�P+����%�T�V�%�7�TQ�,V��7]ٵ���bs���nq�ݕŦ2��,��+����qN~��#�uC8??�����2R0˧�!�U�=x,
��,`�#���}����|ODH٧(Z}(��g�
�Y���]�n1���=7/�
M�Pg����Ii� �9����Qw����M�K����*�+ZI>�`0y�ܘ[���L����Nz����-`��Q��t1=���x�U�wk�3���WYY�/^����%>���
zd��nx�0~���ȬmK����n�q��PT[�Et���vn��_�8ϖ�~|V��c%��/�����#kr~�x�2C�|�i�l��`7�c�����H���`�Z��1Ǻ(k�������'.A�]ha���q��^�������I��q�g��P:�9��Pۼ�ͧؖ��J7JW銩�o��2B�� �_�e��W6%�?���#'\Mf�r@���"�^U�1�Ǩr$!M��vB�y\�qS��.��^��E�>!��x\�@�5��jnB0���m��4uX�2�Y+&��a�3�9�PgU�S+���0�~��Sq��>g����?���ꏩq�?'�?/��7�1��%��aq�JD�;*^Ptr�=��W�����X�'���'uo��ۏC������x�m^`�*ٷ��f��#{J��{�7ϵx�Vq��byd=:�����(z}i0�دAQ1�� �����ȿ����4�d�'��u�thu����aG��*�\�<ҧ�m֧X����,n��A�j��%7/q-�HT��������;6�߶8c���z��c��J��(�6h��X=q�)�.�E���Vz�3[(s<A)%�2Qh�i ��=�dk4��� ��#of�#�,���������؍������0�d�ی��&ȗ��s���ͯ��A��R��m��ؗc譱���2Cu�+�Ggф���:��@�:�<��[��bq����+I��4�ӵs08aj�JB}\�w|�9�L�5���6Pa�K^[�}�nw	+�U~�P�h3eWÙ;�l�9���5���M�cTa��z��tz{�e�r�vp�F 9=�K}�R�ӷ�-�p�"R��Ku[�4�;��X���{!�x��NH�3Pؒ,	��6�3.�E!�B$�kȀ���q�39��5T����ŶX.�*uuVա��bȜ����ב�R}�@�U��4M)���:��Zr�'�$������QO	��-.+���	��5�e�:�L�	%��c�]8^� K�nG����%����I'��U�C�2BA��}
�i�d�<���@�t��i�q
9���$Z�	I�*�!F�~�(���"Ϣ���ݭ�|��}0�X��:���\�V$��= Y��<�K��n&gg��of� ��fH�/ɇ����Rh;�K����x`�������=s9�twScl]Igﺓ`���Q��k^�l�b(�z�E�o�9�,	z@yɷNv��B\;F3o�MfZX�_r*ff��"�Z��\�NOx@��ZQ��f��`Ѽ���?�:��m���J^_�4l�1�t�}���C9WS�(������>�nW�p�;ԏU��-����	��� 1���J��h�1+�.��wT�u�jl㼁�`B��E!/-RMl:ܦw{bw]z�6���B�:p|�g�tҧ��h�S�N</���_�h^�ܓ�e�}����6]56�7}�H��`���F�!mo$ pzn��p��(N��;37��~�� �}q�/�����d^�`�(99�8y��	[ �N��f���ֹ��S�.���� GÃ�8�v���LEZF;�Q�z��3�?�^8[G�fuyU��Bby���0�֭�g��r�h�x�U��$Ȟ���!7<�]�&m����b�u����x��I���_��T��c���*����J\�|��'A3?�Ҟt�6e+�?+�E���|�MR�G .�~�A�{g�ɺ,{��/��wӉ��AD��j�4;ݲ;�`�l�����T�֤�����U��R������E�x-8���H�Q�ώr<۲��rj�w;`Z+�%�	.��'7	���^h7f�v��H�턵����3+!B��>$}�$l��;�i�;�Kbk�6�����M)`P@�$�`����f-�p����J�uYm�����9�����*3y-�*bS��yȭ����ֳ�v����S�4��ZA=�6���j�?���屇�q�*֮6ei�١�0��^a.���sXRL��f-X��2=��2E��@=ٚ|
��Y�/l��C�h�T���j������Cw�5|�.Y��
��򮩉B�5P��K�nZ1����7��V��6F�J"�1[��!�Ω_&�'Y�Kĵ�9�/���PN��-vB9�Ac-]�)�᝴Pގ%���Մ;��V��76�o�g�όU���qW2�w����6�w��#�<ɐMe6m�.e�/�^aX@��=H ����_�\��"������t"Η�z���=h�n�t;�v�¢�i���l4��/��iU��Ғ��v�=�,�44i�*��\��T��7�i{z*c@�uhi�n��h.�h�؀G���ùu-��������ů�������Uh�KUCUD]�so�U�)K�,�&�y.���G$(68-�����#�v� "m�h#xrj<�٦7SC8+�(ZP<�P[ ��@�:��PX�L �SI�9�
@N�\��>���W���k���"!3�ǭy�p�l��/�1Q���v� ��� gd���:���,&�n�vL���l��C~����qH