��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���_c='�ؙ9��2k���:cܺ{�]�=���0�>Ev����D�3��b�$��9'e�8A�$�D6:q�"%
6Or:R6wT^2T�WY{�d��%��]or��q���C�9\GpN����0����U�y�ѩ4�%y6�xfc�PX��|���T`~����T���b��Qn�Zq��ˆ/�m����G�DXOX>+�zAI.WvL�>+��)�~�g�U4��4�t�0������X�(l��:��)��S$�^bݕW�%�p�J*������W�8�q�N����[�]����=�miZ��Q~s��6���I�
��>M8�qqu�]�E� TP9דFB�u)C�����>=f�j~
f6,��g���b2.�|9�$�Q���,ʡx�N�6�g]�@��1Q���!U�U�&BE����}�	7�lk蕷���6L����D��i�#��k}x��L;&�?�����q�p�Κl�����-���p�$�}��OI�n��uֵ�qy@���^�3$y�%D4�^,�B��@��h�'{^ǽB@�ڶ���(c���)����+� ��:�$�0m�X4��T��r�vU�j�T�V�.\�ȥ�%d��Ml������aT���.�Hu���M��	��b��Ta(E�!m)Дr�w�Q�Y{v'R�'���ޟ����N��Zr`�i",p�� ��ĭהs��y����HkV�NY�7f������	_�����;�t6�_��ZK���Y,��p�kK�<���}�$���E�b�
��	m�7 j�z�68z���i� C�y��vb����\iVR�*O�צ����&��i�C���B�Tn`���V �5�`��#O�tDy+�=��v�D��9����.x��!����1$b ȁ~�|�}�z)��q-��4{}EZ��#�/Qo�s��n��j/��U���/	��0:��d9��
T�K%�.BI�,$��1]�,k����+�
�c�NTُ8c��[�~[�b���]��X.!�ZM�*%���}0�kJ�n�'#��t��������zO�?�<f�L�x�	��)2$���/��{���b�LFg�&~�F�2�?O��r�ej��
����*�۔�s	q1����@\ �#{�� �B�{/�}�͸���	B�'%:XT5Y����3�z|�h1k���b���i��ƛ5�b�s��Y��.���
�G��Ws���MP���wgje���9Ӿ+��	�����+U���>��YA)pѹ9�ņ�}��J���h�w6y!����b[B��R�תQRhO��@�7�({��H35+|1���Z�j��A^����0ϝfCbm���+�K�U�T��c�_<��`D+6����6��D�G+��	���a����T>��g��M����ak/��#)��p�= ��GKۖ��ai��S���-�ъe$mWH�FE�c��
.bfs9!�1�\��Af�G�����<`�U� �op
݄Sqbi����9w�����M�"v�vvV�Dp�PX������	wT�I�V}�V;�����d(�>YF�>��q��L��8׳��^F�8�a�^2�ԅ��e�{���A
�����\��F��}�Vײ:@P:�g�!����5�t��L�$�gݞ���y	��!�M����^/2k@טq<^�H�/8�)]�pO7*n��%*��gdɪ��eq�FMjoަ�[8��,�-/�R�ܘ�_���`������NZ6Xi,�\��q���{��u�۫�4b�P�jN4����>�|�l�_|�t�X^�u�Ue�/�~3l
P㥭�&wg�ؤbſ^��a'��3���i�º&V!�3��_^���V���`.T6X<���|�z���/2߮�A�t����ŷ���h�����Y
r)���-���Rr�66RVW�t��:X�1�����x��� ��>*0j��N$Ue��eFǣm��?�t�~����B'�[�W�<I4��H�0�f�z��1L��?���L�����K;�J�-�3vc��甍�eA�P���Ha�R�)e���9�`���DunP�� ��T�!�H		��*���C�j�ТZ$���N��f��!E�W�<��@P�0h�F�jT�{[l\�E��D��  3�_%� /�b��
�Gc�������o�Z�c�UZ�x�0T�~Qy��� �B�����X.򒆝�T>Kv�x�)_�.���O�(���WO����|k�X/�f�fLUO�4
ئ|Dʳ�Ue�'�xŬ��������
B�I��׹��NE8��^GE����t����9��g��C!/��«���h��}>�b��ײ.`�.�=y�{�ʙ��5�Iz�����u�`�/8/��N�$� <��_�:��jcsW�N���ҕ�PN���JW��!wU��B#����M�[w��-Ax<2f?]�t�H�EǛ��a��{I����.?�h�ϓ?��c�ֻ���c[�K��Y)֘^�W�ZH3#���"S�\��:�> h���ܢ��8{��r;~ <�f05B����]���6@����3#�� �T�H�����^v�#��Κ�9����q�G��IR$2q�@\5q��9�࠻s8$�0� �Qݧ����'r��w�=hQ�h:A�Te��ִ�c�X3C��]���9�"�=��������j�l�>`ȗ)_����������t׃>�{��߂�j��7P�zi��J��c�i��x���-9T�+�LD��\��&"��]�?D�[�#�0�:?�(Y����H�26�>2��X���Q���#�������|j��E��q
�qSK�U��c�:|xȻt9�W%�wQ�$�) {���#�?Ԃ^�yS�V~�ǀ�E4�G��oX&���j�o@󺊙t�1���#��Tt�&�N>Eu�A�,�l����\���m��w���\���`�� R����fw/�n�d���֗S9Qw3B���7�1,<��d�p�}�v��@H�T��y�!r�G��~z��:F蕆��2��Y�Bj��`�>��&#LEQ|%���Șu2���6i����<�����H9`k���#v��ס�P��b�.��N�qʧZ�<k�g)�۔�g��Z4����Zv�OV�S��[(��M�R���i�޵~C�'hפ�������T��Y�˕Kvn��dO�\��c�R�������KY$��YV��r}��v�;}Zu�*���c�M�K0z��a�HLkIh9��b�U��v(k���)���n��t�OGc��u[c9�{�> f(?Ұ���z ����̍����'�l'��?�oy�'�),�N��A���:�s�y?�d�.<SO�K�N���b�H�đ�P�jv�L����!7��!�S���>E����r�g��s��N��#<ݺ��0��8=����� ��:��93*V`���$��\���
�}C\��rl��M�P�C���φ5��d�#A�ٱ�}�Oe�}woM_ݕur<59#�k�m��/�#�RAV�`Z�H)��j�$�;�P����ޓ%SN��9�r���Ɩ�M�`��Ev���+#�&Y��5����ռ}�7D���1�
���3@f�Fܩ��8
�wE��s4��R=i�������+�,��s�Yڡ�5T ��IJ'HC�����@MLϐ�-029���\�g�KC0 ����Т���ؼ>��5Ŝ�i��haχ���Ȕ ��;_�����f����{=���U�����ad&�d-x� zlU�⊿���I�"�Om�N!�^�Brź e1�sЩ�����/�	��()܊Pɲ�c�0�Y�4H9.�y������D�(U�;��g]����9��z��(u��~������.B�f� o���C����]��Z�{�dHUV
�<AMB�
��0Z�����3��0� �y��!a�K��2��7K��+��gx��;��4N(��|S�\1Bx%<+����z�J3I!}���	�v�F�K��4����A!�������#�&:��ՕTtJ�{C�g ������^��fDG('�@e{�֍���$5�]4\����bAm?fi���q���9
�m��ߤ�7����n�����{U" u�smw�;%tG���RR_�}z�?x[��1��U��+�v5&s�ҜCX�z��/<��e�O�6ȥ��_|�I������wb�(Ư��4x���}r$�2�n�3��6�9)f��<�'��vJ�����P@��K�T���&W�IF#���S���|���L�d�ڨ�R
`�����/��UM����@Gut��XX���s!0r=@C�4��[�F:�}ڹ���!!�����ot����"ͳl���3	z�r������j������R�6�OB6���;�����$��c�Y��N�|��k�t��޷���
ڈ�w�u�A����^�������Yek�E�ܙ��Wr�=-q�#�GH��zO�4��Ӱ�0`'U*>^>N��0 Nv�����H�oJ~�"qH�P�#�A\��� ��8+�`�x�����1���C�<{�==nh�8m#;�%@L�b�������ՙ5>1���Jnb�+ǋ�X�!n%�}�[2��C���V��ԙg�����q�?b�/�"����#$&�5?�RMo��'Ȇ�D�$��j�񆵽oSث�Ï\��>X�6)��1�MAB��b�%~�p+�6�Α?�μP�x��I��³W~�Z���GeXj��i�R�	4����n������vXH����_�$����\��GC���%��@��r�
��\(����G�2�4g�!���(��U�ω[#���PF�U����mK�Qp$���T`��[���A�[�)�Y7q\.�ۀ��g�/V�� G��
�q�)��O�(�&Ҩ�X�(c��Fef1�ZY�T�$_"����a*��V){U��+�Tz �RK-�"!l����Q�dXF}��JX2hc`AL���r���C�������JA���f�� �љ袥#�>}���A�$=�IO-�ds:�_�	,A�a\c��̥�=#E5��HĞ�if���f�9O�%�9�?&�q�ǜ�Tߚ��v�R���g^��>/�̕��9!*$1(��._Ʀ���%�����.�f���)z��$�4`ǆђ�j��]�"���
	"?�-�I܃"��%#�P���2��a��a��l$c=
�y��$���K�f۔��0�S2xp^�-��P|�*)k�����n��(��{7��}���x�� G� P��}�ZDeC�"1 �Qĳ������q���'(}�hx�1EY݀�ޅ̿k��c��
�}M{����%�����I�A������X�-����H^`���}��]5������v}�^�b(u�G�e0��ǎn^	!�n�$W*���1X�R!�Ca���rA���v�2�D<`W�$�a6&N�:�G�֋op�~��Ǻ\�,5Py҃)\1�>�J|����]�U��Θ?pqֿ��0gt2�zs�Giy��?!G��?�H=\�7#������\��<O;|��4Xj���8,� �� �I�bܽo�aW�n���
���"���Q�yp���,���ƻ�5�F�B �:�6������+I�����$�1-jFI��"�~��{��
6�&����Z}7�Rꭎ�ĺ#�+D��'��|X�W¹�?U�d�'47�')��E/1Y%�is7l�(�L���TR�3�w����cR��*�xu������1ŭPM@�t2�n,��3��yZ�ʐ��5`�vT�Bȱ����p��p���7TZ�A�u;�uag=#���"g߯��	������;%���eE��Xy��eٌXhፎ�E�TN���?�