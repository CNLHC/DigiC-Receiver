��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���;rU������l�f\gt��]/P� n$�q��Gդ�V�/�.��TWP^�4g1��6�>�� #�z�1AM��O�p�*��/���R�뚗^Ř+.���mS�W��aʾZA1^���N(u]��x�@A��𮕜˗�rq%��gy�/m-��F�����7�NƜ�ڧ�5��:(���C%��g�zS�Z]�ߠ�4F���~���I�`s�غ����S)�6��!�ISMM��ǁ���ˊM��M�c��\�a�)QG�	�(�t�����ۨK���:��\��2Q� ƪ�ľj��F��X�q�0-g�KɪSJ�ǚ����b퍴u�?�}���[~�e@��
��"�pAG24k�?Xm9ŧ3KN�5u�0�{�裇� ��3�6�hQ_�T
6�tօ�Gh
ɚ�qP�K�&�9��k���0��v�
Į�}*���kԜ���Ay��N��(��\lOﻭ�"��#3�X�֕
W;8{`|����ɸ���D�e�Hhj�Mq[r�V�[�ֳc���F��ɯ��2b�##��Uo�c��ɩ���<��*#L*�Y�C�Ԩ+X.�U�GV,wa\Rqnt��G��cr�����)�r}�xj`_���&��H�G� \�kc�aQ �7�]5�+T�j�5̏���]l�@���P��~Y���ol_f�m��4`.���?�A{[�Y�ձ���Ox����ɚ�=S�4��>W��9��yӀoƦ�.i\7�T���%���j\��Ќ�s�.Z?8mus�O�}�uRM��.�nE�F�漛����Q96�b7��q�������h�h�}�N��P�u��Y��*�*�d��>"k�ah�QR�68�̨�����	�!�'�|'��ƪ����]�Va8�G��VA���w�@��1ilS�@[��6��/���M��4t�'���Ӵ'�b�xAj�:1a��1��t8�N�{�]���$;x�s\����R�*4�l�La�5�eS�YA������IƷ�}���3���OMp�.�����y[�"	<.ލ=��T���b}���U:<�H0�����w`|�.�7�	i����2���ӊ�W~�uJ���\�&�h���I�`&b�{���f�G�}Z)H��q�΍�Ŷ~y#����Nu�(sX/Ll�O�O����a�)&\�7��L�}�]��㖄�38��d���.>��#ɔj����{�N���c�m $M��o��Sl�B����C�������2�>s��%���
#B�W��pF����mwR*r�hxT;�(�S��[P(�'�OwRϮņ��w�V���s&�Ћ�;�?UO�mZ��D�Jv�^st���vG���]-���oSA ��b>D^���|�
>VQ+ET6���ϻN��5�s���MU���>-����l%�S�i}�^4f��_Y=��uz�l���}Z�ʚ�m�Q���.t�&)L�m������	�W�pm��W���Zh��Ƃ��'N�Jfv�>(]����[�R����N+�a���.�Y^��}��t~}�.G�I]p�k�d���[Z\��e�(�ۜ`M�>� &��]��D^�	�5p��A*f�X-�n���7��*jt5������]��L!���d����(0�I�bb����� �l�-$� ���An{�q���*d`u�r��C4S�0D�p*���������-�l�|�;'���/�w�C�5�:�H\^48Pj.��$�,�t�;%x��9��9���:�u�z|w�F'�ឯ%�sI���	� h��Hi������A�;IH ��[�dJ�	t�c!�i�G�Nx��Ǉ��6P�>6,�����0��E���,��Ť��|
�t�~�bء��Q���t�����!�.�U�cx��Ϻ��.�z�7IjI&��U�}κ��-;ޯ��d���FQ/�v9Q��s���d���'G�^bI�հUgT��k��ИA�F8RE�������� ���?QK鑼�p��B��h���\��v_�H�.��qRǧ @�v[�V|�ʆ��7�z�M�w!���LaZe�ּ�H_&�h��se�����i�+Q��2�M�F�Y����2Y�EvAQ_���o? ����L���nt�0�N��3�m�T����� i+{.J�:Ҍ��y}���(��J���i�<�tOP�,��x��`��kt,��Mh�����%���} �L�%̀b,Ł�6��Z���St�N�v�(�^ �JY�P��靪-�DM@�#&��*�V �.e9P����'|����%���y_}>x���74�ўmi�6>M`�Qۆ'o)�i�s�fX��T�YD�>���۲�'ѳ���Ȋ.�Qs'cb"\q*^4/���o\S'"Ͳ�a�+$��a�JA} ��?�[~²
4o�x#u_�2��"-���|u�$)�H�/��q��h�	J!��p�����y<��R [ٽ�'0]�SǊ�v~d���y�k)�����9�x%^ǥ��;޵Y���Pqwh }�j�������cL<];��A��]s,��%���4�*�'ԃs���=I�iÆ�"ć�u�=d���:D����k$���0ͮ�����>���R��i5xr���[N��d��SϮO'�CP	5�Z�|�Т3S�8:�n�[˒J}��a��_���`�q#�����c(�����G���B=�ֶ���|�(��I.��|�v�1�zNU��7��p�B<�^��Z�N��;_V]A��+ظՋ�@+�!O<0�4��]RԼ�]x:��,�TeߑEv�������^�^�Sj=���*t�~���g��W����x�̚���w�&2]����;�ҋ��NI�\IA���YSsl�*H'F[l_d�V6?D�^�Wa��2�~V&RӉ�7���Hh��]��ΞQ�0Q����e谂�<!��C��T��*C��Ymp�iF������Ξ�J2m���h�����Eo��O"|�w�i7�����Q�����>�׾�8���%��w,����f�Q����(af�������{8�2Ś4k�<f��J�df�h� ��[ί�oGr)�E�y���(2�>~L�R����h�P֘���y�?ĮHDB2��iе@a:P����㵵��_�d>;�S���Ya���泣#�0j��G������5=��K�.g��`F�����j�4�ؗ?COg�b�*��������ܘ.˄�h�p�d7NM���l�2,ƹ�������)�zQ���at'q��1
�s� �orIfr���[�CSȅ�k�f�?1gO��y��[�n;��u�qk.uq���Ndi-�WYnO[�֟\̊I�8u�e���Puw�������B98��eذ�rn~k;P3|�߮ɹ����c�,��rr�ȃF���x�u��!F��`66��O� G	C鿎rk��8D��8<��o .���	D��6S2d`3p3��#xm9s�������wb)t`$~�M���GE�j#�� ���v9��x��\�o�뿿��d	��W�/צV��7{��5h��Ci'�\��bc���F�i��/�d�b���Pf���� *��2��L�[��5�h����{6�w9ʡ�oX��V*Z�$� 12\X'߈�6u��_e6��m�]����'����Do�H3B�f�URt��Q~2��$�vR[U�����F\�N/�hYW�&��~��d4SL[0@
��)�+��CUY.��A���9�Ũ`^&��.��;R]�'r��>�/B��f�tA�0Ļ��,�����؉�`�G�.	�j9�f��ˈ8��.I$�~uk#��o������Cz������1c�!�xѬ�s=�_��JB�����}22T�C��+窅��b�-M���C�3���1�rgX��?�2�s��=6�T�53���\\�jR��G4�<�w�&Z��F��˚����,��,D�u �*�H���?�:�s��q&ߚ�Cw�Ǵ����]�9��&;N����ǯ<+i� ù "��,ai��+��\�Y��q��ܾ}��� �1�;�$h�z�c�鯬���!��5���Y��z��sh|ʇo�
_��������mK<b�t+����T7�l�Ak~ɷ]oT��ۓaЋ���/k%�h��1�h��eii"��V�;1d]�.�l�iń��<q�w@�F���@_�&v-��V@�b���+��}[&���;���L#��6��n^���`�Ĝ��l�i���׈�S�Hg�bs���z�E�y���\�~4���x��1� ��Z^����p4���ߊ�%��I�Q���Rg�b��R.u����}��=�9]K�Y���&/c�éh�T�W�$u?��7�~eT~8�P3���c�����f��>-XeF�2(d�ʙ
� ����Z�8�����݈!�g��Dۙ�ڜ �O�����(4���4�a'�����q1VF��B�qL�m�8k�շ'k����-�O�Rx6_j���}��OGUqU;�~�$�����Y*R��2�Ÿ���J�&C�ċ�ҧ�ŏ��"�u�L[(������J���#{���T^�û��B�����k(�<lb�*\�kp�{�ʴ^A�aP��%D���%OfH�/�B���1����?�͵J��پϓ;4�}='�</`Z�����\c��߆�eu��n-x� ҈����L�j��a�.�6E�)�n�`�+�x�^���M�"}���!����]�f��挣� F��g��/y`5T6��ފ�d���@8�w�څ)�ڡ��e��|������];�@��<z�`�FS��m��paڣ�}���LU�h�W���l��(��,��Z��X*��_�Iq*{"hW� �9q���-)a=u���e��և<��AS���b��P��I�D�:�UD��B��dZ��;/ѓm+U$��I��'�@w�)=�aJ2�u1K��%(�=�{)I��ҟ�W�#Sd����cPϝ�]����J૛�!��^׉�z�/vq�rZ�������m��Vα��H�x$h�,��?�5��;&��A��A����@M�m�Cb��	3����yF��	V[$~oNΊѴ~� �g��#��M��K ��>��'�z,������n��TS
ȸE����k�0T�X�|2�imGX�e#�q�0�~Ѣ�t>v'�D��E�(�>-Q��E����'�r��F�J�~�CLN���;���F䘄��K���nJ�U�m�2Qc1��|0LQ���<���\y�8i��?Μ�P��[3(3UO�k+�1�[iy
��T2<LPK�!1z׿�Y�xų�y�ӂ����A���ZBCpy]�<�m��ح��!�������fb�͆D�3]��}��CN����S�d�#��D�4_����i�-#ܾ��z�~������>��f@s��!|\���9*�u�H�xܕ��i���$E�B��yѷ�sio�Km'=�ɍ���)��Z�����k�(�62keo(=^��ϊ<N8���5}�|�
�Y9��C����'�"���^� d�Fľ�23<��ᕖ���Ԅ��N|	(ou��)�����n�P��A	�g�Э��&P�LV�v%=R�3�M�ڻ��=L(�D���a�0�p6J���1��k9�RS[����
\�6��*�\j(S��K�bh�%����fX����}��m�I��^ea��P�C��hL���Ie�����i��N	�Ӱ�a1S���W�9�$��w�<�$�+�ـv��I�l�6d�w�1�K�yh�W�<:���Ic�z_���0Y1��ެ��Q�-�}��%��*M�^�����o�8����v����
0���.��!8��sH)�T�tF�ox>���fv}�n�����d���ښB��=���:Mt��X�����Ë'fN��ˠg5SJ~ �0E�%��4ؕ�r0�jF���i���GsXf�+����,v���9崕��6�g�d�秈����Ϛo��B��`���4�}uĕ�(,	�m��Y�2�o���Lv2|�	�B��)�[e1�g�ܒ�hp�8FZԜ�w��v0�z��f�\�_#� �?�6��";�DP��!��>�ݑe<��U%G|ʬ��nN2Uۙ�Y�c�ˬ/��Q���T5�]��}���z)X�3Z����x!{푬�3��`��j[Ւ�
������Ibh�O�!H�#>������qo��?�!{�MULa�cm#9C�"0ԲC����?h�=�@��c1#C"r����S'R߲����Ih� ;���4�!��&�+��,�����!�d��Ӣ�:��N�m�K�T�AJ�̞V�=>����ڜ0zF0�Gk&�|l�V��_��1�H��p>�_�<
"bI�F�e׻Ջ��)��N���/� Do��k|~��B�[�� ��H�����H� I������j�������ic"*iȀ��3��i6�"��I��9<������g�;���-�Aobl./�� �]�2ש��_�_��*C�R1��u�S�� t9��6Rv��\.M����ck�o�"������_J" X8�%u��u�9�A^7QFO:�'���0���<��ip�[�:݋�c���!�(�k�D�v��\*WR����>�	��&������n��j�r$�ۘ��
RPUj���g�t]U�'��y�n�L�Y����D��D�ē�q#�y��$5��$e����K�?���o`8PJ��9Ś���Ka�v]� l����8��MF�ڤ��O�C������XH�l�bXgiG�w�	�_P���6�����|z�$1�
A!����.�t�8Y�ʸ�Q-.�׋�� �7,9�Y��]�z�;]r��� g�2�ۦ���ύ�)m����V��u �
�^%EL -:��\� �0�%�}➥�ԈV�fQ'h�Z��Y����!jL2�H�oSs��F'E�q6���c�v��c��w�P����E�"&����<�g@�!�}�� �oJx
�?���>�ppi������qq��F�˟V��������i��{�R�ԧN��.�����\ۻ2v�*$a#L��6�o��Y<' .n�N�:��ƈ��w'x�}��䔁6�}�*��f]݀��92P�+�'��0��T��������P���->s�$V-@_���������R{!���)6iL��h�cy���Wk��6V_B���>��'Q�PL�&PJ�d�"54g��=Q>���F�bف�*w�gn���p���.�;�_ ���*P0�� �h����+X�V���UZF��d/�d�!��@蟛���4��N�2�\�wa�K���5�����,�1��k�3zG�c,_6w�����6��_}Ȼ�Hd��ɭ��@j�Y4��m�4���J3��q[��/����.Pl�Γ'j;��P��\ѥ�}�*����d�����g4s�V^E�2�v�aе~�֔�fLͮ���Pb��L�����#����xC'oނt�>�1�F���dy7 ZG��zVE�L�	`pt��P.󤗗���A���ԅqn�����v�үʈߘ�������M���52Ԩͩ�Հ�m#�Wk:3�簿�`���Q�l�K��b�#��l}r���N�*�Vo��~v������.�:�J�>��C,q/�0dw�L�F���>�>-��X+œ6�{s��.g�Ed������-ޛ�&y{=�x|_��_壅��c��!�"h�����p ��ig߬�3d�FM��:[�^NS_d��~�i��0,˯Q�}x�X�>�q���ZS��a���U]Ϊ�U���!����W*z�F��
�c�%fJD�O������k��K���տ ��#*�HO�2���%�\�����:gr�\~7���o���A���zzJ�>N?���$3h��|���c�X�,J\n�T��?%�Ҭ���U[N�h͆�)X\Og�:��
��}�R�A�/��Jg���	"��w/*s@�{�*��lV"�z�FG�[,w%]�c5�gqc�QËM6D8���k�g�S��T���rN�awV���d���Y'�¤w�Y	�<�n�E?��9�
�.0%P՜�Hz���_HIRoN�C=����,͂�N��P[}���7=�C�@+>4��;�FD�yA��Xg��C=&��
�y��?������ï� �ߤ���Sa$&'Z��	��%f��H�:wd���<j�/�֬��|���Y��ծj�Gn4a;ښ�t�	s�e��Z�P.��KL҈:�Y����Aj����?�XmG(|	����L�PII����$�XE������-؃��m�H"�(��8�x��_�Ϝ�Vf)"\w���WΏ���*4I%��5��{߱4����JIk&4��$oeF��}��(^�P9'2I%�!K$[�I��(� ���w���ܘv��,�|��V|�&��<������x��LvOOɵ�W^��k��G�����d�"�s���Ii���k:C<�wx����LoP��(%�my�(�p��h���9�,�K������ l� �:nn$b�߁I&��̀FJ,0`IK�T���*g���'�	�.�5���;�����)�c�
E]��$C���I�JƿX�8�B�Ja׮����I�?d��#�3C� 3�7n�1�j�c#]7I^4�%����Mԇ\����>��W��l�a���[��SQڋ�=��|����
Є"��M�'L��N����$L����e�Plf� #�v$�#���Z\�q���A�8h��0��ү����N\�濮�9C�T���cpM��V�7� �����t��3��"+��
��N���(�q�Ѱ�e��h�i�8���JZX����e��z��KK �ݘ%ڐe~-QJ�������37Q2dC
�a���,T�Y�|�×��]��P���_ʋ"U��!���c�'�����*)6
���f�������[jf��n��ש5��7-�aG*��RADr�˙!-���JisAjk��C�`��� N8��c��6����g��tMŗ.'�M�֞�r}�����}mC��d�RV*;�:�R���ְ0�7x�,��NP�m�%�k[����t�Q|�A-���'$ʉ~�p�v,@�[:7���AT��;���v6d~���?�v��L�����M�0� eo�?&K�Y��t6����oxcw@ �/7�,ԳA0�~���q���*����\[����ʾ&�q�ޒ)4<]�����˂B�'?Q�|.��������	L]�� S>o�"&���\���*�u���d$1�0L�5��3i^K�lB$8�770WgQ�z��(j����)�a�oj�m���+A`c���X-��T��,�G�9��U�x<�g7%����\$�1�7��ŷ��i(X���I
�v�n��D�5t`�Gqx���$D'�Hh&�<��|to�'i�t���!j�w�^�f
������v�1�n��!q�\�{����g͍�M�4ڷ[*?̱�G�_i�&�v��{ck4_Zpf�j�W�He�L�+��q�a����/!
)X���"�1.�+p��C�
a�{��ځ�!gX��,Y=�(}������UP�c;WK��D�	V�� :��/�R+�Y�b���(��+�.�:��C.@�<(#go�C&+���Q�X"(o��;x��.���M��#A(D,lWk��ac��3hw���}���z����W���_ʺTȱ�Aw3�lO(l��L���?�����Ê�j�]Pn��·!�-~�FѨx�CU��R�!����|�WE��R:��H�_�JS�ڞ��/.��nw��b ����c��)��'�g�St�.'�Qp�����hx�8Z��j����T�'�o������g5g\��^���t"��S�_�Y�䂷|ڽ�{)����;F�_#���r����K�]�J�}u� 8� 2w�a ���n��u�᎔7k��e<��%�MR�όbv�'틳�,�=��ޭD��U��<ы�͖n�Ҩ��'�7�2@ʰ.��U�cI$��m���7��c��~���:� �ƥ������ �`���%*���~t`���qrSue�HM<;Oq���cR���0��n�	כ��;C$���vj��i�&R�����֣>�iR�/���4*��S��8�3�/I({���)#��,�r/��O�	)���Aӕ��^U��W2����9a
'�Kأ�S�X�_ukH���ي���Hl�#�S��B�4�/���{�v'&�n�E�|�قf�
��vE�z�3�%Y�vz�"-ĕEs�v�f���r��� ��8��38�v�4�}���e�Y8N�BW��|�����%7��QZDb��6i�7=Pg�i/s>�M~Ҭ/����q~�W	��>n�.�����ɱɰ]za���,�%:�~��0��(��mɣ���ߚ��U<bU;�fq{�l@��Es��6$��q��%5�Q{���9y�psW��e��S�����B�ŤH[�R�t���ϝ/��val�6�
w�H��=�gͨ�A�Ԝ�H�xĴˇLH���8l\b�y��(���R|GD=xؾ��U�9���>C�A�1�p޺2��>��+R�W=U�B��X$b���o���qǮ6��=Z�������~�P��q)�g~h|Wa�/�� Z �K��:H���1_�̨E���>^���}�V5i�z��0Du@X��gz�#��Ăۿ��"l���(�Pa��n�ߘv�-쾮Ĺc:K�Dɩ!1��[+F-�QR�Յ��F����+�d�2gH��֦/�J�U��Tބ�I=A����$+�g�PB�����$�XFle���l�U�S�P ���3�Te��M�ѝ��\#��ұFJ����,��ὅ^{�����E	|w�JO���6�+E=M.�4'��0��<��
q������>o4le���O��\��P�:��]�w��r�M){Ml�s���7��%P<Nڜ��|��nزg��z����w@
�_�КP�0��m�	��ʯ�'�Lfn���(�s�Î���o6CZ�q�zԟ�����W�����$x�LR�5`��K����:\2��_7J�^�BT�kZ�t���ڪ/���b��s�V)L"�^��`��/�[�r��#�B���`������HH���=ʨ�*`)�ޠ��*Jw����&���9�Y��]��\�rz�
��D�����?�)�
��	Z��{ҭL_nޞlY�ѵ����x|B����ފr���,�?K��`�E�K��c�[�C�i7��	�1��B"Egh?EfqU>(�A+�B{R 2����|�O��D�@1��Y��hZ?��Sl�$7S�&#��*�y;#�w�G�6�|H,rE�7a�?��¸--��9�/;j~O���Kw1��SMM�f����	�oB\rr�A2�_A��E�:9�$�=4����f���f%^�lzo㱙�)��2��ӗP�g��K�[������q�xv
���B�̘���I��^�VY�����d��a)�R�0�^a�&����I��/��F;���i:����;K���l����M��D)�`~�&/�>�}w~h��T���M���0#Eq��R�7��|�ң��O���%�r��A�XB��T�L�f�$dEg�ɜKܓ�о�ˊi"�����P�-���[�u<p��f6�E�N�,�Fٓ��%-���òJ��?��Ǔ5�s�`a��Y9M�}��d�eC0�����m�2��6�g�~H�x_��x���ہJ{wkܺM��C6F���"zz�G��Q���+�D����g��NB�:��S<��T���k�����i�wWD���J#e�eS,4�_��;�K9�3^�����ITB�j��'��i)V�����Z��2���
���:�^��}ٔ�Ғ�e ��O>Ph�aF��\<�:8��H&����2�1x%����'y�rq�1z�G�Q�����5��^d9�(�ϩ��O���h�d���^�o�P ��H(��I�{����i�( Ö�P�� o܅sXլ��+J98��ٹG0y�b^T.M�0�ˠ�����~��%��<[�Xy
$�@���aB���`����?�}�W8����zC�����G����ޯa��&��n�I��	<�=Ӗ��>����Q\E��k�T,ݭI�3��ƛ�}�

�����NgzD�6E=����S<%Z�E�� ~ўy���}�%;��AwT���cM��v��WrF?چ��*�6�<�&�{I�1e��r��&O��r��j�HmI��wh�j����v뻥+��nhQ>�IJ�z=�P���ߞ���y���
V�^�Ƞ������|.��P�V	Y�"���%k !�:��X(�j��=��ܬ[�������#�Π�`	����v�W �������E�㪼�l�P y��g�ɱI(u��Ӝ��w�0��)�|V;�1�;� 4�9�C�\z+�b>�"�'�N@w�SL�\(���ۙ&��D"�%�l(B�V8O��o��4�Pb��a�x�)�~C�I�a&LW��W�},.���<�*vhfm�[)B��s��
��p j>�:>R0��(w	cϑе�`�W�fyWn2$����|L1��b&
?��W���}�@�e����%#��'7�+P[Rx�$�ܝ}�u=�Ɔ�ȴ���x�Zo�S���i޽��U	J-��)ʼ�X�V�oM�eB�3�0(�
	OS�]���]DM!�� ɖ�B���c*#ٓ��8����NX�(CRZ����f�Q��9/�TC9��~ީ�DZ�D�,^,��V�G���<���E��>�Ѥfsj�X�@�[x#IS��#��//$�-�5Ya�I�\���`"��}����D�(h���Pe�� 9�<��Vf}sӧN�^��:ޡ���%�#�� ^�o�	΀�Q/���@S@����;~�wm�yxe���%t��ʕ�VQ>a�o�s;R�UWF��!xL�]�ss�@��q3�;�e�x:ei��$��ah�ۄ��=��@���_zU�<>i�2~Ps������U�~�R�K�e���į�	Sz}�9���jaT��@�"	��SU�Az�?���p�	�H�d�9KCq_��:�f�71}���;p3mJ3>fi����,z�h�v���wu��G4����8��_/�RHI\��*�˵SC�4�F��\��ĚHq�FP�>�f��Y�~�k���Ed>Å�|��y�h*|�՛�{���s���{��!v��[�W�xzQ��6-0��&�^m��I���BA؍�h�7**����5Gl^0�J�IZ@n:�Bj0����	|�.9= d�ٿ@Z�B��|s|����9ƣew4P �����KĶ��j:��W�H�(�.~��;uDKp�����6��
��=2���4��m�q��cv4��� !��@+v�S���K;��>n%'�ϊ�/ �{�CEu��������3�]��y�ƭ��~��y\~�o"�ClԸI�g�k:�C�&��y���4�#vMV���f�x�a�����$��B���'{�F��ABEO�u�B�xP�����[l��+�,��1ޟ���2���HQ�\
��B�׫
���;8pL���B�p܃J��<����D�5��FD_�z��)��*%^LVn�K�W�u��$�4
�ɺ�9���0"�!�)�v .C��_�T��ZS��|��וm�u b�ե�Cy��as*�p�o�F����ׄ3��|.%�~�<	-���X�����ρu�og[	�F���WU��N��hSfkh�-��:����wM|���J$>�� �p�Gf�w-C�fr�o��c3��C9߉'�G5�9�+�N~,�|ള&󏦴�W
@%Z^:=&e��uz����Jh+s����/M̌Wc"۶���ޟ-ቈUeg����Iw��\e�}����.3U���,�׎���\���̤��ZzU3��!��Ns(h�1i C$��Ь� �����$���w��1��J�2P��}��W�s92�ERR,Y�J��?J�w���ݶN��, ����fCyZUBi�J�Ǵ�7�^ʌ#E{A������#Í�ܺ����{6?�;�K7AN���	���Zة�q��w}�K���5�G`D��9�-<'r�Kȗ@��/��N�-�k��~�0eOc�%U0{�HU�Z$o&/���Q��~�=Fa�3Ţ8�8L�o* �I�Ǥ�X�L����!�'s�*2�g����[�N�3�Xq��?��J�cu��1�w����Zy�����?�����g�R���a����*��r� ��ֶr�ɑ�j��4 �����
2;qQZ�v��w���=BFA�Ót�-Q^L6&fT����k��d/ݤ��^�{�A�=�drT�N�R+����q�ϻ���@����aӋ��rhQ���X����o�y��C1]r�۵#G��m��V3)�M/3�gD��	��< 6 9����\����3#T���oD©{C�1��i��*��T�~x�H�+�����e]LG3(���q�����/uA����ܘ&�%�i7 �$o�en�����Dn�8#Jr� ����j���}�@{B���^�-äe�g]o'��/�Iy)�F����
���Nڇ�����׆]�YO�i����^[;LFc��q^�m�����s��S6���3�'T�d�����e������JYs��֌<ˣ���qx�����-:0,��lvQ�g��=Z+ʣ��L�m�D֋So�NLKu�W�姑3�.F#<�<���@�/�ñ#1O�zJv��?���nG
�s��[�J���}	r��";���Ţ��b�P�ZLC�w|!��0��Kn�V�c\���ʕr�J�q����ܪ!y��ZsǞ��V��~��j��,�н=���i;���^?� bV���l�~Ւ�� �	Յ�ԓ@�L�W������́x��S纇�Mp����;�v%M_4�
r_�z��%O�D������A��� ��8 ��l�p鳖�۩��T=��_����`M8G��[���Rb���siNQ�6�}^C��b�9vHQ��=�����"|�|݆&R�T�Ry���Õ4`ȷ?�%��.�C����o�?���'{��K���8�݄'9S	��eĳ�Ua��{���T�����3Ǘ�����dT{,�0�1�n#!@_�"�s�v����?�y!��x�4����T|�l�B�_��v���6�r=��7�];�ٌH��ر��q��|�2{��T	��!3uҍ  RQU�,o9
����MY��+Ɋp�eH��V><Y�{`�@�h��u�Ƿu��#Y:L-S4|pUYê��o4��[!��g��u]��y��aw��"P����l��t�Z��Fǆ��e����w�ܣp��"t�c8}�tL��e��w�|m~�Ki�w�x�PQIw3b�\`w�=���ΰ�� ��;��TW+�j'���p����ĉ�P^u�4|-���ny��[�DKT���19����7�`���w���Io9�����C|��Ͽ��ĝ�d�	IC�^�Y�P��?���ͧ�@��ٱgt~�Q�i�I��� ��WLb2S=�K��57�1�؇�x"Y^�����}�O%�'�/�mS#����t�~�����Ex�=�����YL���h�����I�.a�j.muq�K����?����z�\��oO������D�ʪ+e�ʞ��>�a�#�
v��R�� ?6cϐ"��"J6�{�d�X6�r?�C~�ƴ��z���J�"KRI�7ɗ����=H�3w����F!�-=P]��>�t� �-w!V�C����d �Z�Z|�,�t�KK|)ZU0/ci�|`�l`l�SR��:Nf U��1��c�s�E�ސˮ/�Vm�#��i{�71x�S�F���+B	3� F����Ԗ˷�����w�l��*��=)|�[��Z�p_o��BW�t�8eF驅�f�1��������.I���k%����P�� �������4�M�X���Պ�w�l��J�E�xՓd�5I+Z�o��P�VU#`��E�e2K���#i�E�wx��A ��O�6�~7�V�H�7�P)��@����ԃ*	W�
k@z2�L���7����H�H�k������و(P���
��\x��Ń�t�����>�(t�A�����x'��c��N�D�?�6��no�_�u��ߐV@���BU� S���8v�-Υ�uj�-�I�/�"W�P�a'
5�7�=�������lu�k�(��o��y�3�� 5��S0v�hP���:�O��]b�`<,��|g:93������G��0�Ìk���x�+�}o���
A�����T8�f�=X�EKY#)jHW� ݐ��������L��y炻Y_�R*�,�O��/�A�Cm�vP(&}���M�?h|����v�n�M0� }��h>�Z,=ҙ��tpԚ?\f����	��>^K�z!6h�o�]z|�|֠�a&� X�Rd�muv��$=�F �>������jl�{�/��[�N�8����K͎y��vZ ��+��2�@D�v� �.s:����Fs���[�ݑ)����*�{;��/�8�7�f3x�=�x��8���~�|59@�N��9G��X`�+�͑�K�0�Ń�$�=��4�I�KҒ(�K�g��,4���/\Nl�wx/V�b�x���\Pޗv���w7�%z�@��χ����f;n�sN� I3�c�I#�����v���ۉ���%�fr;�k�r�w|Z�m��9?5�|��a����f�]v��QC`��E`oq,I�0#':<���7��Wpze���kSP��+�ܜ�t�{Y���!0*���K����4q)
�ݾkʲ���VW�z���#��K!DD��v�JW4�K���,{�$�b��ҳ�ӂ��Q���q���&�H�<{��!+�e�֎��@!�;z䩄v\�A�O:8�1����[�	��bJ��[,
��c�9H�il;�.�91ߪw|���Q����R`�
c|[ أ�J��w�N��q�c���-F	n?=�^���f��T��S���u���h*x(i��b_�|�+�
�|>&�l�ys��O|@)N��] ��rŷ�����h�m���+[������l R:�p��Բ*,��9`�3a�ֲ�&YpV�X�&�7s��SR`��pZ��'�:�4��b���툖cݎ�0��֬*"�d�{`�j_�m�+��g)����)�h,��SU�t F1ܻW�k	�NrM�)xB�V�H�x;�s����
�����[؂�,>ix�^�1Yp��ڙ��a���<a��N$g�'V�0[�%����d�<ΛD��Z1��My{�u�#����4���UAn/ADT�)�xC���@���[��������Н�'h-.ÙD�4�@����q{WEPAl��}���?�[�	ג����	s"�aOڲt�ׯ�%����ƐL��F*��)�� �8j�h�<�Gӈ�<��W��h����BM�x�P""6�*~���c*���"�L��9}�뽈"���H��,S� H�%{�k�� �������D�2�����(�6;�F?_%� ���>��T�m;FI�_�m&!u䒲1�Q{
~�@�/���,��'`�_�g�T�;����y�n����XjضD�E�0��u�(g�2���hW>_�Ȱ�P�d��<���5Z��O�6./�]M���H����^�ؖ�g�:.Նe��sWO�B�8a�1q�ي�39��|�S.��յި��V`ﾁB�k�V�|[�ab�$<_���[������Dh@*صm���l�d�0n��h��~���xr�;~�?�N���<.�*jm� �X �S�����_C��6`�nM��H�	RMS.�����.֝!�|3���Gܔ?iy����'��Jl�;r"�������;F>h��z>�
���&�J%��2L۽94!t� �M�ǹ)���IU�L�5挎�W|��9�{Ĳ%�I�P1���=2s�k�jaHDx�m���3 �s��(�����OJ<�j��f<�]&�k���,�1�g�j$�٭.G>�����mV�j ��^��JFjl�:�$�_�3�2��:�>�5M���7�$��;>���a�}�E6$_�rmd��e�q�Mbq��zwǁv�BKyzY!�A��S���NF�1
�u�
B���niւ��P� �w�D�����6� IfiFSc�l����'!�z�k�8!��&��y��6ɋ���dC�]��_���α�РpL��c�n�)
ϟe�	���|a�r���%�/D�"t�k\ϻ���A���*b�,U��t*����x�ռtV@/�IJˎbJ� ����;g�)���l}�5R�8��@��S�4:����#�h�s�;v��nK5C��]������nZ�L�&]�"s�4;D�3���ߐF�$d�UR�^�)�hH|��g���5� 6w�z_�Wv�
'L��`�!�yaiϪ��0������H꩔��[q�#6AY��X�mY��\�{pߐ(�X��[a�&yʼ�)�Q\�zڹ�y�ʽ6����?m��PC�vH�2͞z�:y�R'-�N	�u3�����\~^�G��#�(�,�:'����������[f�G5-��uTd�.���HѠ\��/3���S����ݲP�)@b !R����`���܃-�n����.���/�evH�
Z���6aM�WOv���ǜb-��C�YYX4b9{�nC����W�p��`���G!�i�����溠�'ڬ�JjZ$�ڈ-� �� `^h���E�6C-���n���9V��\�P6�h:��Ɂ��m>��~�qs���|�7�1�@aTu��Ó<"
M�}A��h�IfL���k�͛��e���
xj`s%�`��d�~
Mj�%������ϲy�f�i�
�9O/�vG����������2��'��P Z������$�k{�D8��y�K077��J*���gV
^��+f�^�=����(������j��(��N�);�d�����-�ca�ԔA������%�&tgHc���?��Zv"y�����WB>)~��Wn�D��K�?��O�vk��Ox��3�h���k(���lis��b��Q�٠�~W���d7m��'=�Z@�6N����j��V��V{�ڪ���2��D��m��yD|�]B�ql��2� Tǂ_������mYx���W<q`����ח�F̓��/�i�Ա
T �r5�K	��B��2a_�/��[�����,��)�`�D8��ڣ����Y({���}p6}�VOR'�<�h����݊�"��T��8	�G���2��3k��;�ç*�b����r��H�([�E(�O�^�[�Ͻ�S
�MϢ��>D�/�(���F��(Yp�*���04s��G\g�,���5��s�8/�"�^H~�_t��wδY1ҙ4�Pd��W�;�i药9��S��(��1�h�9���#5}�:F�;]i*>��v&\�I����[^d:������[�Y�g�S�IxӨ�)!ޜ?�Ӗ�B��mm]f�
�wFA������>2@���u!���7$
4YZp@o_j3� �Z9]�B�5�-�o������q�z��vuf��.nPW�3F]�P�ib��(�K����>��3Z���_��4bwٍ(u�� ����܈�*p����q(�*�\�@3k·�NP�jܫ��e+2�����pl��:[(D\8��x�[�R����'G�ƍ�:n�Hs��֚��=�ɯ :��%R�G�$8C��TV�����S�>�4�+H�z�l>�^,��c��(!�o��3�OR=P�ÎR�!� ���{L-�8�^�,��8�͸+�5:�a�Ըdti��eد@�W��6���r�=C�'����E�t��8q�S�4e)AR�BN��D=6(��	�f?�$��G*����_�O�#_q����Gq��{XK�BN����8ߛ��Vڙ�L���w~���df&	�j�$��Ʀ�_�_{���9y��L��z����-1����-09����[� 4��Lb�;�Ε�G�]�� �?�����{��3�Cg^�"��ᛥ�-�qT,~��C>�Q�5.��-�_��o�=����M��� ���UL�T�P.R��9^��U����v5��s({'Rcs�:����� [�d�n?�¦�K�ϫY�������2�ډ�����rG�&�s�}Pr{�<�F:�[�S�)yz�ѩE�O!^��q�j тX�u��h�_(�_2��E��U��� �S�����k�]]W�~�������bͦ�"�dJHN�t
��	r��Cb�2E�`��M��aC�H�6w#�j��Q�sޒ�~��^4�ͼ-iƬ�l'�1�d4ƯēkS⥎����\vz%v6��l#��(L|$���+Z3���Vh�-���[N�j֮��.(�4R�d�Z���[%�]�5L�x��!ZL���;��ެ��g�΅=��H���J�5f`��k�3ܭ�Y]O�^v~��-���m���)�\��
y����ѵ�c�� 1}�\sV���_F!�P���YEt"Jǘ�ɔ\��2�ˀ���_�Zh�ܶ�l-F�Ϳ�1�[��7��N0�-�|�,�;�X56H�ZY?�Yb\��uԅ�xH�QMK,V����!*#�s�k;�nd�����}�5��Ɐs�k�Ǒ<�.��j+�Y��Ί�v��:Q�h��K�M��R�3 ��*�č��n\�W��?�އqI7�b$X���2t�ޗ��6�i����b,5��x�|�,G�e�c���w�y�v������ Q��o���,�nM2bm�Y�;���qi����o����!�|Tro��$���A{�ȵfy�D�pֽr��(��7�����Ѐ��O���8�w�c���;����ቼ<�Z:F鳲|���If ��H�]�R5�O���_��_�8���j�[�[����&�D�ӛ#�=�O���2PgoPcr�[l��Dp�)g(B�x%Ix�Z����)�(:�ސ��GU`u:�"PU4���3�=�R8��:����r ��}��yͣ�{ῠȨ �7fO��7���t��ۚ���lC�C#�~�0?���>f��?�2���ڴI��y8hQc3F!#�!E�_x���*�V��ه��s	�G�	\��~!u.z��L��b�^Ⱥ
��y\Z�*�	�M�bS�X����ˤ��o��9�Yo��V(��R�	Q�,�n��hZ����Dd�5i����hXD4�w�N����L.W��' ��B�m~�S��Z��RY<�98�`����T,�Aƨ�IL-���Y�I_��9�7@{p��L�>({�J��W���[S��� �b�Eצ������0�Tl�+Ss�>oSTZ�΃�����>�o
q9om���W��$k~=��!���~ݟ{~��q��D�9듚���.@#��a��"��'bw5Mg�\��S�c<gES��w�Q~n�e(9AHᑰ]�3�:琂!����-k&pu�z�i&�DŔ*�1b,L��A�v�I�^�n�fo�{�m��H"ʧ}�<j�v����2�p�"��-��TC%cӓ+΅2$;�[�EI���',v�A���cn̽��іB�p�I��q,,�䚏T�C֘$9����.r$��B��@3�ʦ�⠋���RLe8Ҏ��4	o
��Z�V7�O�3�����e��ă�m���z�t�t��h]��X�:m�.�+�F�i.�;[���4��6L��r}�Fik������K�3�l	M-ܐ?�h�	�Dߎ�BF���e)v�fN��wI�]�WK��2L㴠���F^��]�n��r���q��`��'A1�2�T�(�m��Ү-���5�;w������$"8i���Ov��YC�Z;��d"�w�pd����C�DS�Z\߿���2e��nIn�����y,�(J����j��j���p�������3���+e	#au���9I���KCx/H�y�^�e�ך�Rv��
`Ԍ~����z�ElMnZ�ȟp�o)#%襋�O| �?O���r_�y�t���
�|��l�J�o=g����p(�v�\�
�l�X���O�^�}\'�L �i�9�[r��r�[�[U:�'����jjHL�=l�6�{���C<���*s�Tm��K'�i�j���E��� ���孶�����n%H�!(�	r��蒛w�!�4R��7�͵��(?�%��ޘ�3	Z�]Ҿ���E}�4�j%��Y)��K��ӗQx��2�[�#R�"���oR�p��8Fٰ}����mѷ�6��8�$�|U��EM�!�-?��R�.j�m���B�ȮL��S.l\���G0�&��8��ߪ������5���\v�?�4h���8r�ՒN�t+Cu;�d���/��!G�2�����ٲ娬�$��[�j�$�>q��˳oR��W(4�G����m�͈�'6ؔP�_s3��%fMt�
vδʥi7$�l��\��쁽��Zp���C���yC���b:;K�!s��*?��n'PU�1;���c�����Z%�ȃ��"E��{D	��������oer���gtwOI�笔ԓVɮ�C�s0ۘ�6ۊ'���&RxE:��y�t��x�9��n+���>S�����{Ģ^����yO������dd��I�l�t� �a��R6�06"�_㾳���R�$�˖E�Rk�Y<�jS��>Lx9'��ңG�,G=<�8���Q��v�^��UJ���|%)s�AG$�� ��>ު��<���$�Ժ����~}�ʏD豖�����t�h��ܚ�)���#2e�ű@RB�������gE�����ܓ��"��
{*���1)�Yr�DΛ oVe�����h�9<�f��<� �Na�%6v(ȸwwV�>�^i�!9FQ�r #��+��h�����f�5yg['�7ʊ�,2獙��$�����tC����[�D٨B.&��X������ҳ���.,�Ay��U�\6�^ך	�v^�[sk�o�/P[N	�]p�z��Pq��Ȑ���Z��B+q<d���� T>���i��<7J�B��R�RXԃ'�ugb�B(���k��R;��آ��m�%��xZ���}��Pt�g{{�{�S�9�Oj�@:�c�0D:��P9]�->��RJ�fxGOm߼8�!΀�^:�5GVH�pN.ŉ<�hz#�tQ�m�hs�ͻ-�7���	�����g���=���k��ꙕL���7�B������/oa��^�.$VO"��L3Vh;��ު9SF}S���dT9ݠ��1T���+�rM�8o~�����©YmrcD�����L_{����#[n���g�W۠ʹ�B�刿�� `Ց��̇zz��r��stOJ��)̹��A�Թh���H������^=5]�mf�d;��M������Ӣ��r�d<��:)yV���[�V�δ���%�9i=������l!����Ρ~�TE:%u�4׳[�A�/ ����G�#��fo�j�VE���J���j�<p�� +��(��K�e�pM ��!��q�ze���wp�e�_�eM�O��s����VL�֜��d-�;�XJ�c3�p���<����h�����Wnn�3��H� �F�d_��rf��>�n�Hց�܇��@��j�,p��M�,|4*�D�?KbN��^�i���Ϭ���J�������zk�5
MN����˓Z��#�	fe���c���Mv�(��6�T]�T�a0_"���+N����Q�Huz�
��gr�]�W�(����=7�>	Gb�2��qT�����A(�Q>��e��(�����ŋeV9WAD���4'?��R�d�]N1�� �XQ �2�i4�|��G�y���@U꒦�i$�6!�ZW_�r&-Bl�wv��pn�)���� $$r��u��&A���
�<L"�Yu��Uo�}�3��Cx�Z���'?�4���8�y����ޞ�xm~�Yfjv�P]nb8R8@T�A>xFxUo�R���o�L~��CY:Bq���e��e�d�A�'�P!���@���2�47p���1n�!�c�ߜPeRW�P*��v+Ӑ�s�u�Z_�A$׼্�gAAp���'����;?���(L�sͤl����\�wJuO����z�aR�	��Ξ�sa�(�1�M��^�:(H��M)"W9#]H��Ӆ0%͋��n6�� Otu\ܘ�R���aB��BH�P�����x�/[��H9�}*6,�H#��x6�w{�~ 2H�_e�E����z�?l�����`���,(��\��3�����*�@�>b�� <�u\.�.�=%�䇖�LR�ɼ^�t�[��ϱ����W�wo���NͰ<�)��&"j�<ǖ"N=i^o���U��7��$�8;֍8{�g��=�/n6e��!�t��[���6-�S���F��t,=�`�I�,C8������]����R��]J���΂��1xb�Jm��u�C�T��>��԰<�3�jhp�~�Ww�	p�V7�yފ������Ζ;�/�y ��M��.�$��d�c�_�@�q�q,xZA�7j�+c�zݡ�Pܧ��f�x��fr*f~�!YG
SJ׍�^��O�I�n��lN�+��:���8B��g@�#��k��C�N�Z�Σ �eЖ(9 #��;6��8ŦI縫cl�
�x�Ы�r�|��ފJ�*�Q��N$'dlw;�������K4��:�!aP,|e_x)�%�2y�{�Eԉ߃���k�~�Ճ�6�3����F�d�n��@��ϣr!��,�E���k��ux��ж�F>���b�J��nN���ϣB��ޛ��y�KH�<w�b#'���L���,-S����@q�:Ľδ-�4��A�X�Jx�۟>�w=&�M��r�a�r�኉��zd\H��@,A{̮ M")?�IH-�b�s�
��������l��w�b�wbz�0��6{1v��~���SQc����lIxdC�܋m��� xP��}�b�>7 ���pw��s��叮z$��nbTA�����樖�QNv�Ml��cG!�a� ��(����F����w�NR	i�z�H Z��-�����[w�;�ުĢ�q�67e�J���O�2����нR�4Zơq���M%ɼ|��(��2$�M�v��q �6R83[Fd![E���W��Џ�mH��BF]���a�@		_����2�\��(�fJ���Wm�>�㸢��O�:"7t�����j7FqT�υWs��`��GC#�y�Oq?���;�+��[6�>��wMq�+�ZD4Jӧ0U�� ��os�kn���j~�c�����U[��ս ��K����LuA�:�(�qc}
��x)elv,���ڜ͹w13�=\vW�r�P<%����7���;�EqH4��f��q��i)5�|V�=C�_�t�%m��M�<�Dc3���Z���I&�V�QĬ����,.����0��mli�g��*��RM���6gD�@z���F���R�Jvg^Q3���k�N�?;�\8X��R3*�Y��]�4$E��޹�����O���r"B�a-�1j�+��"���lkn���*Q��<��'�Wq�y
9�/�x�O�����s��B)�u;d�B	�4���\��Ju�"Rq�146e��2gu�������������*��T�h��jR�F((���������TQ�e�]�#m��ʓ���p.�8�����t�����
�t��3�����Š@D�g>G��G�l�TL���ӻҔSj��_�5Y@.[��̽N��G��,��X�ǻ�YL	��C��s.hrb�O�_����zج6Q0��]��G�I�8�RT�z�� �=h��3��$��c�r�/H��Yy�C~��=��t�J��n���v�`��~$�[�S/�(�i=�}$
֧(O��/�`;;��O��`��F�9�N��Dε��nF��L� KvHV�IL����regR��N&�o�Yp�<��ɵ�ݱ��$�$2˱�-�@t�w0ῠ�c�㏷pr�)νƒ�K9
�}QI;�y�PZ�h�U8��	य़���mPn��ۋ��rש��X:�!�,OzR�+Im���m�i��_چ���z���Z����$7D��e◼�[�Q�CT��X%�O�ߛMgViਭa.؏����k7{�CS��[�	�ْlΞ�ۦ�F��{
�<�t �
�k���Z�v-��v�j�)�I�l![Χ�3���V�C���qYc:����⬇�n�y�"��fl?���U�HT�\�p��-ֿ_�,Bǆ�K����y�tZGt�l�UQ=���!�_�DX�bJg�W21�,�c�\yC�4�D:�O����H,�t��*�e�Hb�y+�Z.-<\n�����x�P�_��!(I�7X��#���ڸE,'���Z�I��dl�Z9v�ào��_"���=$�c�H+��NNxg��:�B�%�B���G��4�r�Hx�m�����z|��	-�V�}>����}��yo�66;���AXw�K�4��f.�Wacc�oE�Z,��B�K{�=����dƆv/���6N���tae����H U*��`� ��A9��poz�{���
X{a�i�e�@w����b{������<�-Т�M�<���Z�)5f�/����^X�@p!�����o���F��$��/�J�	o�f��	��˸,�j�t������9�H)J�������E&�m�o� �)�Fx*�i��x>6`>���}�\�'�WK��ܞ�nE%+ؑ?¿�E� >_�}���z�M�~/�9x+2Z�g]�<�����ӫBF�K���!�6��lS!M"P��>��1tٖ�!!���"��8����z�	�)I���K��.�xċ�3~�/qy� Y�ڤ�1&;�x�io�`	"��%��8����ݙ��!zkh��p�!8�pk�9}�q���bH}�:�i��Vʩ� H��Y
�2C"]�
֫)&w��C�,`P���h|�2�F�_nz:�� ��'p)�@%�:C���'�����v�"�e��CK��_Nn�����;���v�q��{�p:<��
h���) �`�,zLMܼ�����'\ebFuM\��A-y:W�?����P$��U�tJ�p��.�N�<��N�	u*a^�vxƯ�T���2:f��I
R	}���ɏ��0�*I�x���6Ҋ;V%�2h~�O2N�}�d4��|��j�2��Zp��� $Hpp�kg�K5��%��aԻ�Shw1�x

Ď�|r�(��BIm�F�lM���a�.$�`i��*Kl>�z��r���[�C0�c �+�7:����ywL&�*k�ס��7�a�zdW6�s&{"wby�����_R�G�ǅ��~|�|j9���Od6�:�n�����f\}�����b`���Xﱀܜ�d�����)�s�hi���S��_�"�l��W�VS�۱l(>�M8��w�"��8��+��Km�1��@
�i����ŀ�zs�ҕV��R͍=L�݄c5�H��������f����dѰ�f�o� <��x�T��T	�7U���sA1H�����?θ�I�ĵ�!��xHgcڦ��M��@��k���E����g{䉏}��P����^�%4*8S��?H�t�RĽ;֯m�cR�Z����#���!CN lݺ���1�{�t�ǘ�j��_{*��kA�ޭ�� >�Ox~+�h����
/Ӂt����zƍy�C�s��M����sҲC5Fٷ�L�'���o�l5*�۲U����Q;m�*�+߭�������������k+�g@&��f��O���;�A��x�r<*�M�l�ۦ�E�A��W�Y�� l��(N/͠w�Sݟ�g��5ꬶbL9��v��1�K�L�eb��X4��e�r_-2�~9,�f����p1&*�Դ��T'.%=R����W�=��	N"�E�B���&���B�B|��:�Й��<�
�#��j�����&_~]]r����(7f�����Y Z�Ck��l�_�|�H4�_�i;>E<�V�H�2�Ֆgl^u�ʴ�I�B�J�+K|��XK��!�R�ɺ�cLPH�p�u��f��'�-Śo2%A�]V����O��T+�&}��swF�&����e0����ʠ�K��bCX�q��N�÷}3��59Iդ��u�<��bϖ4�sP���'M�j��Ύ/X�=n$�Q�|�1s�?)*(�ϴ��O���xb�^UJ�HF�kG���w��<�;E�tʤ� r�'<;!9�`��j���9��v�,�౩��7��}`�K~�/W���*X�p ?�e��������|��`M8O��}0�6�aZ�xw�܀$D�3� 6\�2P�J��RtC�����U C���ۄ�Js9�1^��(
>[8���$J!�P��:yAn��c��z�~Hm
����j }�x�f[2&��mp���/4�d7B���8�JR-�}�v��	���v�){�fGU�o���6`d�5n�0�&y\�;=7��)�W7[V��傦g���Q�W[k5-��ΐ
�(���2�'�ϐ�W� �nE_�\�S,=�(=���*����;��N�K���L���굿ڸ"�I����,ɯ*�S�}lv���T��a
�u�ph��c���p�
J�^��ۥ�u����ĳ[�]��|�cn�G�}���'��i��R���=��N��F�ߠ���7�y�$���<��R���t�+�r�-��"�<.�Mɦ��GJ�˕G�*
4F E�~��%'�{NZ���� �rz[79�5	��{7�|;BP�S5���4C�qn`�wO�$���E��fN�o_z�g�8�ʮ&��(�c�h�$^6!)���L���Ţ|$v��粟�����Ն�B���.��k�*k��QE����EO�����3���p�S�U��!�r|��U�9�v3 2�y't����G���Cl5>���o=~�����N��
����s7ɺY��܎|ʼ�?��T��D,cP�? ��3����=ĎB^�!�\���9Љx�ep�k�ZgGq6ѵ�$�ZU��ys{=C����`u���vL9�G���ֲj�0����P���=��f�U��<p�4}�r~�e#+&u?�e��K�����˻�6��<((^װ��B�8I����5�?��_���V|�V�q(s��S�g�mGg���1�GUS�f+��P�:V���Y���'�ڜLo��P��]�Jɝ���=+"#%�.㯝�.$|�.��d�I'�+������8�c��h����L�HIX&����s��Z�c���B['��w�b�[��j�;�潼&�a8��Y�5��2shũdq3�����yc�#��;�t�7;Xo�E��"̸n+��mIb��)��V#�?�H�ug����R>�i>�d��7~f �	;¡ޠX�ԁ4x�g��>3�J
�8.�9'@
�Xan$E�1kWÖc�Ӣ��SͿfmm���F
W#�D�X&���o���
>�+"(�xe�ʥX�����b�v���H	�>!��h:��}��փ~{����j�Å����z�S-.��-2��/৶���(�XB�s����o4o�dv�6Zg%���t߳��,\�?5׭�Aſ�`��B��-]!=dC,Fƀj��x�4@{2��q�_4l�M���b�v'��Si"�t����CZ��06 �w��S�	���fm�XF`UUj�tf�M�����x�!�ɷS�i�CVא8a
M�e���Z�/����>�Lp"Q�C��C�^���j�NR���{���D&�(�=�1�S\4N�
�1�{���z�$����'��YD���2�&a��C��L$G��I�n߼�|��v#kȚ~��A����&DJ7��_�G�t����"�-_��D\���� 9w�!E�~:���� �PY��!K��+���9:�MPJw� �/]Y/N�)6k��k����%�P���5�a��K���]���
Yj�a�o^6�0���	�yN8�����z�����Þ��=>`��2�yPs��c[d�O
 Y @��v�x�%w5@-	���ٸ�_��.�o�և���Oo�blD�&	g)iB���AIH��Z9�;��Ȏ-V놡0�`8/I9S�L��G3���Cݘ�o_V�a$�	Yк1�x�aM_���mX�|�}��H�c
(�"˱Ɨ�e�}��S?��)f;.p�q�NK�� �H��I�vz�C���lP�������_��HÂ�"� #��Bx�P�7S�����'a��Nb�G������]tg�d
���$U�Z5�ǝe&	�����X�)�O�G�PB���V�q��F�C�TJ5R.�ʐ�*e�;�n�ؿ�Q9�c��?Wd�r�Č�_'�V�4P/�$��k��,�Yj<Nƺ�T����-F�����sd	^���͢X�A$~�AKz��\�2���|͛Y/8��xS:"����a���$��҂�>}�N:^Y[z���2�K"`>�>e�+��;=H|EJԫ�d��R��#��*�p��2�;�4#���m�&�Ϳ�+����<!�������)HT�[��S}�^�<U1��b�?(�U?�F>�`��*�r_��miq͠��}gpN���D��9��;n�j�IGwF��)�~�d�?���`�ڰ��Zn*"�*�?�&*t�j����9��
Z'쮝��2���<G�!T�)����(D���'Ҹx��n���\���)8��Og����ϴ�*ܳ�)���āe5�@���卯1e>Q�R��J����, �7e�\�Z�u�e2e�_{��Sv*���@Wtv����( ��ܿ�/�p"���������b�/=H��Jkg%�C��o�/{9-��,yLG,|�fi�O��d�5GoIA�����U���TZ� �d��&H���ʋ-�~��`�����nz����6�\=ą�^�Y���B_���N�r���<�p^���J�1��ί�噅����i}ka-��!$����	@�:�,�A�g�N�)[���w*	��0�3���j���;�HC/�l��YA&�T�L,��E��Ǩ�|)+�4�W�E���m��,�{�������:&�moK�1y�~��L�4�WV&���fn��z������	W��v�n����׭�aVp3Mܖ~<D�;d�-��И�_
"�u�+���΋��ue̜Z,��] ���7��a6K��Q�b����6A�IIt졫Е���̧�7���>��JUv��1���ǜe����4Fp�V�'LV�y�- $=]9�!��I��Sa���k39�nzh���^�6��@a{�����^��Q��^���>���6��f)��}��VFn���qδ�h7eD���BV;��/5�0����jb!Zx$O��>�>T�k�������N�o��X�	�
O̯D��t|�����̚C���=+�o^�6�ֈV��|?W�M4��:%bm���eZ"W��A�&\�-�d=1��W��P妙��
�E�|~�V�N�q�+͢GHL��>�1�V$�_OX��fw�����O��7�X6Gd��0l|҇O��b�3�a �ù�S\�D�>V~@X!s#�@��Mt.���l��eeLg�w,)��Y �͜�1�?��bc9Q^��� B"��ex3��fh���z��O���Ӳ�Qi�/<ˡ���Pg��;����G��þ�%��
�:W�5�}Zk���#�#ػ�z�H��߈�S��[:�2+�� z����*�UYG3+�3@ �k>7��vX���?�D��F�̝W���V� ��XX,�C�0�G����q���]~$�a�r�O��`�#��%���R&l�Ӗ�W2����c�e�ͩ�j|�C��'��O�ӳ�@�vf���jԱ�+��_)/���KI��'�;�1���-���CG!!����F@W+W2��L
A�`\T�;9�a+�C2���(�o��A򫎥*YF^�?�ep	 ��L��
�]ȇ߭�-��m�wL��NК!�� |�J�'����rݦM�a��[�&�s.�;�W��N��5�'��k��h&��?����0��|��$cM61�P�`�*E�3a�|y�����-䑡`�v,�Xm�`a����b�<X�U*߼�w��k�O�YK�xړ?�_n�������c�v��xd��H5���+^�ٛ�2�����cǎ�J⪬�nk�5Tk�r+���oB�\ʽM���sZ&OS1��LatȦg���l���'�E�+�d�ͥ(g2����rQ��k�6����Ғ=2t>K�P��߯��q���TK�
D�)B�O"b�e�����[�9`������L��0�U���g;q��idz�%�o[�O�����U���Z��t��C��݊�*�NN�n6����ϔ*�.`�m}�H�h	>�C��"Q!��/�=���֜0TW˶�2M`?�w��2��<��8g��A���n������M��9�����KwC�"���K痉N�{�B�]���9Y\MM�:���4S�a���Y\�&�hA}�Ӳ��`gMP��<˝���>$6K�S�y��<j?Y���9'��wВ�ŕ�$����+Paҡ4����:�g�F�ܒ���	E0��`i���E�քDe�Ud�O:���;�r�� �������~�u-�/H�	���>n��v{�<<������'��3C[��m��A �O踣@�I�[~�;��)0QH�7{��R����6i��0\�o1�oc��tF���Wi�2ni^u\	d0V5�(C(�쓄/	Y�H]~?��cǻ���)�Q	M��/>���^c���xA���/��<b_ܷ��xbGi����e���n�di����>�:���C8�/�1,s���r�xBޣG�G���2���jܾ�
�E�����H��<���n<i#��=��ܡ�����Z߰m�?�q����I���}�5�2-�)Z����Yҧ�`��6f˙Ͳ5'�c����VWW�]���󛺔���5������I���f?=YjHx�bWbb逸���Z�`�wc�|��d��������lܪ%�����<T{��SjiV�iB�����`!����(@��ƻ�Y�sRH����ӹk0��A�~��=SW�䤙Ѻl���z���/�r_>�1�<��h����m�HX���R��U�6T��v�O�z4�!���>uq����FD�lΕ�q��[ؘ��Җ�h�hi�0�_���^Aa��5Ӊ���5��61��|�Q �DV&�A	_���h���sT�'擄[�Z��\�I?"l������LB����@��䨙���U��2�e)�Uo�oa�
�W#��>��[�*:^����ᩕ�<�ܨ�kJ��Rȉ}
�9V6E6d�bO�����T�>�O�w]0�k餢6��Qp�J��'DV�Y��:�"�ʾ��nF]$�KZ�l����Hn��n\1tK�D��/l�rE"�(�� Z`� �9�g����H�?#�a�O�������Ľ5�=�H��r�,���>.	l�#k�+-��d��5e�?X�lm,��\��9��J��z�2?ɞ�H��K��JS�� 脜�J��i���UȜ_���xh|yk���*D5W/vڂ����y_�X������So3�Ri���xY��5����ʙ��yR� p��R%6�?>3n8�H���.�`��?4: Ϟ�e�Gt�����D�I ��է;O��!N��|�Xp���N��#]���4��l��Cʆ�<ՅQ�vy�p����N�����4��O���O�3ԓ�W�X��b�"�?A�	1;�
`�I�°��%7��l�P���p�q�I��G1� 6�����Y/�&�OP�ϗ-��Jwa}��(\E�xs6�X���ԨZ!o��x�sB�S���^�HN	%<��|���i�ޅ����p��(��u�%5�զ�J�|ug�E[/�poX��`c^P��@c����ŀ�����޶,q�P�z�2��L�>��o�J�[��2:�����0I-��Q�li)��H~9�)6@z���B�{��'��8e���\1:�69�����|��|����.��&>ZYz��A�f�: �2��l���BA�IG�l��.�y.tk,��s�����7 ��Tw�uG��+���*�����:��(8͍yT�:��[�v��oA��]w7J{Uў5J[�90�����Y�ޱ�{��*�}3t������E��L>`��de^��>�&߀	}(v?Wc���H���,B�/m]`���kd�oZL*{�_k�P�}���Lw�f���ipi ��.�'/>T�<(S!�2�伌ZX3��Ќ�\Y�� ��e/Ն.x���&�/�a>)g��#�U�����p�|8m�9�r|��Rt��ٳ�YM�ܑaz(��BxS��*�2�x� �W�6���@^�����S	���r/���q��yq]�ޯɺ�"���ȷe@#8�갹,d�#گ7��$����нJ?.�����]�q>*���EF�[�\7S��A7����Z�V�韬�8W�*p ��sbS��Sa��\j�������#�Q2��?��?��}݈}����|q@L���q���C�(zw{!�!�>��U���vE�+E�zԞ�>�ok�^E�0d�>R�HLV|P���e<�=e�7F�7>0]��%�$�I�:��-77�o���nB;���8�3��+n|'�=})NM�����7[�r���uC�dJ�IgeH�$����w�@����C�?/&�wlb��x����2F���N��]��9(��ޜ�+�0�~��Ӱ,?n> �vO3wj��M
0K� 2�/rm�
~��Ӄ�6���6H���8rM��e�fB�qQ�����:&��,0.�d�ЧLaf�ޜR{�7����Z�i�7j!�6J�ͣ]�-D�D�@0���n3��� ��.Dr�r0�C�>V���1������\�}�{���Q��T�.�ü��{G��sϚ����NvU�	� 7q�"O=s!Z�r��2���h����Ʒ�"��KUI�NZ��2��K�gg�����(�{�8����
i�Đ\q�]~5��E�f��i����QZ��m'�>
���wI�����`K�8���*���yP���4B5Bm(G$^�eGqLb�!D��앐�|��b�\��
L#����$��@�|t�8k�f�s�F�x��<5D#�6��"���y���]��=;��`�KJ�U
�/-l���劧NF1[�"�����v�M��a�╾�=��M���g���$<�_~ `��i�f�%���z���g1fI�p�u?��|����-ݭR��[}���|��^�?�L?�����dY�U$L��1>����qe�f��`����s|��"�N���/�b�����S�� ������
�� j�~��RF��"�R=F�ڥ�a3�G� ܶ��*���u=gq�E�ʹ�G2�uU�M@D=&�&�>��^��%{�Z��jb�L�ZI?�Ⱟ<�x�B>���<>Wgn��p�K�ԳȮy��&����<b>O���������W�#������pjfh�
���0\�l����k������b�B�&�Ti�{�ϵ.äCRk6�6��['/֩w^K=����g�n�����
r�ԫ:��!͟����AZ���>�z���U΀����)୓w�(?��E��z�Y5�؃�v��H8�'$=[��[�s��_z��.��ˢ�fLfF�=���kwi�*ǈ3"�r��R ����0����ԥ�e[xtCLr|$ȈL���%:>?����B���-��WT��ا7U���u�?fϡ�<Wm��6�5�i�)֠�~���0���Cݛ���XN�bM���!�ʶ���֎A~�#�uC������4�S���ډ	4v5�$]�a顄|\��g�t�;�r����ތl���/eu�K�G��*&g����q&V�����:Ό�i:��>�X�\��OL�=��Vٮ�E������*؊���������G`���S���}�. uf2m�E��Fj!w�?��PHP?���t�����[M�>ָ��GܫM
�O4�m����9g�i����� ����L����c�Ӓm�n�-�w�$�dc�7k������4X]��I�cS�����x��BD�r����x�rx���KfР����"n��'��9�1��;?f,��C?�Ծ���8�Z�B*q�����Q`�����vH(�����~F�6Ku����9�a�X�O�f�^�S��"ҽ߁��O��"e4@������1�"��[�<F	t�E����ƽ�g�	���yR�"Y�W!��;ɒd��o�;�w����#��
��K��P�i���-�9�U��͜��Sv>����Se��"7i��@�(="%"�d64��/>鸆������x�N\y���;B�D$�	G��J�A!��'Φ�`�ń�03�1��S����F@�O��n2����j}]����R�6�p5�EJ���u�l&�؛\F���ee)�i�#i0M�o��/��g|Z�it��{��^pl�$�L$��k�{ʿe#K��([� �*���roA=q$O�Y&.+̞��FZ�_=�=Hd\��_��o��P$]�3�F�GyYr+m
�����V�hE���[�]6C�W)��~Py�2lŁ4���m.�G�S�>2�b�o{y�I�z.����$鍂u���nף���<v��	��#C�Ej�Bl���n%S0�%l��g���������6�����ۚ�v]8�rH��$�b�x	�+i��r���F�6�Q�JES4~�X��ccn��B�d���1I�����E�P�j��::�m�w�b��z
���f.Pi��;
+l�����\REi��ŝ�ڎ�ʧ���p}��v�9t��H�e21���[�P���d��MiX�e+4��2���jQ��z&SkM��Uiz�Ys��X_U�%]�]�,�Q$����}�p�� ���x�V@>�$I�3���1�=wc��O�����5����c����X,�鐦�1�[��~ ���.h�n]�<��*{}7PG�d�J���!x��3��Ús�#j�"f��.�����$l��_�]D茤��O�:��Bv�Ayy4�,q$�
�z*����l9�R� �Y2ƍ�B�-#{��Gg�&�(��i0/�<�A�
w�1S��I�Wխrb�y��'�j�BT�:�n�)����s��c����CPwyŋEG��V��7S�SŘ5�QC�TN����pl~�8[#���y��3��Wm��1ڮ���߃&|�2����Y�$�g6�s�2���b�9�o=�M\�)�� 6+TTe���>�|C?��A��#��HL�y���ZDf�д��ޘ��T�E�n,�����o26��e?򘂶aD�1{��ī�7�f	q�)J���D�"y_��i���S���\�<���YV�V���6�N�Q]��$��p�=v���E|j%x'��Ӽ�5��"�NH�QG�@o��,QŅ�8�K�i>Ր�(���Aオ恥���C��x#45d4���W		��E�w�[���%*�Z;�@�G	˧����_�0���<��[{�&���v�%�p�w����0}���16-����b��ݻ�gW�qIGf�Hds,�K�ldL�j�,Z�����W�4��\� �4���h�'�.�?�W�'Mm���9��ޣ�����jy���S��캗YQ�O�/;P׾��u�
��ơ��
GK�'M���{����9r7y҇~T@���iĔ~	V��J�~a6��E&T� d���]���@�,0MƣWؾ(���p/�O�H��!��S�7[q�w��q�B�.�U����f�g��"��\HWo{��K����1��1�|)�.<��������d&s�"��÷�3荭��Z$��D��§��9z���V���o7Hsɐ"(k�jjd.7������AJ#�?vk"Wr@�%�9}���9�&pK�H��IGx�A���7�&Զ�r�z��L�ɆǟnO6k6���^W�c_�\���bk������O��:��,]�~@�j�i ��6�������+ �H�CO�G�
��Ju�3	r�I;�#��C޶���`:i\�8�%����ݻ5��d��R� BY�U�/X�� w���r!��^#�����I4�w��-bvi�Ì������|8��ƾ�o�lp[{|�Ĳi�*n���~h���ULv�}�!T�.���'�ȕ>�_}��J�K�Wom���Hm�p�0)Gg�]X�4���8���RV��E�Z>*�����q�>1r׵˿��M��}V��sF`n�@��#,��P��D�y��=�Йm�7�U�T�Q��d?`j�rn.���''1*���A��.���1��f�잴��\:���4,����=p��5nxbM$fg�$"g�]m�S�|O��h5��l;��zW���:�у�i�DC�=G]ЩU�� ��؇*���u��傿��c��B�~�q�������s0�|`Iz�c$�y�k�����­+ȓL1̊|�T�ar��-j+�}U��c��a�������6;k�EBOs�}Q����(2�˄t��)��+$v�V���E�\Q_��2���F!V��ǐ�Y�f��2�a��������4�W�p8�Y���6C	gU�����݉%�H~	���覑F�Cr�{���I=��(���Ą���MTS����	�W\����퓋z�y�;����|��f+u�cv@�{�Q����+�;@q��׸�gWb��{��)�,5>�ZA�&��bD6���uRg��}D�]6�@�XS��?�v�t឴��8X9�����<k��i�阻�f g�4Ck��Wk���}F��¨����<�V����g^s�F�'�.��f��1@��I)���և>8�<#��T�J���r.$��U�1��ʇ����NO@�Y9gߎ�y�^͜�
�П6���aX��l�Y�O����K	�>�� N�Xq<o������3f�}E�}���XΎ���9�K��'I@��G���}�3��*�iNlp`H@.p�mf�����3~{&���= %������a��DE�C��n߄�U �W�#�������Aj��@� x ���E�頲e��Ѿ�p��r��=�����v�g[@�^8��^��Lb	7�T��R�ƖK����~d��H��u^�ݱ���77Z0�Eq�Nz��{��h>�tE0b�]�gc�֫`�"���3ʼ��k���Fag�=6u�-,�p �⠷p�HԬ�Mq�8DK�]�Z�?{W�˭���q����7~ݠ>%�������qF>�3e�9ԍ�ݚ�j+��)g�u	�$�aRDP�1�#�� `/���_��@�	⍝m�{�i�;���U��C��1�$�?8�6/���E�~�q�@J6�$R^�k�O|p.
����`�כ,q��	��<�����a�yR,���U�ΠӮ�?F�0�?�W_�,&�~�M�$�:�����R����4Tfظ�j��=ײT{U�?��C�SZ���[.FW*��<�o��^���AM�bD(b�jU�+�!?�+X�����?���x�l�N6KW����6<�"jB��*ᱨ �0���9a��-"a�2�ٞ�w�K��$���g^�����]���s��5zo/���
��c@|݃I�E�:�/��҃�9�=G�H�����!�;z�W����i;Nϥм$#Yk�%��]���\'k�C��\�@�m�u��������Q�q�G=r�oq<,�vkT�A���&��f`tp,|��㐉h�m�����1kԌ��y�y&mQ��P�y7D���רI<�K|�߂�N��������l3��މ�����_�nN�������´�z�*j&G�2${$��H�'�psK9X3���_�vM�X����vue���΍��u�Rވd�~�a�ڠJ�/]&���]��|[��{��G�`ng��X�WW��,�HQ�i���x/���� 2\�9�O	yr��hb��X���ؗCy-ىs`�;�K	��]�B��l���,�>�Xލ�����.ï���;وyܧ���xrH���)�QGb��]6�&��k������7��	�V�ӝU�38���%,��� ��7�����	i��ku��mT���ի7�8W��tFDU�:��g 3k�q�����[��g�k����-��j����*�qK�5Mj[\�RyƊ��z�R"/�����������/y�Z��|�p�x.�9���{���P�ÜM�e�@� �B�����m0�d�5Y�x�M�"Tgp�?�T]��r'��+���pܦ�G^�X���'��*�:��
��j���d�o6��E�Vu��&=�)�A'�>E��ҥ���!���LWB��a7/H�� �!�C�y��n���t}Uo��� l�{ߔ%M�}��)�K���O�/�]IP�}���zo�S3t��<�p�gA6��'f�[=�h���|bT����"�rr�m^-��;��}�#<'��taثO�$T5K⹫N~���9�.e_�x��8wT�yC�Xp�H��
6KИ�uf�����c��y��>Qo���^?�d"��
Cu�m'��7�^���f'7��m���	�+��
Ⱥ͚��Ky�oU��+���c'�T=_ n�I�dP�2�e~�Sf��V���[C��E��j�q+6�߱��Qt���N˽�9�w/�t��X��@)_�F�ź;�y~M7�6�"l 2/2,�b&R��&]f�A��I<�ZaG��v����7��0]�\��)y_�:�d��|r�Ϋ��A��qQii�C�G������L�w&
hJ�]WUB��I�B�����[ܖS �島4� �"1�'3e���bv�YQ�#��Ļ��A`2*ȱpЎY�5��Ep�ᡗ��XΎ�G œj"�����
���4|P�&�6
������F9��0�H��L6EԼ����g�?���8,
iP���${R��~�֒�'�C��v2�)���JzMy��6�>.X;�^LU�e?5�j���dX��b��ɪ����S�{7�T{�)zPYZ$�/�DC�U�;1�\l�7u-�O�`��"$╄�8���\�h/�l�o��*�0W=w�.0�O�u
u���~^h�y7�A��`W�z���o_&q��.J/�PE�*��QpjVxs����S7�8�K�=�0���$�V�aϻ	XL��AkO��׉vH"Y�"�]N%t��P
�㉄���޵.n�����<��R��>��Pn�4���^}��]B(�_�<�۲��J~���.�H�����eN��>r��:�ɢ�f�}�6�M��B0�NF�*�+k63Ѱ7�
V�6Y�_�-8��|�_�w��5ouz7���ĉ+���։�:X�}!�4+t�@�V	W-���Y�����<q��9��9�w��Dv��- �>-eڴ(�C���✇\�c�.ƅXW����jʭ��+F1x�́p\?��R�}A���-O��ͪ��'��}��=ʿ+�d�kUx`S��%l�9��D�&��	�3�kD�۪]����x��-}E��׷�h6��-\"�j��mNN�a�ǔ�t|~|�m��`"xUfz��<W�e���H�\Ϗ`/��DX����,-?�(�,�iA�Io"�Sl"{A�Z�8c�Γ�����gǡ�gg��f���~�&}�?����a��{~٥`��������h���L�
�������ŗ������b�!����!����G����T g3��w��X4sR�Qb��Ltb�I��i~�bL��t���|��i�rS�E(qg�iʲN�.�mZ��X�j�[�����#fP�KWg��:=~�tf"ՓX?"�Q�jG�ްK&��H>a��6�o/�f�ς^�f��ҋ� �^?s����Ԁ��?Th�Fq\�n�\�O�j'?xXt��KV_	�P��Z��p*��*��f*(S�<��[��k"�y/�+�^���������?4�cs��;#�缯���&�m��᱊NBɧ.
�,.�ͪakB���Y��Lr�G��Z��E���8��f��i::�祆-��y�D���k��LW	~fz�\G|R ���S)l�^�1�:]� � %�#� ��-����V7ܑ�T���< D���x�H�xK|	ML��u��������܄�(_�$կ'�(�:��b���.�o�a�o�y&o���oX���W¿������(%��ݤai���Ϯ���|�,��ʗ>m9�p#�4���0XK������r%��~h|��(��#��T�Te�h���vk���g6�b�Jfƾ��v�q��:�����W�N+M�h�f�[t�J*4����u�ψ��(��pY%A��s(;�Ó�s��%_�*W6Z,=�rxXF�!t�:ʶ�{U#��ڞ�W��~^M��Sw�R�w�r8�g3)����k�!�[�~8m���1H[*����IH����/�Ze��G$���w�g��ߘi�5v�(g`�HG��k��ף���~�r^����Q�i�⒠�> �>��n���=�`����vݼ�8S�y���>4�kA\��i2P��g�?�B��f!zbӴ�=�8%e�Y	���"�i�q�q�&��]?����l�z]tf�
�運5�f�:�c~��$�#WQ�����"t� ��X�Td��^C.�^�h�М*�a�,wu���8��3��]g�pD�&$i�����Ę(��2����")�����{Db��HE0��1�PI�y؅-X�q���A�3o��ӄ���Ytw
�s�%K��E����:%���l���%��apPe{�y 57&zӐ�0�*(��s��U�p���ڄ���_'e'1e5,�U~AH6"�L�+�P��cS��QQ��E�"��2(F��sM�X�؄l߬)�øE�<T#���Vv�|�vV+/>d>5�q��#�?|�a��vUg�-����o=���-�2#��
ď�:~�!�z�� _���)?C�Z���i3�E�!�b+���	_羺R���q��L!��)
�M�!2U&P�R*��1�CV��;��h<R^�s3��$ �� <S�K��l�X�ɜ����aWj5���a�~�֘�Q�*��v������+�TƂ+��� o�wʟσڰ�}�1��/���p�����1dfe�/�A�]�/_���:�]���<x]7�@�}�"s����˯����"��w�����ɡz-O���O���8�>m���C`1����88�$�S@���{Lb�.�][g��:2�����9�L\��x;J��Ԍ�?[��i"d&Z�|*��_�7����Ã �:-���(z�:�e��מO̘^݌ �v�_E���m�Lz�M�6CT�_�s7�, ����f�t�T�s��|1_Y6'\������gS�j���L��$i`Ͽ�M1n#t4���i`s���US��A���v5^��FB��~OE1�Gf;rxC�(����cG�w��!A �	*���!hw�ՠ�G�Fh���^��߻}Nz@~�
��d���@���V]�>�����/k�y�Y�f�)� B�R'D�O�IA�����z�W85�a�z���I��zE�e�B 0���c�&��Y�i�! #�+D+�08L! ��V��`��30�1T^O��]�(z�A�)��f�^�UԵ�Զ���E,0X���N�6�J���^�&d����x�`L�%fh,��/�;)�H-}|Zj�_�˞�����w���5.�_{�D���~���<VS$���5��(�UY4��s�p�+u��<�9�F�9m~c��L��`��/l1Z��O�)HX@jr����<3���g���E\ǉ�|�yZ�<�zd��v����j��*A�;���_c��=dJ��2.ߊ�Ψu��JO�
�{��I��UT��ڸ�K�ߤ�v���l�2��u��6���U�I���������dǓ{��c{ի�'T�fbd�c��V]w��$`��6Diɹ���ԙ�y����@��]cB��׃������WA �xi���	�xE�C͢���*ˬe>��4��/�~<;R�/��T��5�̒ͮE��%�_�@��%0#g�>�`,�!r3�+�*lǗ�b��W|�C��*����?T���ra�z�E
s��cL׽�`)B��A�O�r6��:�Ƀ��H�!�cf��3�k����z����T�:."�y�G[R1�IlVE>'q���+}��-*���B,o�N�HY4�7v�"F���ǲ�,K���כɔ*�9����Pa��mti�i����ᗯ�g����f�ir�[�.П;�!	�iL����������-��J��$R�P�t4��H0�v&yY��u��5��(�6�h��t��z(�@�W��F�f��g��P'B��9�~���j������H� 7����/��c��M��Y�˙�<�����D�(I�f�����M1~���>L�g&�B����l�4���!�FI���R�qX�f��B������uN7 �Y�AH�	��1.�A�0�3��JVe��>�~���ױ�� �_�3�ǔ��4o�\1/�RmEЪ���ҙlS��voaٯ�0�A��7C<f�]wJ�@�I��Xp�0���f�0�/�96�Kn�� �sE���:h��cϬV�s��Zk�鳖&��؃�A���	m��9��ٳxS��$_ܦ�ϗ�׮�M(�]��&��Y�J���x~�^��:�/�k�t ��m����rc���>�y��E1��_����.$@b�B��_����5
_��ڦ�)~�4��#�9��*_����I�;R�G��C�p�h>-VZ�EC�wgED
9�̑���YNa���K�yCmp�EVW6Q�pE�&�c�P�t�jw�4m(�W\�"*��W?��@|x2��C�~&S6���>ᥧhLZbpZ�#J��Q	��,�V��E�Z�@8g¢�|{�܄2U�pmr����ǻEo��~|Jq
�Oh%T��>��y��;A����W�>����Hj�:�0L���\=�8��o����n��W8���|�z7T�B�S��������גZ�=�0��kf�*"���J��ӱ�"k�J���VV"�pG���식A��7;Ne�I�B^6�_k�]�;\鱀4ol� �<|�?Ij��S��i�D�o�6��^�]S/�/%�]��P�iO�e�N^�4�(��>�st%����'S�d���x�f�I�huk˔�
n���e6�/}R]���}�;8e�5uzUʽ�����s~����~�p���$���8������iؐ�C�ҥ���V1�x4�-�a]�V�j=F��1뛑��i%��;u o��5d���=�='���$���RیX��k�<fJ�	+�o.w@��6�ۓ��
L�$Մ�o�!��.J�b\�����;&�	�]��}[O�H�&=L�/�ť��Փ/Q��E>W�kn�2�NI�Z�R�2��m�����8M*���;m���^G��w��� p�H����"�i�>܃��¹�dæg�6j���&������y�!�NO�`�B»�O{��A�R�n���~f=�c1�|�q���`7v��F`�s(�6R{��\7����#tFX�㴉"�T*n㽞���,2�V���5����0L_�2:ul��.m�L�ņ�H������naQ�l�s��4I� � �]å���"��,���k^6ѐ��x@W>���'M�!;聬��s�	��d�/n�+�� w�?���'��ɻ�Ê9�,To
�"8P�#XDSa_"T	�DK�$��M�� |����lOM'�fz��������G�ј��Q|n"_��И͕�����4��I�K�a�R�p�.���L�î��Sg�7FL3ꜵ�����i��l�[�p��[ 8�^2_dy���F-e����Y�X�z�,x���?AnR�-�U�P�B۸ә��	fbk�Mz:��dP�:�G��K�]���A77A�C�/��a�9���u���|3�tS�Ԛ�!^��U�b�#���:�_wb���g�Q�E�r�+E�1���=�~��8հňj��\��S �x#�_��
���9�*��φ�Y��Wң�Ж1���ZS�����T�A�)F�v�L�T$�<�i��E�8�[y+����R#�i���Wُ�R��:�N?�����jq�Y��R�����|��^aɉHq��F�d�c`�s�$�~�̊*؅��hMܪd۴&�ƽ���cwXD�D��Er-�F��*);�mvw�U����ʭLhM�T�"��������u @��p^u��t�͇���p��s0�q�:�z�ŭ��Ch� -B����o��U��_�'���.V@q�R�d%t�{��(ޒr�Z����V�tQy��4��_���)"�Mn5�f�fLqt�V�"�������FNˁ�I^F�L'�f���j�+���hp��ʬ�8d��i���:w�b��#�ᓌ�~ݟ뿣a~��9�E�0�  bD�R�R���v�P,�0����F��Z�j��;f�~���I�>���U������`���k�� /�hx%���F#S�R(P�n�T��U��A����pO�&]b���*�Gab\��Aݴ\U(���A�&]_ѽ���@QzR_��u���Go�e<βU��Z��n*�|���!-���� ;й��l��e�#������W:�	]��yE�l��?�y�9��%T�RP;q��-W�)��a��ǵYc[Kր�%K��lpphR�S� `�v^,��[�����E�ڱ^T/7���1���~A��!��)�?��R�r�����8���K��5ͼK:�v��ٯ�e�)GA�OcF6YR���%9.��ӕ�)�F���1�۵M�Sљ@�o��k~���+~e���m��-�7�!��ZDTn��nӎ"*�_gt�hs73�]�ߔ���nNg	�XU��H�q�����5{�y��Ż,�9�io�2�e�լn� ��G5,�	2�iV=�1�)�U=[�"�[�^��O�|߫K���9���W�<�Y	�t�Uӧ�xm�%�c��������[ʼ" �/�NJ���T�w��Hb�$�e�O��F�B*󊝛�׻���M@^@H lvpqH����m��j���Zrp/K�|"��!ym^෠ _0J�d�[�׾�<K���J �mD�愃>±�T-��,}���;;)J�o��cӨ̴]��7W"��`���j:� �5������ے��������@��\m�5Kd������b[��Y�Tw8WN\}��' u���t�0�}���q�P+���z��.��qF��Z��?x�l�C�qF}�:� �d�!���	�b(�@q��~��BZ^���L�4I~k�)*�8�:}�"L8tv�A~j���P*�䢞Il�%,��ÄR�n�
N'C=�*����MQ~���P3p�� t��L�AY�C�/Y�*ܸ��v)D���+Y�¿���L�M��~g(���3����:[�i�C��^ � �XA}y�P�豹���B9_Gt��/����F�E�q1�����[�B)�����W��?LP?��˛�n	T�C4�1��I��&qsz���%ݖ�����`�
hG�V��PtLL��y8�uZ�v����g��7-�����:�=<�'F��no�A�'�@_
�~O���f�n	��OX�ĉ%0�X, hr��?���(�(@�Ӯ�t������]�\���{����kr���kR�j�e���g��67�[�ξ��RR���r�0>���W�X*Y�f�����R�bk(���6���-�s�^�D�/{#-�����:뢐�N��s��h.KY�cH��D߫]�0U^����'?^6�ɞ�@PF��C��X��d���~�b�6��\�,�I����|������U��d)uՒE&|�$���:��0�>���8}cWy�m��-w��i>o R�x��w2���KS����!�� �c՝%{�0c�Ԁ�j�#�<�=�٩,�T�!��zR}%���!|��O�A�
�a���VT�K�^�S�OԲ���k���" "!���`癧n㫸xU71��U{k�>��T;���_�0'�a@�W�MB�1z��I�td����\K��&�٧>mq'�p�/���`�R��^��"��b�8�\~��w���}s9���U���"#��λ[oo� =��%ŭ-��A�:�ADI�$3��Z�x�"����z.�\+wB�sG&�x���B�2�#r{��~o�G���#�Q�-\�k�L=��$������,��h@�+f
��,�`�>����j��l� �O^5߲5��O�X���f�7F��:4�{���/�c�vK���7s��ͥ�ʵ�dY��8�[��J{k���9g���N�anw�������؍b-��{��sP?\�`���Ⱦb.��6�(�*����)�%�0�Ͳ����}���F��_��J�E�QD��3�k�p�?a�8&L�K.
�p���h��hg�L�b��O�;����Hx L��2������w�6��	g���;�?�~��y	f=z��^�4�,��m>J���o�v.j\^�dM`2��n�n�Z���.|׈��XטE��y�r��
V��w�.%!l�j��ZC$��Rȡ��Ж���b
b��✠F���G��H]��V���qE*��x���rtI��0tcq���r���y�:��q�r���#yW����%��&�j��Z�8+�&��_��y�1�m�m��Y��?�,�1s0��Z�n㥽�e�R:N�5�r48��͟�S:V�wbo��eN[%�RҜN�TĀ�m�����*�&�_(F(5�tv�V��ތ$u���FS*:�*tJ�s���؋ S��+��h@877ј��Ь��4\�(��B����/��'|�n��?��c���1$�op�L0?�����k�!����{gf&B�(@GR��f-�N5B�e��x�Tjo�|�I�|�Pc�9�-�}'�"���j939NH�մB%�/Q|[�2�"A�%�gr]4����@���)zs�����u�1����`����7���M����.Mg��Z�����az#LG�(/�'Q0�n�����ڡY~��25U�^V��T�^'���Ë���3r����q�w٩ �7�B�+�4�d��^������ǝ^8p��瀜4I�՗�#(�Si����\("K^��Ô�њ��J�^:3���ќ�#레`���� Re޽����3Y�1�Ȉ��J���Ę����:_ ��4\����o�ρ0	9pk��Q��o�OD�]l�5��i:�������?P�E�K���聘�zK)��%uOj
�92�Q^��H�j�ől11#�T�쵆�'��*k�6�0sS��ZF�>�(	��Jk(��~��Uzs��6^S.SZ���)��[�u�yk�ȇ�*Ղ�^@)�扼.��9o�r��F�S���e�xH�gZ�Yɥ�eog�Ҽ�1u�u�.�y�G�8d��2�(�� ŉ6sy������W�:�vF���6$w��R��Hz�D�l��C8�j�I�,�:������a���۪���ۚ(�>����	f�c�H:Jc��_�?� �		�!�qqtp�klI!pr��6��1�#U\��*�lN�KD7ݳy��o���0��O`8r��z�f�!ڗ�$��zy_�^@Q�:���J������W�c:C"��M+nl����>��.�ƺ�'��f�1��p��s �z��B�}�)����.Ր��g�!����p[��Tl�E�v�;-
������}=A�����nq����E_�0YnMY5�	I�,5�P�MNd~��"�߮��2��
m=&���O�����Y�sފy��1=x���V�[�d������z��X��o�s�Y+�^~�=@���_/��et�N��׊*��X��4)��7&���.��U��o�������d���QV�ӧ�MXi\I�`��g�}�BU_�B9�[��H��N�t�Q���	�ʕ���<
��%��c���ׂNb�5����>	��Kby�=ȸ���o�6b9��3��IR��8l��S2#�~s��|�t��/u
K��=P�����v�� ɸ;��}�myv���^?���5����y�ًgFECނBm{!��/������Nv���^�~�ޔ�;׈�z�pTH����i@���T[�93�^[�C���D76��%����/G���%X@n�����r��D��pL�^8%��1w��+]}2|cw?fIL���͠�;{�.��OG4�W�7T>0K~���n*�b>%����['.���R�Yk�j��n������`-��~4�|�&uxFR�����.ً�+�j����@F6�,28 �WXuK���.�ςX�'���2�_A�)A�(3�1���+�N"��ؒc��X���nѧJ
��T�91�tt��۹:��(E)�v��S�J7�9v�y��}ˍ��T����ƍ����w�NXZ��f �i�W�
�m�gyCqv�)��b<E{�L�j��qtf&���>ĭ�����	)n��&�#�G�����L��~SE��E����ݏ�z�y�lMʥ�~���N�M��hl�eZ���D^�#�뱻@�xlޒ��R��s�9�.�mC~B����8�V0c��o0�D��� {��My@��2�Y�O&�MF�C�B���.�?�͏��!bL���rV��n'Д���qH��]�9�?��Xy�J�q���⽯�n��&���=���Ņ�HE�ǃSCH�K�0�b�\�b��e� ��{ţs8T���E���^ɥx�0���n|Z�7�L&|�y�7��k�t�D��_A��Ի+�2���'@��a�L�5��I�^���v�~6@�f�d��U�q��T��[����Of���0`=�Z�!��Z���C f��/U'�e�K�j��
��V��кԤ$%��]�'�S�R���c��v����Q�HKo����6���)ӧ�7a��'����FI��9��D=������4��?��V�r-���r����L��L����*'���p���8��ߤAb�Ke){QJ-ŋ$T�$�c�BL��_��:�LJ���:�1��?o���e�+wzRAFi�ͥӐ'��%
 �g&u�02����#A�6~��Y#�_�`B×M������<��2��-�w��A��4h=�'��^>�e2"R��2�ۛ}��`��
2[4\�Vt�}���ؔ��_�0��_�}�5�R�Z��e�[X���]ׄ�c�0�V��'�|k^�����1�g�]||���P��N�j�;�t��s��I�'�`y��H�5����C1������FA�+P��Tw7v��?+	~������+d�C��U�`S����~]"�� ׌��HߏGY�*d��T��4ػ�̠e�2)�Ӂ���w=�ݨ������lg��+�ֱ:C���'o������e�m.�WP�i��빋�۠����(e���2�����*�nL������h�y��c��7�D�Ŵ�Q�����N{ ,���:V���6�uO뤣˸����B�$3����ui@r���ɘ;)"F`���+�f������t�����	���=��B���4�<���bP�F�(���e�*�'����,\����^�����70J=[u󞉯U�`AIٴqT���~���7v��0���n�Zm��#q��)._\