��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ����X��ߍm��zѨ�`�ۇSw�����g��.��%M�:׀��T�����|�n.n�W�Μ�v\"6j��V3����W_l��ϗü��¸���ꈰ��R/}���Q�)�4�#������d��� �ɪ��Z�%���mT��9��T�3׵������b���|}�[�on��29�#p_$&YY>�m������s�{�R��L�=�S'1b�a�%�x�~�
sq��H泥3m�$����iY��G�1���YK�8�ڰX{D��I�����"T��e��*xY�:����KQ��T�}�v�����ւ��t~d�������*���Is�[L #���!�6o����V	�O����+�n.�f�@�Q&*��!^;"��g/�{�"ܾ�PX0=������/:�NF��Yj
��
I�k��K !�i���,DAA�d�xYT
�t����!I� 9¬�펦��CK��Y������._�����2�"bCN\禒������,�EԌԂ���p�����&�NQ�Uc�DV�]���cYZYn��э��S�5�hG����Z�'�Z�֜S�i�E�h�0X��|�إ�iяD/9N�,�BmOiEm���2?��u�E��pۍ�"g�:8�#��%���Y��tw��N����x�j^�!0���M���*��������gf�\� y2-����u�ip#+��kS���P�Y�z�`A���/�c�å9Üv[=�0`��y�F�E�$��2X!�d���)'�x��%BQ�A�*�X�4�%�Y1�����|������؄��J��{>�>��H���&�A�u9�W�H�*���~4�A�4�oN�mP�Ǜ�#3h����*�k�?�&�bV�G L���m���;Մ�% �.��8�Ξg�����o/�IA4�DhE�
6�������*���R�m��U�^�w�����^\�}&�s)�:rBQ	���������~]�Ě�(�Q�kE�uO2�o�w����؉�M5���]��[$�w�
������3�*������|I��/�3��J�� �o�*,dr�璗 �x�;S��kpx�uܸ��E����^:F��/�T�����L\�)o:L��G�F����9��Z=Ի�;l���+\Ͽ}�ZXM,�#R���e������p���[(	�ni[�@ ՚a����������B��b��k��6"�̯�|5�Ɨ�����AA��yǃ̏��i�/���,��A;� f��7�YZL�^��;Ppoe5�c64�M�c"qP�����@�N�	�GŻ�tr�k�= c�ixc�i�tTn6��3�>�]��Ĭ ��&��q��"���ͫ���0���ծ+ʕ3�3k\'C�Uۊ�%^�d�l[�^es<��n���o�I��<f�(�}�h*��?�n���ZBkq角�d��x�����̏*[����sG� �(p�=2c&+���WdI����������4m �E�e���Q�:���@��j0�B6v&�˙i��-��QoV�������H��X�2�n�E�j"T��ɫ���w���Riqv�mZ����7�{�Lՙ+�!Î?p�{������O:��C7�w�7p}�yn-$rj�C�(4�Ҡޡ�9}��ӍE���ߟ9~��Yv�4*1����j=1`��[��S>��'r�w� �7MhҎ�_,AU~���3��͏�:~b����4����WC�;���o���e�40�0�sK�Jk�~0ٌ���w�i'�ej��n5���n_įs3���k��=o����V��9��#�#�@�13B 6,Z�{2L�JQ9|��8%�N�F{�U3��z��^)�N��Q�y,���
yY��!}��-Y$�Ko�-:&�|Hh�]"�}p�wg P|c$鵡˶,�7]Wj��;J�_������M��/��#�����N�:t���)�I���t�{�4��S�@=ls؝�<����C��,�j�W�z�E&`J���	!�W�U�&G#����t����8�*��V7ҿa���'�7�qgh��$�G��.���s�ξic�`L@��>�CJ<p]G����m��.Z���j��2M��蔂#���o�#gnɝ�}�ć_��ssQ��g|D��������D�߃�������DA�a"���ڟ�jUq�~�����-��|Ʉ���=x��U+m�lC�Lʪ#�F�bP�e��M�6��{ �~ͥS�k%~n�|+WmQ�K�]��Ǽݞ�#h �Y��e��(���QP
E=,�e��U�b{=, _�%��V("��;T�4Ta��c+���/n������ezNq�#�З2n,���G�ԺW�'E�����B[ŭ�����r@-�#kA�2���]-�G )݀xw�psF~���i�xp�KkA�����@Ц����G�A����g�r+2�5q�P��Ѐ����\M �,�2y5��9W�I�gy@3nˡ��-�j�d΂�@"�S%�1�&V�D;�v|v��U��'�sW�m���=Q��O�� �����rU H�T��������Z����c��3F��k�:��[�_��� &�B=ӯ|�fEV�K%��$� 	���F�bT�ĺ�"����_ke��uAA!k�����d���ܨ����}�5bA��%a��{�c���(Z����bР�� w��<ʴR�:����p(4�Ooթ�"���k�x��{��'
� �l %_Ŕ?�J������?��-4]n���_�Ӝ�=
��p�Rz���ӕ�c����C���1����̩�V�kHqr4��)�����Qa-�sw��$��cd��j�eDv��=�c��Lxx^�F���3���yȒ��+��)g K�.�K��{E����1�N��ZK�B��J-���EM 7�٣��Qw5s�S�muk̺�������E�J��U��n+z`G]cNש.T���^��g{!��'!�#li��E��!�)k�W���+8�fl������.���!ap�5�Ų��q�FY�/��^��6�/�,CcFs��-�1#wݬ8#�ǯ�����C���e����lL�G���Q��*�DѻB�%�i����!^��"�#ay����ҏ>�B+gޤϭ�Wrq�M��nTi�Nu���1�� ��F[5�k�D!��U�eU1���|ӱ���1oAX�d�oS4� ��� $������E�w�f���P!���QtD�e���R��/�dC�7�U�� ]�o��΍��c�a���g&����r�	�^6j���H\��|:��m�L6j���Y�����Z-xo�mr��ُ��,���;hs�q�0 �s7d�`F�͹���삤1:9�P�s�b�
|z�9q����n�G-t���5�3H��i8K�!3v�U�`- �I������VJĥݘ�$-̞�{̍�X��[t�ʹ�p��*�Um���Ѽ��/�z��a\w>I��1LМ;���c�t#����ƪ�!���|���Ⱥ�Z����h����=�UL��#o^^~,t�[}��D����]/�1yȋ2P�1��a�Z"!�=f��L����D)TƃS�pW������I_X��m�P0?��N�����i_pvB�{����J�t�N7ށ4�#\���~�bF=n�zW��8��(-��d�K��*�̵���6=~�_̐9q�M<�C�y�S_|��Y�q��R���e���<5ݐ70�����2j3�I���R��������}���25Y�p$,ҳ����7������i�4`�j�N��zڃ��?/
ξ�3���D�͓�o�,3@QX�����{{��%�S�o^L��g�L�
ހ�����I��n�Y8���'3��s��өꢐ�و|f���rxE���o��6�H�Hf����d�*^��0�?�I������/����O�f)u��o��T{�휀.
�=�Q)����vV��e���ܟfyrs�0pG��0�b���@�M��\�OU)#4�ዤE�/�[�~����oe�#
Х�"�a�������甠�\��b�V�ZM�pk;J���(�H���呕X�ԠWiaPj��֮��P3T@_a2�r(
-s�So�g����n�JR��=/�um?����{�-luh�Hڀ�:ڽ��� ����b9�qE���i�k�d�6XjqX��Ś)e+b��ۺ�T畝�"hW�3�(��n�|�@.>!�x�<��{6X1�����Fu8w�mn��@Yl�m�7w�N$�^�F��𘰉s��\b�S�Լ�d-Re'�����z�Y86 ��TX-H��?�n􂾸��I�lk��1je�R��xH&�K�P�
b8?�"�"Gt>~U����x��	%�+���c�V#㢶k��E�C���m�
��G��vkN4��e#T��:�G�G��Lo?a>v�\8���B���;��?�x���I��GyP��R�H�S��Y*�J5l۱�ec;����2>��b���!��R�3�G�����M���<'%�
$�~q)v�ਙB������`�11V;�Ob�m�y�W��S�ۗ��U��W�����4���{8F�O�
|l�~�2C��D�|���p��7b+��O�7h�Olt��O�<����:vh��x]F9�!@��T��)�_�&�mPe(�Zهo�3��l���e-VGo6�]yi��V_P-��Mtq��Cv�*���>LL���WaX\U#y�;�h�9��g�O���j�L2��dnƊSs�:��<����
F6���VH��E�� d;�i��_�o*b
��2�m=S�*�0�
J��6��|�$�TV�b�=���Jt�����ٙn!��4�[��߯�7$��Nh����\�l���F.T~��Kܔ��XM�	ܭ�����(�ߋ�o,%X�y-��A�b;�l����RT��#��?
V����=U/���<��a��3�ؚ�r*�i�>����U 
��R���#���e& ��WL��lb�y�	dO�����W_�r�0W�$�[ϵ(��1R;2��x����n^�G��k�_��] ��T���m_S�ǜB\$x�x����v���R}��!up�f_��z�k .!v��Gvy�ꞥB���r1}t�jD��NQ�A�;�lP�q����	�%�n�a�\�DiSF!7�5Tۢ�G�NߋU�M���1���
mէ�'�í�:_��D�e����"��l_��Զ�8oo]�p`kӡ$��4�K@�nb��p1�'隣h�����.!�*%�,$��+��
h/�l!��T7�������Nv�Yy�Qu�^7�	�-ogC�	Lo$bX���0����M�Z@#
�}k��L��Y>ȸ�S�OK��^������OߴAS�/��ʜ�*�2%=��z��j�v3V�g˕Y:�3ߘ��	۰dPǞE1)��g�ՃK�[���޵K�0ZG[՘S�<n�ier�(r�5WOo���a �gJ����p�N�/���c��QP��d�uy(�R#��?;@R���s�$Ob��9.L����\�7��m��G���QM��� .���J(��l+�ы�L�=�tӖ�&'�c�d�r��?c�z"`�q&���*���L�Fm�2>�+97/h�L�1�sFf@�w��x#��?Єrz�k����Ǔ�+Ϫ��ڿ��/���RB�?�Kq��*q����5`��G���w1��^�Ճ;4j���$MT�O�BS�!E���Ic��A�"������i�7��u�Nc��h/4�v����l�Q$Kϥ6��Hf ���� IF�jnо]��PL ��[SK����Kx�&c�AUp ��Y�>��h�5�ky�l�~�e���ϰx�7���P��=�r�w��XQ�i34�sG�@�������u�j�J$_�>1�|+�x@�`8���Z?�
�MO� >�E*Ғ��6�Ne�@�s�Ġ����gqaj:lv��.�ډx=�J�`�|1a\F}MɊS5�d�k���.P��ԩk�FȈ����[0�gY8mɬ���� ;��R�+P��L��s/�mT`!Յ�^��ϊ�d��l,�� 5�+��ӉT�A���������8��m;_��.�㉒��=3���6�����u>����4��a�֌�ӭQ3�z�O���ZcI��-���i�W�-��Lw��6��O7}ѯ ��}��l.�Ba�keY�r��R�K�Ҷc���$|���?I�MV	5k���!�͋�MO��9�;Mq��Jz�l�	������,���/|"���SsB�[��!T$�MQ��_�ܤ���29O�V�>���q6��F*`	�4| ��l2.�OvU�tA�������2�kom�򼭱ڿ�kC���$���N{i
*���n�8�'�$���.G���0<o~�xQ�pd���U8�ǦnL\����6r�'�a�$sA�{e�ö��s���1`�u(2�YD�8>�T.ё��.�Z5`�V��g��ߎ�i���k�Y�p �\�%�>�����b�l*e�}9����`8@i�HP���۴��	��t\K��LUcU�U�+����j:L]~M^4�$((�c�)���n�*H��C=�/��c�����;��ܴE"v��� ܦM�8LZ�S�%7���OqE��6�����1"�P��ga�-[�V`���6~��&\�7��{��H�d8��cT���y$�K�����.ٵ��&�~&^��������	钱t��_k0[Q��H�HIU�]a#����"���S=c��X�G��vt��KC6�z	^=}2$��8��/�*��B!I���zD�vF���/�
�ˏ�wzfj�����q�%S��?��.UA�&}�^&j5�!�l�#��N\�r��2$%ҳ�P��2@ǱP3,FV"#.���$��,�B�O���w� fC�ס}5�o��ˎ3�a[�1���GL2�`&���H��u�$���f�Hb82�2<\��c_I�9Vr'�]�
��[ D���V��= MX�l�|��G�2�'�v�^&'�n�S�Gxx���wk�E�]"B���,�u�Z��t�c�H��$4������|��A���.���W%n@t�fb������y�K���W�wy�xѣZq����@��܂ﺿ�G���RM���U^FѨB�������z�yɵ�4�?�� �m�(���3=�QiS�rѮ�L�&�b؆v�f�x(?��_�/g�yiifbùGI{��6޵��:�BC=lj!w��O:oa�x0�������x����-m���,NMt�lYCO�'�������ch��O%Z�a ��߿�9α�O��9Εn	��g��4=��n�9F�Y2��)'d##��E�<*��� ��GW�Z�͹���L��#��7p��5ֳ*��_pD��<��aD\��L��XD5�S�/\�nֹ�g8$Q�0=Mv՚��&�"9��6n�ԡ���?�u2}O�t� �+��ۨ�2�b����LC�4RT]���C{?\��tU�d��׌r�:/���}%�vq���΀�W�=�w�[�r�7E�T�יy�O���ʬ 7�6��ޞM,�6�+�2�X��y�ۮd^jlۅ��m�r�>�1����1|�U�� J����n� ̹�b��W5��(�m��������a"����YQf]cQ�`�aD�9m7f��rء�;��&�d���H�\�K@y70���'R�4�9B����Hò���I�5�K��b>Ƭw��#d��O����\)x��6 3����R� A�5SP�`o��f�|��P�z9�Bx+�T����ߑ�c�r�@��u�E��+_Z*�Nk�[b���K��Mr�!�4>\2�=�hs���L�)l�2Q����7=���>��P�4��h��;����3���cӡ�U��]h��vp�Ӟ��6��a�E���m^�M�/P�[�A � �s��;��O!ٲ$���x���*c�gc���q_�P����c�I.�fe��G>��B�T&z�,X1���*��U����<���=gՆ�#�0IO`36���R���_�>���S~�F��J��q�����s:�Cfb3��4>aw^��3_5}F0_ǔ��ȓjܧ��U�Qr��u:4/�|�Gk��ؠ��������͛�6U�`��KCmwR��!���_)� ���-�7!�g���,�26����B�Tb�o'����XIG�}�B|��R�@�I�P{�n��h)��ގ��"Ї��OX½�-���n8�()����8Hh��"����KB�cs��D~/�\I@`|/�=<�
���=��W�$�d�̓u�ïsi��WG'�ͭ���?�����/Q�dj6�
�eQZ@�;x���	+�	Y�:����4,�,2��	�_˹LJL_\�� )t����D�,��t����F���|��.�Գ�3^I���Ѩ���H�C����C���Ƥ�!��p�A����Ɔ��H�����s���4��yv�s�"v�-�?����~I!���]Lu�R�VI��>>RB3F]��C�����(;����Ov%Q�Lӳ�����L�ZI��x�����oS�o���[�n��b�ߦ�������Z ��τs�1�)N�*��D$�%\zo:��u�G�� 'ǜf����L��㛑K-��S��Kx#a0IQ�0>"�CߚA�f����$J^ޓt�w�h��j�L�=�x�^��Jh��i.�#[�!mw��1��Cu��諬ۗ�C�ELq��	8K��`-b���`}E�� 0�I�	�/r��Gq�pp��ea :�ua:��##��<c���W�w|z(���\ Nps�Tˤ���.�Ȑ�\�&ǵiY�Z��*�V4�,�[Nr�݉���:46�r�cV����V�إÛx�؄�U+0�M��r�-.�墫��he9!،�	�����g ����Q��MU4u���i���3p�F�Ł�<WGo"�}0�$ ��i}��>k����`a����������V�a�9=L��0���1�VF�i>7�L�{���=���Pc�H3�����[ P!�����T��R=�~�V.`�M}���!@�e��|ܫ�}x��
�)E�b����Igux��E�C��i|�h�$ݥ���_���  3[e����0�@��?�۔����ᝀ�ѐ�4�Y��2�%��������І	nЂs��Sf��ȯ�F<y�����6�j��A�D�
�YMr'}�}<�,�N9�h� �/��W�B�*
Z
��ɩ9mP1�wՙ]v�je�bb��C��ߠ �����t���	b�$���\z��R�N�=KW���ci����1?x�\�O�k�A��D 9$RY࿫Ǳ�c�[(�����-ނE���ͤ�h�o$R����`��Vb��p�L��%��.�L���ݚ%��
�J��N����v���Ȟ~یXK&N.�9�:K�Ҕp?Y��O�?:|V"������[�ԐϚx�OkTV篜$�1�
P����osb]���O��Z��Uٯ��-���nL��ƒ(?�$X\YȄ�����_��-t�ʖ4�7�,��0�f�۲c�(���tp?3�]m`��Z���hԼm�MYHɩEԥ}oOq��6�z3����(�r#�7�O߽E�뜬��B����7J����&�s %�B51���*��jEs7?�X�RHXy���7��_�	:C����Q�M1���~��CF>�itA�4�q�J/YCf�G��ڥ�;K?�rǐ��{wC�V���(.�J8������B%4Ú�CY�v�-}&,�9N�m�Z����M!E1���ۤ�%��'Nk�Z�n| 9�g�N�;�L���w�0U��s1yq~��`c?v��q�V'гP�
�� �K��bS7������Ȟ����~�k��X������l�Fߪj���˻B��6���4O��:=��
țI��$�.��>�m�q��ΗV("�U`���a�O���y1��Kod�P����['�7�\ *E����Y���P����t�Ǝ��<q#0V;R��"��^YJ?�d; #%~��F�"9��6�2����Ĳo���]r�hsc��Ь�"���>}���&�Bƙ�n��hE�.V�P;�,�������K�6_p�D�8'ÿFЅ���f�Y<��k���㊖�S#@ֶ_	�B�R��.|��A�3��8}��D��<*rS���IU�����
��ݻP%���rQ�M�]jE!�C�1�X�_���ZZ�3CYy#���nHT��PQ���'���g���5K�mk�%Ӯ���@��X;��0�+�Ww�e�4|�̓���òM�^h�MisW�8ӧ�uJ�jؖ�a�[f�G<-��4rC%qOv�#2�#FH�����0�8�@y�!�͙����Fk瀱5�%�ɤ�4���B�u^۪Oތ0���VI0�η�"��N�@�&���|3K�I�8�ܳ`��� ���>
��VQ�{�X�����hB�[�5dи���^kЪ�~�Z��M�ndCVk������Z�Юbc*��(�C����ˌ8���6�)A{�Iw
�g�D��<����΍Re��#�`h�&F�CH���'���q���B4;ߋ ޣX����N?PQ� =~̎r�gmyf<4���n><ʮ�����WΡ�dC�DQBR��<�6\�.`~(<��߰;�^'��܄�Mm�m���Oԓ{��a����`�eR�2�*q�]��)ۡ�1��[³|�Axm�xH��p���	N��eaw�n{4]v(#?�t*��˺*�bX��v?rlt�;�$5Ά2���D��=0�_�`�"�f���#|�w��_�6�/���Hpʬ�̧�����h ��I�+g�XE�X����v8V�w�@Z7��<ӻ�fzƳX�x�1r�@�f�$6�����p�l��b����t�'�<S�~;Q_ﻴ�ʕu�&���߆T�(Ð����4ݩ�Y��9�g�7���� �NՋe3�zG�A�#��HT� #&t��h�bM63"[�b�ɂ ���>�����'����p���x_�K�:�E}BэA�7��Wŗ^�=�&󏉢���ܴ+R�|�p���メ���P��nz��<0��=����$m]/�_�ƫJ�i�紫[u�^�q��5�bf�G�ބ�F}
,$�k�����"
�wK�n�������.*��Ϣߍ��S��s�׎%����
$16Ycy�ֽ |��lÌvI��	��M����[N�'"�����up�٨�	}��?����O@c�/ ��Xe�e�|Ld�|QEb�}|�NW*��[�,.>}l��t�	���N�0#������~?��ySPzO��>�-� ��Z�]��g�MbRloB?�U6ty�$!6�7i�̐��_�����0�=�]U!��R���"1\���P&:l���n�`nu��M�cT����yy|�j��� �����>p��r6��͠�'QZ=eƉԨC�*���!�p5�Gk�u.��&�<�fR��J�1����k��T�1'2Ծ�*�fv擁�b�P�,r+��z�&��J=�0T4,F�ڬ��zi@���zv���x� �I< p�Jz62^��O��,"k�(-b�����
��l�؅���G�
}n�=H�o$�#�;�8JE4C�nc�̰���@ �'�@�3�7�X��1G���җ3��y�՟S�Az�e���ayF*9�n�i �w�+?��.��Q�,N�}^3r�1��NM�X]^&���e<��>K/S/V?�qm�|�&�3-U����>U{p-{�"�j*L؝�|K:P�<;�`Gm�u�3k\��H����:+�-P���;-������\��K�1��Q���r��b�[oI�L`�q��%�M ��l|�/Td�>d���!_:1�h-�5��n��*�{�M���ż�������x�+��gU�l�?���%Z����X�3�1W}�����#��1J3A�5��o�@�t׌���d�-��b_�K2����uŠK���A.͐���d�V����&a�dO��Te��l�.�8GC��kv�T�N^ıo\\�B%.�g|��jB��5��T�R���������^�9���U6'fAk��U�]�;���f6�
dY����>�N�,%v�L�Q|cC��[/���NJ�����u ��dH��R�U�-Y����Y��ax��S|TZ!� I��[P��~��x]�k�8흣P�������pp!��%H,��.��s� ���<�����XD�=���&�ҭ����Y$�ӥg�*�I�t���|;
����?A�j'�3�o���Q�.(����+�ձ���@�ź4tV@R|�~�V��33��&2����d+_,`t�����`*�ߛB-շ�c<i�ط���&�~ǳK�9A�g'Uq����i,��'�wpNiS�6�mMIO���TP��������`x�6-S��& �V_�[]p;�*T�D�h�&&�d�5='��g�ʌ���g^��+��@P�x�}���UiWd���5	� >�K���,�gW3���9/a[�"x�Y����G���.˄ߋ��,4������v8�I��o{��-�����O����寏�L�C���א��c�>w[x�;��l=���]�)�W��}��	��$1��T5��L����M>5�&�:]��l�1/xn�e7�F0�r��?��Y�h`�n]�wi�*������nR�,�x������j��V�c��8%��*�{-z�qr܄W�V�}pn�;I7���G����� )�/1��/2ΰ'+���6�taIB!�w��Q�6��*Ei��X��ȨƓ3��dma��
	��B>�pJ�+ P ҹ�U�T�F>��=�5���W��L	�w�cQ%�}���c1��!1�7U���)?#��UƂ:t|�#��nkm �[�&n�eBsw8�}�U��'��k�豑�%)���x	f]&���"�N u��Y?��icfRy,�ݷ��7����p��7����FQH�
#�Å�!=�gH�I�L p��n����q�EV�H3�[�_Hgz�?�>�m����tCJ�C4����.&��l��������M�b��:`�{H#a����:*���	����	/՗��_�Ru:-���9����3*�X��s<I�8�"��M�GЖq�\�ZI�"�E��S��[^�x�j�?#x�2f@Z}�i]*�rk��ڔJD@P+M��^�bǨ���K��nib���Wb�#s�
�`���?��6�#V(�@	m�5;�x �U�>R�;1���!�Qб^&��Λkc	� 3�&p���@��-g�0���ǿo�$o�i����,�����?oˑ�S�k� ы��ϲ���C�[]��DUU��`��d�z�ҏ���9�/����1� \�����a|}�y��*{�w�;}���֮<8��"�5&7^�o�</H�71G�j�K��>�%�շ۾Ӆ�-rO�Z �},S+i����%}���$sW���"@�:�`z[���a�^GBJ��3
]��4
`��Z�g�[k���Q ��3L��t6���h2�o�����熫=c���G	�F�MQc�͈j��9eLu%�K"��J�|G��%mVUm��c�e��"�Tn�Ɲ�����|�Jk�b;?)ѱW����Ue�en\�q�8n����V...QR�
�WP�N�R6u
��6���Q�њ��M�f����P+@����N���i� b���c�`�K��_����N!0I溰Y�U������99�Q��wJ�I��0Z���|<DJ�Z�2�ӣ�UΒo�F�wsȟu�J��ի>#�����E"*��f���<���V݁�T�K=h��9N!��c�
�F�� ԉ*����p���z�S�Ǔ�:��BG�_DC>�/�*��'�_�����(�Zj�jŌ/�a��*4���i~�3
�]�T���U�X��P��VV�AI}�˴�~e���&�E��+�����$����Y�]1Q/_-�,i�}J|���z��
x�����_�`�0��IZM�uº���W�+l>2$�<���U*G�KV������F�a�\�����ڕ6�����تbV���q,ۇd,���G/yg�����߂a1pK���2%��d��M;�?�]�H{�����#D�2M�֩�)sf%�J�J	�Ec~c�X?�.N��g�V3(���U8��|p$�c�ҙM��v�kp�4LL�׵��2W�M��@��&���|@�H�7����~K�M���� UkQ-Օ�}Z���@�v��~�*]�)
Np�����i5dx�.��e\���� �"��=DP���k����3�|�<�X��b�IN"ci�#���U����M�8��$H�f��&�퓱Ġa��S�9Q{��<�5�B�)�k�S�]2+��19�R��x����EB5ϢoE�)n����7�赆O`��sr���a6�����)�1٣#�=LX�i�1"Ӟ�ɦ���h#:��(���\�5��ہ�}!���6Z7�O��p���e��H��B���=._�h�42j��5��w4T��V�i7�d:<�*H��8-KI%�J�k0�>E�� ˷��i�i��6v?����0�݆=[�aF�5���f��G��ќBs}�H݅�$(n OúK=�Ǖ<
��A� ����}g�	::">���Y��.H`�#���}h"��������晶[����y��E~����4fY�UO&''��ؽ��*Xc>���KL#�)vKp՟z,���[Ӱ
��F�c�3򂻦"~�b˂9mʡ~��KZ��.�� d(� ��l���{�(��iZ��-D�R&N09QdlG���F����LPk��5�i��8_�l�H�����/5��tu�^�+l�%<���Hu�cF �pnt�g�����܏���;WM�v�-�b�o�	��wcm�p}��w&��Ġ�#�30�)� �e�A����ԓ5,�ظS��"u}K����`ڎ������7G�`�_� �5E��6�j����-��p	L�3$5��P�!sa�SV? ��/��V���3j��}J����.XW��� ��5[�=�)X�R�o%,u�U�L__C�|G�,�N&Ua��G�9��'����jrR׃������}aܽʌ��e[��
\L�i�-+eqI�� ~te)��B\�N:�[�Ǒa�G���Vo͗Z�m�3�{��I�p��Y�Ҁ)%�����|��E������o�M�<�)	�����5���<IaB7D"�\����d|F6��<*�V*�|�E�;:�w�ϑ�ƻ�S���&�V$*�쭄`T�:�nO��9��d��'���A����n��m#�ij�b~Α�u����fc� T�>�����
�F��}m-��~ ��V�`n��#b{��S��L��]L���Q�4P�s,B�'&�wg��1��?��rA��3.V�_�n<Gh6�v֎���<�pa5�/kǶ��T�1��l�"1��4��	aNa�r�U��kb�+����v�~�	1N؄Ơ�/�\�pg���V����D�/U�:�D�y.4�S�A�=�b���]�yd*x��	�G�$ҩ��9&�I�,�E�d&/R]�,gʃٖ��Lv�_�\#PԮ��`���xs�kʸ�c�Q�գ��È��*�$�iͼ��y����g����(VP�`�U߇m��=�%�����VT��zͽU�ջ�6����hA�WI;�Zt�|o�pO<���� ��Xk+