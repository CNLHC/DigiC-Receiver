��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���P<�%���>�e�2�H����^3p*�ˆ	���<���ꂸ�V�8 [���.��I\��]�<(H�����$Ϣ���`��7�o?�_��F~,�%���o��s����ޑ�
x�AWG�[����q��-�j:k�U&n'�ͣ����^�c����]]w*��6g; 1)A�ΠU�_D)�s��B�<`O��miӪZ�^ޚ[�&&��^ɴMɕ�`�6ڃY��B]�iU�[��|�3>�d��}'Vbۇ�_KJ���H��x+ t�>����}�=�֑Ǻ�L�S���Drʣ�=��3ƜA%T�X:+����S�f��XvA�k*�",o3�wv����T"	@Ui�W���\m�����_�0:]:��m��V/+58}.2c��/��!s�K����;��-C�j��ġ�d� O/D[��$�c`�Nn[�T<l�E����9�y��Z��M���0*% �1�{�;�r��3	`Z
���-��P:�4�Q՘���#\�'lD覼��V`�ZЄs/";"��d��PX��<y��/Nkc��al��t��;�|�^���c���I�zZv������(��܋�c[�,��p�
����|Eb��hoT]��bp�i;�\I������0D�G�M��MV�Ja����u������45�gjPf���0�޶���M=�&ޏy�:���񜝰V 2��]ך?p������n�%u�d�,�j
69���T_$w6��&�?�Rg\�.�)<z�u��zu��(���}D�\ ��j��a��t�f���T���4��h�5�O(���m���Y���GV�	�;?�������rb՟�(�������	-�:��%���ҐŶW#��_��s���z�L��Q76'h����$䯢NM�mK}4Q sB�R����P=�&,�M�}+K��_i�G�vu��J ��Ɵ�I�JP6$�JPR-�e��'�d��)i���URۛ�į����/��lE#q�Tkv�Ϋ�6�	e���Yk�{�T�g�1�uKK����c!�A�Ҳ�r|i�#g��9��lF���ٳ^:]I��������I�?QyaYR��h��A�J\W�\m��M4NN/I�mT�>�i��+���O?�²7yx�%�ҽB���\xB�Om�=[�%Me���-����ٜϛ�Ҍ�cM�«�S�E��0�p���k�e�FMZͿeW�cV�֋-/�$3�6����z�9���f�Z)��F,sSAo��6�_���E����MJP��VHQ�|���vJ���'�kF��	�.Ts@�-��?8!��(I���,At= �>5�Ҥe��C�i�����k��z�/s��Yh�� ��3�9�;Jֽ��Op����a-�=K���*���O]^e}�='	�T��P�z�`�b�_�� *�G;vt���K��ޓQHMrZ���BK)T�mb��~w�H���m�#��Td��5��� ?��z��Y�d���y>q��D*�ýx��b>��g	2�����j�+Ur3��F�:ӎ�[��;��q�k�l'oTM��������x�:N?c�ʌPv�	�m'd�b�7f�PB/�_��]z��)�/�D�fb�V�q����Z ��^��1g�k�	|H�ƼI��e�?�]<��|�Z��	�������,(���Sx�!��2V�F�o=��&�4��+sx�����^�J7��]}�+8�DR�R	p'��.�!�����,�S	1�X��|N_�R~�"��U�UF���N�r����p���3�T
u�/)R0O2.C�@���{��[l����ӿ~���P�c$�9}nd���d�L�e�{'c�ۉ��8�5��^ᑺM]v7p.���������DD!��y�����X�1�Q�Լ����ڵ����y;�4�� 䙊Dʄ��8�-%�1-+4g�H5]qt�[0����d�|���S�o�A-^�{m=�n��Ɏ�����I�*��M�{�+N��G!s�4��u�W���ddAj����j�˖�{þ�������d�bo��S���f�C?�$h8�DӋ�,��TN�{>�o� ��c$y�6!{�!��B�*l�ٺ��E�W��si=n�"鑓,�@���eq!?�ܱ�-�e��9�����u����E�ON��5#�U�..��pɢ���Bc^]�k�p��a���u�.RJd��IӞb^wV��(~I>Z���D�lܮ���A��Z*S��������M>#��qY\@�|��`�L�y�����ީ���j��<k4�����
���H��t�����
R��fK�����R6{N�-���9N/i�&�b��F ����v�;�����v�� �?7c(tI����H�X*�ւ@
��v�]c��\�u$�+-q5p���W@!$S͡^znĈ����0%gj�RC�O-���y�j9Y�����"��琱�͑, ����|>>^�aLۍ���
�|�U�
��F�5>�����a����8|���B��W�95����Kț��r-�,���*���ި�{A "u��HPq3k�uO�;8F����1�.8#+;iߕ����PxuM�6\����Xٚu��̔�͟���&|Qt1�����$r�4 �ܧ�`��s�H���]G��&듬k��(L���3���sI}q���C1�Ϯ)�YpP�U������0��T��(ڳi"��5�b��\W�nF�ph��N.��hzHAYV����U�����y�����-p#���4<��B�t܏�-xQQ���Z��j�J�\���K�E�4k��H%[��*��f
����z�aF��Y��׍�Ȧr���q��o�RF�Y�V�7��dG=����z�D��
�|l��$�yB
��2B�����0�H���V�[>�A��(w:�u��Jm�҇��貶Bf�F�ͺE:�3lȲ�.���v򂅪���ۉ��7�$+&a_E0e�{�~#5&c���B
��+���ĝ�)��}�޸�b0��%�!Q?>t֗��is�?���O0��oc�0�7LHV��iLG�Ζ4�a�@��Xl�0ԌFOc�@�f�̝�����]�B1��ŁE:Ye���g���V���u3d��\�G�#S��t�`�_�o-~�����;Z�d�Rɛ�q���Ӌ����U�R�60?|΋Ԏ���dX��F�^���(�''\\N�@v'nh���L%�Il�L�ca�~�m������e#&�N��7C��pЩ��i��w�m�bO���O$<<a��m �c��e�9�4�ۊy5��=W_Mm�۟�\è�cJ8���3�(�`�H� G��02L�9~����υ���VP��N�z��=n��-U�}-��8=
�m�F�(aF�F��K$��~7c�{ی@4�
��NΟo	����_�ѭ�"l!1�w8�ar>�{��^5w�U�xmF�8�����jx	�WF�]U@��=�h���]1��;����#'�����r(Β~iz�s���
P���oZ������S�:�$ߗ�j�(�(8=i�����z�d5�m�rb�a^����"��J��b���'QA[t���V�qF7��V9FObI=����Ⱥ8�t۬��땰�W@�Y�ũ .�ʋS�<L�4�S��*�&�f�x㤙��]��MײzV*�p�w:���=��+�{����G�Bٵ�O���!P���M-�M[�J:B��xKL�����A�p�c |.&�l\���
_��<�Wga򻲺������Ϛ�5�� �_�==|~�W��Ʃ1�y�<�z��%��W4�w�Yըn���*�P�'��F�p1X����XT�Ji��*̬>L���E&���h������wv�yI�n�0�s(��FU��c]I�\�!�P�MK���$�V���T]��A{��>�׬2�T���'��5a����B@�2��9LsbK�T~�� �R�����Z������-$�_���vC_�y�G2O��I��E��c�3C�?�&{/�������Joe	k�Y�%#�x��Ф���]1Apn��o�(�.*�|T�RD���<�:`���݆88�L>\ u���!x�@����v�T����bP��,��~??�^�Rܵ)�v���Ӝ�J��!�6Q:S���ɹ���"�r�{?M���=֊�<i�(���ϥ�|���=G�IX(EO�Yn�s��&��c�C�e�K,�����N��E)����;S$0f��Xn9���h�+���$A%c����^�:�s�9{K�ס���
�\g�A����JH�GŲ�/�8O�������`cN�_$B�A�UR�V-���3"��Y���@�I���x9S����"]�e����iB-v]��a�6�:��H���	R�|؆q������l�	~�O�{Rts7�-U�=�u�Ʋ��y��<�A��*mp�|*.F��������e+B��(M����+���=~�;�m�%oD+[�
���%j�'Rn�xɍ��6���CZ�#y�X=SrÔG����Fcp�-�pR�A�:S����`�Ƥ��\����V�/�u�$�s1e��=O+C.�}*ρ�f,�=���S���?��9��'�ɠCbָ� r���{](0�GAA��<aJ�+d��P�f<-OD��i���i��z'��i����!͊�ҫ_��IpU%L�ˑ�\`OLQ�"V�Cڻ�����@6�`��8WZ�t���7	��ǾC����-+SE������xK�AA���J>�ع�rZ�\�9N`:7wX7 �3�7th� H��Q�w�]jxY�vm��x����aZ�$8�]<�1���b_�N��V�	C%����hSzǠ�u�K:T��Q�`nzp<�JF�^�0�E]��i�v���s��j]� ��9NH�}Ҋ����Fnt"m9�������VhF�7������o���%�BcJ-���a�� x���T��B|�}�*>��� ݮ�g�NF_Wv�/��乿�G�g`�v���0[�����mt�H�zjR ���u�]k�\�����{78��î��|_t�������~l�a��/�n�q��𤔼���O��,w̕���b	��I���fQ�����ﰢ��o<O�A�*����s�O�wѶ� V��,c!���(�՗��� <��4$x�����>ty��7��-��u�L#�b�m�������^��+x�-�r.�Ң�8�b�z�Q|8��#�G�U�
}�&�cR鏙��S��y��!���IQ�v��@�hˢ���V.7>*�*|*� ����QZ���52�Jh�L�������.��݊K$&FO���[�5��v�-�~_j��/�k�2M�⡌�_���/Aș���?aR��{�k���J؅�In��i�7g���z ���i'�u�7����}p$h?��uW���,�i�7���D���q�d�D=<���	;0��H%��d����AڔC�񻍁��x��� I�y������bQ�%��[3(�J�C�c^+�`Ƿ�W�u��YI0ʂ��.^��������a9*�Ż����i�s�����R�ڐⴃ������%;�&7�/�!�l��-��,���v�n��ٜ����i2.��NX�E#Q/t����7�52������~����ƉPJ����ʪ;��"�O�J�2\�E��M�,�+a�U�1�x��H����զ
!LLd͚�t����&&[��S8%6ٙ/&���,͉ͱ��!�u����*ۼq��MI`���d��.@��9�,��{+a�&���@��D�3_@�����x6����`�|.~��;M*�0킑�~�-�D�e�O��Fg4��EʔC��{���kЭ(�P�PG=r��_��r.]C�����7���*_%�����Ʉ�&!	6i�#��`㟃�.�9�~F�����b�
�2�
!�A��)0� 0ςv�<�r�8S9�E�c'�v��J �����Sw鉏�&6�C"?W���fd����b{�_x��]ׁ&��ǌ�>�3w����U��c�WXL�$>�p����ӕ���(�0�f9(' ����E�M4~�v֯��V�F�E�#� 
	m���.�Rpm3�]Uc��r��b)��$���P���zF�����Fh��j�O*�ht^��=`��ux�(�3c��آ��$bu��.h��e�O]�sr��KkH�[����4B�*dm�+��#��jJ*����QL��*B˴�T���{�vva�P~�� �]ff���s�'_h���i}v9c}�z��I;+ps��i�I�X���u�a�S~[��Y2�u��K巜UC�#[ź��ҭ�&<��-�%[g�A� �瓗��؁�J��� -K���������wja��Vsxyj�!������\Ȕ!]�f�_DV�mH~�r��VZ�f3@��3Ό%E��ϟ��f���7�*�g#���5$<��*�iL*�p�(�MR {Z�\P���X�fȝ�p|M�#�g0�O\(CV��\�i�����Od0�d��e�=��"����xb]�G�=[����g�r;(�[^h���H���g(���k.w���ֽQIR_k|���j�(P�
.��s���r�����N���9����#dq�;�	�0Ib��eIG�}��@������M�aI��`	A�M3�$���|$��D��>���&�r�ɧ��~��>�՟`Ya�� ��;�qǃe��z��z��%6\H��6�'!�-j��<I9b|���+��r�	IP��ϊ�jv[d}C�دP��`/265��AAP]]��z�R�@B��ʄ͹3�q�[��_ic�3=��G���;D�h/}ky�z>�y�}����Z�	��X;< �kN��v4�Z؄��|>?s۾�3��N�G_ �2����=>��B�$[����������9���,E�8�C0q�wު�4̙�3���� o���ڃ�bǇ��$ϡ���X�����㇈���Z ���Z�ZӌJ5��~YW{w1�I�g�R<��d����H�ʟ]�5t�Y��[υ�!2.|]�4VT��s���$ȳT���i=��Yl'L�t�� Iݪ���}�׵@� �1տ. ���=0��8�\�8|���8��1BD���2������M��_�b*{PC3~~d���tFX�	�����߻�S�B(R�i�Ɠ�XF"D��B��m��
�.���ƺ	(L�I��kf�oB2�ӰUR*���u"C�6Q�[\����Q;ڍ��~��$k�yC�rVz��v�<H���:o~9���ѱL3�y��x�B5Z�ETf����abT�L^����ݕ6����qn�ͽ�Ȥ�H�]�����*:T�m�`�.NŮ����!�W�dRh�����$�*��ofzo�JE;8���@�>|�<J��gw	�"�h�C����g��R�]�mf5r�l�GPz:ɾ>��'$�_3�o$Y�,F}{�	,d츧�MF�^im�������F��2�n�}Ks�wX7+"��J�M}R���/70�RQX��{6�>�o���vݯ �bc��Қ��nC��� r�ñ�5IM��h�`I��bqqv�jj�qZ���َ��a�[	���eUw������%b�j�_Ú]<+K�4m��@?C���{���馥�D��4W����|��m0�a�� ��7�@�`~�ZK� ��P1������S�aQ�܄R�j��G��}��u����SԜ*�����	���.Q�y�<����<��J~����Զ��|IK�L�kO�y���EI�Ǡ(R�;z����������2u$�}~�6/����X�H0=82[���X���S"������?ɝ�d"�b21O�������ɼ	���k�wIn��g��a���K	ut^���!�>Rn�qH3�Ak�r΋M'l3���$s*���y/��J�F����]UJ��Q<P���6�oE�Q�����s �G��qKs�������j�
�I4��`#��baA\>M��1��{��!�F>:��8�$;)XE��j.��������`����W��鳘]� ���O��F�,��ȩ�$D���wtbm��D�-O�o�j0���i�'.Ck�E�"�J'���Ypv��9�4���[:�+���zp��&��C�J�=���q���{[�o}칬�5�����J�:H����'��19�e6�::؉��Xxe����rq&jp�]��������Vh����@�Ֆ�'��$�^DK�de��n�<��Q[��i٠r�kW�����i�"��ؔ���T�7�.��
CC�{հk�9��8Yr�u��7VsJ�B��u�R�l������bp�4����f�{�3�����N���jzH�n�'�5�k�x���or�E�]��iP�8���uO,�OA�)��/���-���}�$���8(��:��>�B�O�X� Z���Wb�����s��Fk�'"�c�j#�~C<��(���2f���TR�<�� �T�20��%�I�l�t����ӡrڌ-n<,ߎ�=�x0��'t��٘n]�9
�H7��ԯ���֓���~Og���.�d`�"�󐽠c���X�_�\c����1-F�d���ˏ���t�\��GϩK8�J*4�����_`�����q�]-��q����x��*�� ]��}h;�k��Y_���ɥFUg,�ibѢ�������#�`^$r��Q$����Ho�z��U��'�=`y�:e�1��
�
Ѭs�����o�"( �)o#*
�8OIh*[������E��;�x�Y[��*�!U7�8��7_�z0oQg0�����s���:���k��0U�%��A��I�Lm�v�����B���]&T�#$��~f���75�I3�a�7�>MX|����B��)�@0	~~��q����徫�%�P�� x�MhTU��t��oוS��=kW�ʻ��͙~�$���>;}>��D�tbV���� ����l��ݯw�������ʀH�������$H��w,ۼ��f�y��ц�鰟�P�d��.#$	w�iM!"�^���9</=~�ys4?3����m(���s���#[�]rd��j6�?�����:�2�x�01�	KG�Eo6�7�)p�+�@��V��������B<K�[V��kǖ�����D������,�f,�z	�r;�	�&0ֿ�S	2������"}�pF�Ϩ�8��1�ahQa��y�R�~Pz�Ng��{5K����(B�^����ͯ�3Mn��_'b!z��E����H7#�	�ġ7����]�qe��O�����'��qR8*9~2ʂ��R�>4�_D�f�����Q�wz	bK����`�R��F(���
�H��� ��;±�̑����T�K[�;y�cS#�qA*�7��t
nQ;^%�N���\��{JMY>��ġ�Z��o���N:&�h�y���C�q�Fy�g(˖����ƖrE��CU ����;��8��>^���+ŭ�	�������^���Fw�{�k�Xv�������z�@38%�]���$vleeb�^P��!�uguN7��.v1=��j�6��	������~��N���~���E��<L��Y��obi~��W�ջ�L�5�Qz�vx�S�i_��M��19}�z/�x	�F�jL�����`��b�p�;��=�r���*Z��y�D5��d��T�]��4N�tY:��M���~�A�<��h%��Ĝ
x���e��=ΦݲU�{q:9���~��Y���������<�'�L]��9�y�e�pP�X��Ϳ7�Ƒ혮*�HPtjϘrK�f��/1������hP=�$:��ܶ�	%��W��\����j�5����u0���$L��<k�´vB2��o��|���C��6#C����X4��*�#1k9S�l"'�Xrv3iN��}#)�b[�Y���[���]~�(�7t	�Ĺ���a��G'������XD��NY�������
��/BN���r��,��G��g���&[��r�2�7@D��c������1�$0D���r8�'a�G�WY�>����{��L ���䖬��xZ�����Jmq�b����'�c�H6#�M��+�#�g��oT���2�4�I�v�d)��7��Ф0ｏ������5�/�Oꁝ���Ta�<�ПN���a��7q��;��|��V�A���M��}���b�QW��(α�t�kT	V�#-&�R#��mNAj_���e�mt��L)�G�~B��b/F{���4z��Iy�oq�Y�xR�x$�Z�p�{з��'��wYA�B��13Jݶ=�P8��8?*{��iA��,���U=�F�Z�j��JV�V2=x�CHϸI����ܼ3-����Z�*q� �:�~�*\�4�U�kg��B��j/���;�l��ob�E_�C��]����%�Ͼ���K���= ��b�����i��P���r�b�tG�fٳ!]����#e�9�mk�b�W����`H���z@0��*˳���?\���^����������BYC���\���f��ebK ���Q飉ud���/y��f��A�i�O�S_;c) <G�� �]]�nI�W�͞h����#k�� �mڝ8h���Ѫ�o��QV� ֈM�!0��nf�ܷv�7F��5�3��9�#f��k�%���\����
$jq��ldn�`"�ļ�~ܓ6G^��ϼ/Xl����Ny)=��V�� @\y`��Hl���a�Id_�|Y�v�Q,,�ݘ�m:�&p�<C�&$o�+U��v|���IK�/.�����d���ʞ�Af�]�Ȩ����wN��̀h]!����6ݒ��}���g���5h���k�9 #J��L���7��U3�i�����}%zklE����P���i8�n�
!j�g	��ǀʵw
�y�?rx� b����wbn���e`Gg/_D��k�j�a���`x��vj�6	�U��ra��"� `�R���piLh'�?�9��)��e��`�e��j	�;eI�	�=�M�f�gV=4��<���uJ��/`,�o�D�E]*�����e�����<�e9��{@Kk��ڌ��*4:�!m��S_E��	5U����h�~�F����Fg���68��Y��~F��L�~�)��;������&R�8n�[h1ǘ�>ު�T�6�~=��յ1��:fR�:ړ��k�s+�G)+��v8����g$2?eⰍ�|�{4+ o9��P�l��BF,eKoE�BW�㨼!�Sy=5奃��ސ��ә��@)r�#�������^����W��W���z�dA6����ɥ3�q\I��_%gI���ڠ�p_��5�1�@N)8�r�{��6��W�.\ǥ;"�,Fq��ـ]�����X�;I�q�&2�
���Yٴ���L�'���YxVU�a-��N$���BO|����E�����%7��*"$�dt�wd~ԣ<x�8K��m��xp�gf���P�t���ɮ�twʟf��o�S�x���AK�-Mj)��Ȩ��	u��N�:����p
]ߒA�������T\X��P��o~��}fYX6��`��)ۛ���Ҙ� �pP������⪍���#p�bQ�W�|�2ZO�����?�n>�ظ�/��I;������j؋�-�yZO+����:��v���@�:"Ѩy�V?����$[e�B�'�|\
�:2z���_� �<�:#D��3�/>n��@�k �ɜ,��	�����#�#��yS����]UƩ�ԁ���^+[����N֮�1tT�
��Y�L����[w�3���[��4�Ec�\�O�c'�cdгK+@~��`���g =J�(��uxMs��ꊍ�>�$):��qtf�6FU�����݅,���K���� Q��0��o�h�͠p��B�e����E�Dqᑡ�﷓?��B���l���N���s"rkK�D�ܞ)�����n�@� ��n�'�Ym�E
��¶��m���$����yp�j�+ /禙���Y��IgΎl.��5��4)�T W'�W�VJߴI<�I���)�T����ϛw��[V�'Z����Ǚ8�֔��P�W
�`�<�� ����8�~��I�Ϊ�"|�!�8~3�
��'�u_�����������H�?������
^h�f,���;��Ehd� o���4+6Bn�6Λdȅ��d5̈́&��AB"3�o�0���u���+^�'�2H��{+������Ϲz��\���ј)�e�Z	5"�jb�dO�R�3�ۮ�-�j�|��	��[i���|���Y7�^|Õ�ƞ�;�𩯍/�`�Y��
o�T�J���y�[���������Ⱟ��u,��6 ����|�O�9N9�Q�<ؿ�ISY���q��R�K^:=�6���"C3����co�=0I��<|&=K��Q��UV��B2��п)׫ ����s��YRx_Oۣ�UNqt�&���U�>s��R��μ�#�C2c4�9(θ��x�+��hJê�>���F]���M�Q���`g���v���G��4��q���qhT�Z�8V��O�d���臷�O�i3�i3Mnvzc���#o�P�^g�a<�{��kBg)o�%y����ѯ��$$����i#/�oE�ڪ>U��������pP!�n�q?_�\TM�.E�_d���2�lQkY��3��;�[�,G}�����%���3'�T�@<6#8�Q��9+Ƽ)���s�PT?C�Hn������;�bu���J�!5���D��N Ч.����������q}�L��AO&�Ft��p,��aO�{��k��î�՚�7��{z,y���F�S��oQ@K�72����ڵ� ��L�K���?�֨�u,e��HC!�UU��Z�9F�r�q��	J�e��:qmvZ��" �� lo�*^��W��]Ǳ:�FջxF�%ƀ�0"��V�ɏG����Ǥp�΁�@ l�e��v�4�#���\�M��Ҵ�6\�Y�#�����$�]��O0��P�KC�����_�h*�
ɺ��.ʠ��HߏIf�'G��"��9�Y��7�lܐ�Qh8��'L?�A�.���d�0��m�~o�T���W}�c@�d;�D���A儅n��~��֘�'�M�}ąԜ&Ӏt�@��DFR�����;���!u������3Ãv���I�)s	��V�?[�y���z&7��K����:Tb��-q��|} F���rQ�d�0���P�^��%�^��>�ӮS�.p�0B��11ĊJ�9���L����iTd�ǈ�����4v�]���?m�H�{\5k�$͹߀
n6��y�*�}�ջ�G��(��jr����K��F�~hd�h�݁�˂Y�6�4Q�G�瓱���K�<�@{�+�DgbwP�V���Jm޵����m�M�#b�{�� Ȁ�u�?�ٿ�w]��|?�z7M�u 3AXH2�����4����)og7����᝼g��q��E��a&P�e�a��u��ʣw����	w�B��jƥ��r&F�e>�^����S��MT�wQ�+�KG~2�{	��BFn�Eh�s�H���)@<N�<{�O`�L�\�r*�n��r���p�n�/�O�NU�3c*��׬u���{���L�\��d	�.jW�9��)G��MN������OZl��`vc�ˮ��>}]�I�͆�}�����	�Ӆ�A�c��pk_DEod��GQ�DiJfa�:����3"-=�+C�^ɧ�d�8�)X�8�]'4�l��ԽUnh�7/E!�F����k����� yM���:#��{ʽY����]��Z�����_��وZ�����0%��y�5�`�	��|��j�}��r�Mm�R�Z��Z�S�dh�4mA��^F!W�լ��V-�-D�<�����P����dNfv7�9�� �pT����Pr��(B��Rى�g��&�l�vƬ<	���V �e��ɚ��D�bn1�ɐ	�jAk�t���;�����{�,cK�-����/��i;m�Zo�T�g��-*������r�t�/�����MZf�dK��"�ZV�d,���F�L����P�t~)����^�i�b���i�?g��oeiٞ�{�rIR10��HF�Qd"Q�L�F0�\� �p�?w�X�����4e���HJZ��R��2�r�6\"��pT 3(1��d�Gˑ���� �Fd��������<�O�(�1:���|*볏S���W9�%jWQ�M����/̈́���`�_>$�Ii�������n��-�Tl}iC%�.�wB/=�
�_�}��d̼ �6��wj��$�_G4�Ld	�a���бI'?�CRƷ�\ׅ��3���\ �UrF���UM�j�a `+j��ykD������:\ݨu(��h}WoJ�F@����̡W��-�d�\�ǿʂ�ĒU��'��]�)7Tͼk�ϘZ ��a���=~1Ul� �|��'�S�Ѿ3���?���
k����G�k���.���5�B�&��(4��F<�T0(=���%1�G���>"s�f���j&T�:q��@n@H�h����?��D���Q��ֿ�Z�D��YĀ��b���@1�Xy2�Ə� CQ��]T�Zn.���{����ݪ;c���^~�3��[Aid��:Ml�+&�t��GrUf������^Y*�=V�9�R%��k:�ЗD�!y��;t��Wƻ64jl�O�y7F�4,^�����F���d�>��7	�j��AD�%Y@=��lU���~��<j�oW}.9�f]�?w�����X# IŐj�TG@�\x$�⼤�G��c���=U��<��+U�⃭q?���cS�%;�U��iHM���X�b��~���uWh�-��#_)࠻V:��>�4]�t�Ã>��B8�d�*�����Z�Y���j�Y�ln(++�K��~���o��y<�Xz6�uJW�wDB�A6��A�L���'�a�.�t��H���Lx2ޒ����`��EMp��
v�]����T�o��������ބ�R�]�������R�S6/�;�{����:��R��O���,N8t����o��E�����Ĥϲț��O�Z}����
e�Z�B
�2i	-��ն�flP9x��e��$:�8�ʳ/!��3�/�KE�-a(�Mo��0��)K2��l}ւ�D�D�x� ���>8l���V��_�)���Rq���������T"��, PKq�G��
p9;_�<�{R��2N$�E�3�!L��6���U������#0�Ɣ��	U�ϕ9;8��=�V�|/��'SU���"?��'k�A��g�}�GZ�bN3wm�i��{�bI6.*�Czؙϥ������.c�t��J�~���+�ׇ�F�o������{f��Զ3�9�?�����Þ���*-�r��p��� ���P��԰�L�����~�b$lq�
vK_<�u܉8c;��k����5��rЫ��:�G�ȣ%��: �Po�) y���oӽM���n�0R^��'f�� �ͽc����g�������n�9�C���g��Hl�P��{�:��۷ �M9wG������t���;�WBdE���ߍ����I���1���f��!,�S	{�Ap,�_Y����.��3%�����p�S{�B-n!f����>�3���Թ9�##G}��×�f��Xw��m��ؤ�*�u�ѣ`�����^�2�6_5��wh�N�w���OW�A�\ô��{b��N5��c���i�9��d�1������Ɛ�4դmXV�-D;�P�!��\�>�����I!��Ɉ�%�]9�����+1`@8k8x%������'C��ȿBq��O|� c8� �a<lFj�Ά����%[s��co:�$�VcsҌ�9�j_f��V�.��#�L�sE 6Y3Gwb�ĥ�o$��*�tA����x
�p�H�;hV |��_Q�3B?��G����6t�H��	�4�J{�n�G�V�.�,��������7�k(��AhU��@��;$0N�)�6��7�(�p5E�6Qn��#뀉��X��R^����+���A����{�>f� ���d�M:4a��M�y��f�ł�Ύ7�?���V�e�r |��K���l�;ۡIGRJ����C�GޅTM���
��~����"���4��ȉפ���m�3���=���On&Y��1�]��TDS�����<8��I8Tj�2*��c��"^���ԏ�(1�� �#�7��5O�͆� ����֋C-�9C�6,\.�E�����l���
M4J�(xc�9M-^-g���q���3���m0ԝ��y� �x2� ����>5�\j3�O�C�r�_�<3!�F����w\M���n�NE%��ޓ��!L#�m]'t�����u�AaZB�dvX
��#�d+��Q����˗��%�X�Yc6�������U�6$�����AD���U���2�����#����o>�~ �"A�ڝ�)M���~�*kUh��P` �7	\��d������`��2�-�؜�N�a{�9&'�O���-O��8�xΥ0^���C�lK�����O�	]·�d� Ϡ�S8Dh��?��7�� �9*�\�R����i�w;�R9m.&>u\�� ey'K�����Qf6�9����A�l钲P0�l>�;J��-;���>�T��ȃ �+g���nBǥ�a�my�F�_�_5���pk|�ȘO���iOs{?�grmdpG��'�.��pB_�C#�8g��
�D[-��٪Q���&�<�ᇂU/#�7�y�u0�����qyf�>�!:[���,[�([��A�BF�$_Mײ��gq���q�����zlJX�"��O��f����R�MowQ�� ��_G/ؒ5�c�Bl��eo^~8��o�}�.<�W �~��j�y����24,�=�C�)�¾���l�}��,�a����	�vV�ޔ���B�f𥭴Y���5t�#2j����m��3�TJ#Ko�m"(Omc	� X�<
����U_���<��5ŏ��m�= $˺�?#�ռC�hQ��h-*�6�J�`5�D�f�~N���{{��`en�q5}?��\��qm�q��h2����ʕ&��N������{���t�,�4	îx(<�.�	����՜͜�k�	8�R%Ο5�a�9�_��Ɓ����±��!Iw��)ٛ6��{Ȯ��F��b��:�j���D�
��}̛=��?�����,�[�r��neٌ���4����:P�ݒ��D���;��o���5#[ʨwuȽ���CCQ�q?b8�V3г����R��0|H���6z�|�̼�8��.��^J���C[�J� jب��p�A��8�`�d���=�埈�����|ؿF��om�"��@Ԫ�q���P��K�0�4��)��ȃ'Y<���TQي���ٵ���V�y� 0
�9
��;XRXEi5�.l�).�O_��Z�	��m.�����n���TzC5͐n9GP&�E�Y�ug��!z ��H�D���Xpo���k?iD�S������vO�x4��>���,��:���B&#h�H񄩯���ʃ��Uo��a�aY�������t[��p������)s����A*���*���_�f8��G��q�V�! �%��
p�t�%q�[V�1���d�Dm���)iF Ze�8���a�6Ѳ�oJH�� CHA��'�58C�+CBC���9�U\�FX���}Ц�%V��O��	���ǣ��%s�#jC\*P�/5��BƟH���Q-���
��gw7_��y���=JH�q��A��1��GƊ�@��WR<>_�ٕ��g]��=�zT�X\߂^�-�kL�n�؎OQ��K2�7XW�)b(uQ	{$��Z+O���<y/]��#��o$���s�t�3�0PHX�U"���R��M�^U'�����Y�N�x�Mw1d�!��;�?�#�چ��!��ezW� U}:�C3�?��`<�[/��A���m� ��1ye�>v��r��r��my�O��K���M�
�KbH��
f�u���飭����\�T�D��D��.S"l��Z�]d;�������\N�[B�gbyH��a����sb��5���	C�1GJC2���DrQ����o�W�,`x���
Xq����c�� �6��F��\R�&��ՓԻ��gsj�	rfZr�E�Nҵ-@�6˴-fI,1�"k�{E/��Be����OJi�na��d"�
+j@�r�$K6Q��]Gˑ�w8�������c�Џ�(�������bY�F� 
j�'���k�kEp�m��[�ED�ٓۅ߹m�"HZcR4|�7�e�����[Y�*��DY���$@����F�b�3А؆��?�5���P��^(bn}I��;�`�GB����qW��E]��p�:�a�׺�[&�M$��`�=�=� sF�b��YACO`oS5�Y��?����_]��ǔ+��ѽf�i� ��Z��C�8{����E&xy�|a��K����P��yD� �Zl��St��u��M��4�UN�*c�?���]ʔ�FZn�ào�,�9�Ǫ�?�g��-�k4�ɠhb?ƛ�˅P�������}�{,,p��=� ����v�� ��a��Ϗ�n=J<cճ���/�>^���r�@�[��V�ѤmϷc3ʬ^�є6��m�����TX�%'d�y�a�� �Uc����\�$캺�+�=��@��y���uv�����8����z���K"�,(��V%]��n�p��UĊDvf��+������7��:���H�ʌ��F~J���^�5\:7X�@;����ݶ�b��<�qJ�68:9�J\���Gw��.e��pΰee ���D�|�%>zg�l��l�� �kv�'=!�L�HG���j�cC�-Y�12X��7l�3�5R/;�+��-��ݭ��&Y���q����g!�<
���������|�il�ƣ��Yv=��֮��V{�9�!�"�\nI����s��]?i���]�\���R�r�tj]}cafe}��:�"J�t\�xXc?r1r:�愠���xr0�N�)b�cvm�R�)D��!���E�dj�폙�𨆄����ʖ��:^XX�]ǰy���vh��V����Բ}�B��X��q�8��v�����������jE� ����Cq>�X`/�a����2B$�&��"�v {=F��םk����	�k���J
�?<���p���uCN��-��uL�Aᨓ����2�&�q�ȭ_⯯��&,u��(~��#=��[�:1�}K�]b!��^�\���7?2�d_��I��}3,�@��a��=�L2�D�V���^���@��+�-+��;`�Z��n-���tg�m,���9��hU�?7�bz�+�
�-wO2Vf��%�����v~y��O+S�$��)of�4�R��QLd*x����^w����K?7�D���9����)�B�?SP�9��a�1�*�K��	��֧>T66ٲʘ�_X���J��(�M�"��m�L�fw�O��#��(T`@T�*���CoLҦ����
���kZ���j� b��<g�9Ԃ�k�ys,$��[��I/䲋�B�6�� ̚�d��fp����
ɽ-�S5)�P�	۩��I~��<���n�� ��l3�B�8/�8�V§r��\�:F,�m ������o��$lv��]�c1�Q�ko�6���3f�Q_aP�>�P7�]����J`����5+�*ߥ�7��Ҵ��r���_�r���tˀ0��a��Ul�0t�ۃj�}&��bSpr�D��쑆]9=��}��#���-�6�0�xl�6�_��k�����2kf��J���nh���Ŀ<��i:)��h0��Ŝ��V�\�|����/6�*p��`�V3�]��2�� �:�k �|s�ʷ7v{
��|:f�=L ׾�Z?�1I ��������tb�ͼu
S!����F0_8i|*ِ	�D1ni���zW�]~2j���lH��U^\��q�
𳍹0�9�ۍF�e)?M�O�v��(a�gX����۵W;���Z��(!� B����rCO-�B_�"�Q�j�Q�c�s�ߴ�\����v���ge�d}'��-��j��!=�5
�T�M@H���:�C �Du/E2�l��"4D�^�+)���~<�����0��*Kټ����Ե�����^�h 2�댦�w��f2���孀����o����dr�}:\[
k�����"]Z�Q##r|�	�������;H3]�A��%�R�T��]��e\��n�!	F(.h`�����{h�(G�ޤ�")��s{-�w5��e+:f<��ӕl�Rٿ��\��G{���3W�����޲(� �O�8�a�-�G���SFD)$�v ���2b��Лt��,}�����_�?̜p&��CZ�j@'��o5.�p�Y��S$ߚ�	�;n�����uY.�N,�b�N��o�zˋ��w�R;��9��-~�b^�S�á7 5�.'�S������{0�ǁ��k����"^0�aֶ�Q��t��
�_��ɯA�ȸ��Q�%�^
EY��l�7��x>�L�l��EO	�P�ÕE{�`�dq�s|��0����F�¥�ek��'�m��F<yl}*�o�Ș���޺Q� ��kgO���9])������K��c��+1����\ҭQ�����S�s�q<ԿA������ݿדpF��͎���� ˪*������p��)K�էp^��,s�-Q���wE	��q��(32�?jR�5��� ����"5]Z�cc9B%���i���`�5�!�|������*�c���w�n�:1�Jϣ���]���[Ƕ�9%n}?)_^�Րo��iGP0�9f�_+�hD	�S(BG|�Y�� u���:|��`�47��S� ��?3�*I�S�ֶ�
�6F�9qvn9�0����.�u�HQ�͚;!�.�pt��4n� i�2�7�I5�;��l@?I���u"x�h:��NZ� �A���tj�}lD	�ܔ�jKk�L��{֊��}��LZ�y�t]|�Q%���>�o��K���'ք�3���>]b�ֆ��?q*��f�p$��;�2� ����;�X�$v�㆓���N���?�n~5����܄�C4�wac�ؐ�V�w��w-Ŕ�`���PD�)��C_����Bχ�L���pc��2!0����l��	�vW�w�l7bѨb�����4p�����X�rBp,0�}hG@-�Pl��FhO%n&�vt9�־�����G~p����d�0T�o4,�0j۳zO�����f�ƛ��_���-��28�/cDڲ׳�v��Fsa��.�R�+�Vd�.vJ7��cI@X��������Z-a�[�����˹�����I'�V��Љ,��W7�4��b�m�^�m�T���aݭ�8*��u���l�a]&��@���?M�Y��?�R����gVt�<�j�aX�
7|��[�q���S��EqH���-�����`"'M~5�AN�L��fc��Q���q�%x�-����r�fIқ��Μ���ۄ�ƉN�f�J�9�-c��<�`�- �-�!�߱��T$�)<p��O���>Mi���Qw�=v��Q��J�ʁ�e�!�9��(�����ɰ�2u�C֥"m$L47���݉_���"ւJ��{f�� �?��:8OK���S���#
��М���U�.��痐_������r)�:�x��4�u���Nl��$�ѧמJ��duXx�j{$�Ά�]��-�s�q�h��$��5E��G���=�V�^�RW������,���9�,*����b�s^�<�h�l�J4a�)a������E��u�0���*���ᐼ��͚����I��1��+�8���}��)�ఽ~Cߊ,,~���])�%�{)�����)�Y�d��)��1_P���J�?�-��)��xJ�Ǚ4��E�1�,�Ӛ�t��C~�#�	�q�EvBK�#ѿV�����]���\��xxܣ��ׯ˰=��Í{b�㡇�~}�0�[��֯xn��b��J����ϧ!�˒q;?�K�Q����`���Tj�b�hh��m�$k�E�� �<:f�7��e'PR���*ò��E{�Tj]�x�%���j�4��%��cp$-pw�,$����9[�r����B4O.��LϦ3~��j��+��P��4��I2v�t���V?�9L��׃��3��a'� �"#����ǐ�@S���U��O��*�VU&8E �1S��@�#VԢn�hg�B�k���2L�T���᝻E%�h�"ju\��"�z�]����\�=)!���]|ך���K*�n��X	��V�,2�)
7m�|������l����Q�*6J�jI�}5�Ⱥ���>b&:K`(x�ԎN��[�j���_��H'����,4�����TX������Z�mȃB9�~��>��nN2��4�_��?VQ���h����-X�n_�c����\���1���=l^"$�Um��l��<��L�O��{E��VA����(̛5R�y�f|��#��o�ϨCd ��7Z��B�Z߂�*4��#���a{��ш�Y�\�ϻ��dJa"�w�u+rJ�%�g��s'��3�5�i�}�>�����!81o�=�����"�!���5:,�=��p����L%?��%,��AޭZ�r���n;#��qf�C*�L+>C�oU��
�m�%%ތ�S�ldTr�� m���%���S4E���@����^����M��᳾f�`��*�h���r��/���.�צPY��F*��k�O�\3�[U��N2����)�`�7T�|��91=h�1
K�r����6%��q=P�Ҟ #��c����`<f|x3���V���GQ5��$;���O�6�+l�@��p��>cqi����e�B�3U|��q�/���3.�n��r�\��h�Q�QU0k��;_D~�KJr���ͷ�7�<�F�RYK��()��O~����L���7�ٵ�����)�v1��j��{�`P*5>6� �ߠ9�p$I:�V&���\}.P�ncGvG��s��f�-�bb��,Y�
�[h� ����ԋ��t�m�5��;��yJs�T��O�=���9�tPO��{H�B�(���79H��9��VY�Dg\/��g�}H�d�ӓ��f�Sfr֞����J�흏��)�ː��q�[���n0D����L���4�N�l���<�ν;���~�'���/\��I��a<�p��>%e�����h��	P��_�5�	<��Y�n��Z�׎� G�9KLڤ�>D"q^?�.�]E$�\!�0Kcv,D|�Z?&E�ujO�u���~�`�+���==�-���#"�f�tq�&��h��]
�"��6��z��I�#n�$��@iɚr@���6��e)��'���
�aA�	��y/�I�7��wZ E���;�/�p�F�שA�N�u�Y���;���<�oX�)N3�Þڠ}�f��Jsy�۲s5
q�yhO Gߑm#v���f�*B�SP"*���&�6 K� �`@$���v-�%�b,eW҆΂��J����k�����B]��~~�w�h�`4[�4�Kѩ֧дe�!�K���8��\p�N�ەU�X�D��������t������;��ʵv�����{;�p���Ѿ��+r|a+�O��ަR��J+�D��jo�.:)���Z~:Q����BJb1P�ø��>7W��g�2/�^Db0�D�\|3��&pXc<u�z�f�����p���a��:���!�4�ʺ0��WiȖ53׏�_;ύ἞� o�Y���
@iO��(V��jKJ$��jˢw�{�Z�(o[j ����:�e
ۙ"�rYJ����v9�6`N������;3��o��>g���%`Q ����J��uM;̭E����&����b�6�~�g<��^!����.����-p��!{I��o%ߜ_���G��<�	�6��~�m�RL���N2�݇�%g����j0�c�K�N�O
�^�I��|�&�3���ɰ�!_k����Lb<�ȪD���7�wULُp0��(3-�����+b����3��.�������=��5U���r�F������]��0���ȍ]�:fUƁW*�0�u`��XY[ɺu%D70^�*2yt�ZF
a���W6s$9��l�A��%�F*�]ܵ��ʎ�ݰ��I��ϗ���1a��FT����Fhտ�+�P��"���g��n�� ����YI�{��1dV�OvW��K��Lݕ�?�_��/����ЩL��
\<�Tq�E���v�G�s!�������[&��B�X�Y��