��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ������
D�5��L�k��Cؿ�vͫ������i0�k��c�1TX�� z�<� F�I@��q�
���O'�?6��Ue.R��3�պ�6�d$mx?3.����{�^�7/~O~N��Q���5�V}��A9M����j)�R5���=���=W�� �7��-4�d}�3�M$x��nM��%��2/��p�)ꋅ�>�ܹ��yxn�w���d{zE#�m�ɰ�W�32��:	lP�F�p�VQ� �#']�
�mnW�/ݻ���T�/ ���䌀��L^�lW�4SR�m�l���utDmvi<J��+����+>�5����s���ro����\7��L k�G0mb�U�5϶��QSr:ܰ8#�zƝ�ͦj:h,6�n�B>�!�^Z�gf_���=�f�!�X�HL���u�@LX]?��1�������0HC�����������%���P���>;b<���ې�<U�^��!j���,Ԧ��I,�Z�2kl�V�O��ͬ�	��!sL�4��Sa7�;� sj��C3}�Yc�_S۬j��/�iZ�܍+�_
R�苤�N���H��]��~�r${�o��4_&?�{�}�w��cff4I�AH0�=���b���%#�&��	��"ؚ�=��OL�ЦXi'�C
��H��{���ω,�b�A8����r�K�b3�+'o��O�"_v^���7S����K��R4ks��}���q��W؂)�?��榮�Ah%�^�}���H?�2��/�s Mt�_B�-��N�י��G����}�wa�kӵ��)#���9�${��E��n`8����t8+��74矮MQ���ƻ��%Г�'lhu�C����o�1����r��8��wr4	c�
odr�(�3ڷ��w�'<���;��@��mI"NxAZ�b��v?�'��!q��&��َo�Z����G�����x��½v�q��%"�>/|޲.r�r^ᓜ�濺tL��~x3+�5�v�Po�_������t5�����?Qx��3�k:���`���)�GE@�OJK��B��W�]#�`�^YÔ�K���4��xa��M(з�to���a��L��-����^�+Jt��8m4L� $��I�1�[��m��k�D1ֵ�N�WŶ�zc�ء�1�.�����2J2d�*�7HY�Ƽ��F���>���VG!�� %MAV��+��Ŀ~؉4`uH���:ǲ�¾Ix�+�� )���������kT/�:�/��TT�Â6)���m���:#��nZ���{���~S�^���|'~�m�]��T�����G흣!j33
�.a���1�Alr���'��k7�	�/�h��
@�.��%��
RJK?�����o(��ή�S!�$z�}�	��G���h{��$?�����ԤsUO����z��т���sv;��Ĉ0�����QU���]v�W�Lb|��PU:C�8ಥ���(�	�k�GwE1�]`�RSp�)�"4;Q"�dֈ�{�&ƭCFe*���8%#ܯ�];C5�8,xQ�����]G[�r���{f ��J\<��v����e|��S6�)7iK��{�jR�y��_%��r�f�6�J��`�.]�GT�:j(l����Y(��m�J��8@-t����/���	��eߠ3Ә@�E`a������$V�	��j�#�t$�]39H����_�C�razG��+oJ)���5Y8���7��)���,�oH��5Xaڸ${S0Wh],T�[���dE/<,rLn����+�)[�ӝߌ���̷1��g�Y��i�qy�Vw�8�l��3���S|e�o�Q�P��AdV����+s�
�<�tZ�3.�� N���7L�[qX:r(5o�IL�`�Aj��6Hw���h
��PT5���n[�sDN�PP����nb�A8	խ&����W�dYRN��W����v��R٨�G4p3~yϴ4^�+z��`����[ڹl�|����t��bkgw�A+��=E��\K��*�y�q7
z�eNC�41���aj�*��2?����`��0���h�,�U۱�e�L�~~��P\,�.�QH�8���$2s��Kl�a9�.�J��w���7��~��_m�v�}R=B	�ʦZ��e�,Rô
G�.�N����"���%�.��p�=e�^�zCN���a�5��%A�e#8���C)��8�ێ��?��~v���6���Z�tlA��W�O����C/H���dV�! Ew>0.��Vz G\��2��z�\��܎z$H>����hf"�%�،������V"���HpV}s����Z�U;��<Me�m� ʦ��%�e�]&�j�BL�+9�W���9�\��~8�F��oR��0����\1$��En*�m�6Z\S���F�:[>��#P���rN���)��|�pʎ�&�^�V�%�W`����]���IB�����F���Ұ�q{�@���F�m�Ph�F͍����c��/�N� �O4��O�97�qJ?���*��TG������&g83hXf�<撗�ׇv6��^�_�Ĵ�������5佚ڜ��$8n�f�mg��M�#�K�b���N � YoĴ��c��q����Qm�Ҙ�e&�DS�V�����z���%r�������#\�}��ރ�`�R1C.�H��L��d��4�AFزP����iAoQY�)�])���Z���[ب)k:��j�f��r������D�{c�84�
$8)�=ĽUV�"Fy��Ů��p��������gJ8�&i�> �Q�f�J/T7`��w��
��E
g�P9¡4v2�Q&G�?��_w56�W+ ��g��Ԅ��f��XTl�zH ��e�7a��"A�,�x ��n���&5g�S�#2�<�'%t�K�OUL�tv?�
cal5��0,��Y^���rge�R�C	���6~ޯuy�}�����*���Y�wcI٠ P�S��i�"=B����!)V�n^>�
�F��v�AL�:	���R��X!�T��#��{摫ċ�u������iq��@���kP%��b�J*�*~���sݎi��C(O��!��s�v�v�+x{""��Nw׵��I������@t ���>�Q��i������rF��r8�_���/s��*�.Y]��I�/�A������
R�m>�J�֨��/q2�h;�\��Y��:�R��_�s銹�*ii
�0/��Zw�Q��?�a!���sKt�*�-1-�앥wE@��wJ7����˃#˛�h�5�����!�G%3' ,j��Q�/f��T}.?�\��ӡ��62��\�<F]��y����t�췗��q$��UϹ�j��V�m��riկ��9��Y���1�flǝ݋�`T��&Z~:��6���7u	I���p~q�g�L�嶧�Y4E���`��[��HA�6٨/$�c���g��85�;�/.�7�3��l��\m�$z$;�t�D���b���F4��W�]���0��Z���i���8� L�Vd�����@�,�&�M�?J>F��UT�֞{>���H�K:�VMH���g�ۜ�dA`X�3Ù�T��}�+b��=p
���㢓~G&"i�����8���v��}�+T�1�u-���g����\�!��/��'d�pF���!z�5���v�zК�����F�Gz��$⥽~m)�p��Z����/�n=JnNk^g���9��2������ ���bǷ��>\,$�7�y&n&2��w�����j���@_vǫ���-��(
���M"�Av+�fsɋ�����6�wd� ��1���T��~vV�=���e�2g�LA&ԇu�4Υ��֭�,,�[��"���w�F�x�ڗ��%�j��"g�������xn�u�G��������bORP7�n�WCG��M�z�Z�Z)/d"x\=<g��j��J��s�Lh�a0�l٬���n�����km�q��3�# ���Y�.%�K����O�d�LB�>6�n��g�W�C��p_}�gr؟�#Eۧ�Y���-\TV^Ż9qB&Oj���䡝p3��m��4;-�#Ե�T��(�J�A���a���̢����x�L��|����<��G@E��q�t�����v�<�a�ijI������H&�Ѧ=�>!�*��2�m�ĵGn�ǐU��ҞV����=o�/NL�)�]?e�w��׫E�9a��\�j]��bfv�%R6g$�h�[��L�Ի�ؗy����y���P�ÿY�<��7'�O��><Kt�Q(�mT��|F%��������Z�g�ם���1��(���4��h��ҩ�D��	4O+�x��vsje|����f s��g�	 ��q)�[V|��$�i&q��!����nQ�՘���F�avo�m7�柤I��֦��j]�kܾ,�����2i��;�~����j�� �I�h)�v�}�i��~BՈ�G�+�������Dm��q�l��;w�WVoZP/�U��_[�L-kE	QrҺȗ	z��󮨻�k#�6|'�f�:>�C���:5�@��R�@zk��ߖ�B�E�hI+��y��7Ұ�
�9�,�����톢j�<�l�Jx�����Ǖs��s%E���`�9�̼g|��r|�H�U�lt����-�]ɲw��rg�46{-N��QxL"��t=���M&����R�B���ӯ�p�
��d[�����^�;�K����W�95������SvmO�{�Fv��ˮ��v>a�֮*b�p�u��RZx�LC!����C�t@3+�J$v��Q#̘D�`��4l�,�*v����YLj?��T �f5�]��]{=�n�gI�J�P�[O��r۶�v�fɱ���)F�:�E d�~���Q(���C��.W��u1*�XU���h(:��H<�:���`���N{<��x�.�K�c����w�&2u����,S=`��[��M���������fy������"}�����DU@,����on���W� ��n4i��r	d}v�~�x�M�����g�ycZ��qHK"�mA�Έ���L�J��}>�
�RJґ��M��o�cY��P0��\~��A�e���r�ގ`����z,�s&��d<�I���L��Zr��6��f�]�����i
ݜm+7�\�)?��OU�6`�:�4�j�"��CHƅ��g;�X��N��qB�fb�Z1���1�	���GK$���GF��:�3'�}�k�_qg�F>x�n��M˗�쩎�؇GS2I���(� �J�����+0^�s���^z����}�z o����ߵ�]�q�Y�4g�;) ��r��q�D��p���6�J_i,tF(���JR�°�J3L�7:'F��u.{:Q�\Q�e]��1{u�/o��ڎi��n_���7�R�g���!0�F})�u,�e�ʀ�T!/-lYA$NL!�d��Kd㵦����EU˄������*�M���d��h�������\�>�8Dl~�0������4*2mjM�b��-�腻�h��c�"j`2��Q%KS(w=%��_�c#����5pd��͑���St�"��s�d�ّ?`�[j�)у��#A7��9�ԮT�g@a��V��y|�U�}\J%N���h�&�J�5�9�cJ3Ow�53�����NY�H�Ӭ&���{�ǘz$���%�� U� �2U�?q��lg�zSiⴝ]��ژel�633�d*9�2U1
q+�9�!J[B��/zV伕�Q���OT�ۍcD�����64 ��,�#�F�풎L���!g�L���[XR�oC��Ab%af�0�x_���Kl	 >
ϙ��'���_ ���PƗ��5�HB`��c�.���{��_7ҹ���4�@���6�o�s$�E#�l^�z��W��v�sS:P<��I���D�@)�O�0>���J����eƋO�S��'��i���q̉���3rH<<±�}ŤKZ1_�Hg���""%{EY6��}A~�z��s҇�،��<�"��
q5��rND�k���ژj�V�W�����F+��j{χF�>�T��.��T��w�F�M=��q���cq������9<W�鐓j��jyg��͘+�Pa]�|��������f�(x����4�y��~�Qpi�9�q��=���	�����xz{����Φ(���SN�V��NL/K��Xluת�z
�G�z~&��zX���ڤ���
%�V�� �XC��]�����q�5Ԍ�S�6��I��&��4�����0��x�z�������rA� $b�~f?]B
�LS{Ϡ@���my�Tʕ��x���Q8,��2J5���>�h�K��	0P�b6*��l��a�.���J�M*0"������2:��2�w����z��+�	�L���d��pibd�D#}��
��~��j.�49�g����l~�Ę�'���V����Qu�a��q��#����]�mT�^ؖ��w�m�����PDz#��.���v�Jƈ�#����g}�^�`��ƻ��7%����m?�P�m4�y-���($ƀ�" ������_���S�l�㍮��:u�,��{��)Z��b���QQ·�N"�6&q5�yDo�A��Sn���ZObGg�߹!��0�墐T��J��7h�U��(h+\��~���}͛�Evb
�ʈ���F��`�Gó�zǔF15����ýoc���?%�ϥL�?t^a�T���BȑuM�ʔ�`��2�x�͠3�h-֥ C�V~!�VTyD���N�&�����/�$!<��
^���\�����c�Q	4�Ј���ֺ�N\��D+f�s���eZG�i��4��7%6��AR��d;أ����F]}�V��ir�!7��K��K�F��]���Y$�5��ۊ}�B�m�wR)e]@�/��#�;�?� kOr#�Y�6]��ZBJY%8�	�0	�����{�3)�=��uq{�f��:� =I���&�OK�_��v4w|����Չ9�q!ʖ|&���V���y;�ν4h`Y�ay|v3��Up�]R��˗Ii����f��"���b"4�A'2�'���׬f(�C�C>I?g�>��f��f4��c�n[�Ux�2�7W|<��1X�I����RPb�wi�taR�_�hk9����X�4�����WJȬ���y�l�bLp��6��tF�3�J^�n6�!�k��3�-�v;����̻)~�j�)pˆ`U>z�'_�f����1*0*��d���i1`�݇�bn��l@ː�HZyDmZ�G���q"�����F鵢+��9Q��N_N��
_�˿@/{(�!�Ԅ�~�l�ِ�����^���?mExYT���P�)�±�eOy+ŝ���I���\A����� C��`���t�:r� ��C�!�1��b��IVpzy7<�8X�L�j�4��-�RR��+�&�O}=a5׌����lR��Į��q��͌恍�ҭߦr�H�nE/�%��,e��l0�11W��-�v�+�ϧ�G�S?�&?�����]���SQY<%�ew��"F�����Uq~)�����qa<���̽�b(�B�u�������k^�����6Y�uW�
�����Ot��ltEe^x��
'������ZUGP�U��^� �ʿɏ,)eRf�F���rs�N�-Ff��} p�;F[DANxӅ������G��5�^!��o�|`�lS�ǭʄI��!i�O��������P�wPr�q7frLNn�P`��A�Q��H\����%�MF閼^�b�ڣ1Tl�yį$��P��K�A��0%��`e�[�-D�X�����\y�hW&~M���@��Ϋ���TO���E(��:�{������h���s�*�L���L�ȏ�2Y�Ѹ�5�2�(��9j�|p�! %>hc���S����g	l�W�bǲUZ�c1��]���J���+-A�|��D�y����.���&������~�r�5��J����
g��0�_X�E�|QL{H��&*z�	�R)\j�P�j�����k��|�~i����ڜ j=����A�;���2��#�;p�^�,��<(�M'#�uY��֋��;ߏڡr�63�S�z�� {���q�[oDS��b
XK�>�����0ͳ�W���jC֙�
����6����k��3m�Y��&��{j�(|���D3SE0�n�+��3gK4�^+�c�b9z��{��1��+D�%���~!�[7�~#?�픧��	%��=��+���!o<��͇���>�>�4J�[�Ơo�㥑��������P�Lo�]a����@��|�ؤ�Z�I�����J$)��Y��ڠ���`� ��~ڀ�mʷuɰ����oU���T�kx���Zb�x5�q�xgh4?�&�1�8o����p��OD�[�@�e�bƦ�N�0�,bʅ��DS.@����d�ui��&;�lX����s���wF{T���F�[�}J��R��@ܲ�~�Y�z�d2^����� �Ǔ7�?1���B���s�w�w #�+x��s�Щ� ��ѣ��9����Wϝx���[��db6�G�VU�z�۟?���'u��2�q�#+cL�4t��t]�Un����e�����:�#�~_[��}%�=
p��w�Q�O�V��L?@����VD��.89��9��@�#�!t/�<��h�\���^dp).mh�l���gT8b�X�Tw(��=e�xd�:Q�٪[s�jj�Y;���%ȱ��'�8T(��<����_8qSe���@|
`�_�NNgwѧ����v:p��{��s�����װ)#9�M����n�Y���gN\4D��7�(�2���Ɯ�g����k6~��>ԗ:X[
���lXs�#S	�"
ų�V�K�W����W6Sl��1:�B|���ԛa:��_��������//Vr�KЙېgFqU=�=�(O�)���w8�F$���ãGȪ����Z���b;�%!~�!Z�.���UK��`�������Yv��S1�����HGC��h�B1_c�gӽ��%x�T{�f����XḊ������`/���!����a�Z��7Q�ø�e��C��%M,�'��b|���,~�mL�e������KB%ukQ]�bAZ�Q�'�I/��iD	Y+%����;��`F�l� S���#]�=��m��+Jn��=��c$k�ke�k�m�+�8 M�L����[�i��=��C!Ax��nm��+֡��\C�
+V	�JBS==��t�al���ٴ'���,��>f�c)MÓ�d��hNX�ɯ[�/���Ff׿���e@���)
b���|x\u�Q�����5j�QI��|�{i��x:=u_�Q�T�^vlNtN���f���%�������xI��:�3��$��g�4�Ц=\����x�+"|��"��-ձ�JC`�J�]ɹ{T o&*ʍ��;x��D$7c���������\�DA�A�$�n헿�E�{x?�[�}TgC�Aؚ�uSD|,4�C���`c�+�����!z�0�;�-�$�"���fI�f_��n^D�Ӹ�3k��$iM���A�b������cVT;�:~��_wS ��|�"�e�{n���22*G��tBy���ߌ�SLy��J�	������w��p�
�¥�k&�`%P��LO���?��{�ts�[� �oL��R�8Z�pYl�B�xD+d�id�4��
�4����݉?yB�bӰs������~Q5[I׻��(<���W65`�tcF�"��ÉO�#�N_�^U���h���wS���h�Az����*EۼT�| ��q%�����d��Z���iJu{9�f"L�Ej�ٷi��<t�X��ŏ�&�6
6�.ȅ�a*�؍G-���rw#P��K�v�d�"-{�7������k��HlM�ׂ�u�:�gCJE4l=���"�Wg�cG��&�� ��X�VA�e�E���� D