��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���N��`�G��^ ���F$�(8��<M4dG/q���j�(��VP��G�,O�}��è�
u�1�ê��Y&�"}:$���`����INmҌ{ڊ�|��M�v�S9�~�H�����E�'�!��	wv �.nя�J��urCP<�1�D�_���ҠHP�tS3��$6�sq���}������ތ_�
p*������3y����L֭8���ESE
��[�����].�.�NgҘ.0��O�
��@ ךj��lG�&�%�U����Bt����I���Y����J�8_�Ն�`[�h� kgmTJ�Ah��-;�ƽ�D�"hC]N��nQ�[HA��i��u
��g���J-Ҡ�,��6js��K� �B��}mqn�<�+'����3ƒ%+z-K��
D��l��K�D��fz:i��U�ޅd�'��_�TPO��h�PO����>���s��`y������I�F�Ա��u�dP2E�岬.w������BB�e7`fe�ځ���ÑHYKړ�ח�nv� �3�6ګ���-�	Hjna���RE��1V1{�8{�qt@q=D~/�Rv�M�� G��ŉ͈��b�b/�Z��~����Ko'Lߟz��h�2���#+��+�B~�!?D�`J<��j�(Y�#+P.�mۉu!$U��#� ��q�J�ڵ  Œq�l�r���<�����/�ӀG��L-7#dZ ��6h!;N���s��G�tq���I��Z���tU��n�ajf�!Yu��۳T �Ͱ��f9�����\|�v�>p1�'����m���q*�M���N�[=�o;����xˣ��C��;,O��ۯ�
z�Xop�p�ER
+��Zx�$�#s�'��X�w\�K�I�(ה��s�w���� �������*yt��4E��zZ��w�\*�\�lGt[�KO�g��;�;����p������yФw��{������F�����.A<��ŒPW[4��Dd���T��;�a��8�||�� �S�0�P���Z�؝9��n23��bڰ�o�&"E�q湍��Y`���ϴ���n�1���-�0��9�I��l��	���<���������$q��Jw�<X��Kb�N 	�����|M7�Y�0u��F���G�_/pe���(�'�l�K�s�Ũ�k
�?:ézTL%��?״�����F5�e�>ϒ��ۼ�"f�:�/_f�w���@9A��!@T��r�"���ޗ.2�F^��3�Eꩶ����c��uޏ
�6�ۉ�>��TIE:�kx�[�o7���P����w���s'���*��>'��{�Vr�au��H��{uP�zk��;#�>>�XC�H^��*�h&a��D˓��?Ws]B��%���3W���x����r������af&{+�35L�<=��k��mrU��ο ��d8BY&n�	�3�m�6,�5�ډ���@�Eޠ'��Yo��}��a�;_����?ul�"hUem��I!C�G��&R/K���V�ێ�<��Y��V�h�6TvyLj�
�U;�h�(���4 gf��&��`��@���)�5�}��l^B���+�D �זv��G���o�Z������Bs���r�~e����e<��j`�ۥ���;I�TX�ü[d�p�$�t��7��7�*�2�}��Ύi��}����}ւV9�mH�����f�o���"d�l����/9��en����1V���[Si{�(�rw`��DP ��ujh�����F�?M���NZy�Ԥ�F�w�ܞI��<-����y�0���k8���O���[e�pÔr'|� y�R����9�\�<K7tک��u���8�t�)uZ=i���A�������)�v��yo�h��$?7Ԕq�e��*�1�ٽ�|���7�^5S��6Ϡ�G�5��OF]�n�T-��m�kX�U,�y���M�]}k�}����8)�������g���#`[�٧1�X+3��������&	:(0���zV��4+j�"D����9�l�d�V�&K;��)��{yNu��]U�Ӟ�w;��Y��%6�ˣ �F�_+�m-Ō7�0"��aB�
"?��	�|���Ow��1���/L��:�4�$�]�|b���*uA�0\̱ۥ�nkTM�i���<'�C�E&kPg��(�7JšԊ8�.9�3���Ev�FХ��4k�49��:A�ks	��H1~�IYJ��	g�*�}����!�{T���bX'��ò��M�V�J^��`�c8`���J�M�e�
��[�61��WQ�!QMp|��-"�]�	: L`Ǣ�x�mv澱���e�v*_]�ȣ+�c�8��t�׳�ɠ
����AEaN>~�M��Iyj�Ԫ��8�kc�9`x �2������HQ��0�`��}���fm�KO��������+�AJ��zWc%�+fNַ;�xbe�hz3a�9.�8.!�U��
���1M$���2<a��)pT��"��"��r�0A��.�Y�E�)8a)�E;�Y�`�#y�3]ˠz fd]��<X���?]i=�h����l�,�)T���.Ჶ��`kr�oh�d�Ww�dwa�JwߧhP�)��.�����=�i��ռi��Ձ��t�/��[fЛ��1h����ff��Ѽ�������Y3$_��3�`���<)��m�DwJ�#é{�q�B�Š�-?��mBM�c�o�C�����6� �d��̣�AzG7���}�\MPV)@��=��s����b
8g�v@�>����P��hB���o�hi�nX�V�f&�]��]ܬP���$P����������V+.��{�4�妡�3)�"����$��tbL����y4z�k&�����+��i�5��໅@�v�n�|? �1?�J��V���~*��A؉�t�S����JU��/��!?+�����j�zj�Ͽ�g}$�PJ^f��ja�$[� :av�����j�An�H���s�yd�!�N��r����a�iq�u�"	��}�f&��;	�������ul��aH�u]�D�{N��^��?�1N-�({�cH����l����, ��5ъ�	R�����&o�ˎBˮ�t�~�����^ӯG�c��{�!I���(Hy�쩄�Lo%jՃ��*�_;�u�+��	oȝw�(�
Fv-˓iho^�r�`�}�4}����U��vռq� @��kl��O71q�)�n�����?�����h�:$���Agf�NC��Q�Ejܗ,�$n9��/�kh���7��קp5����d�C��Eoen7�2�������V���U���Ձ�NXlI����:��;!�A�0;��j��'�%�y�+i}��fF�U~�M�����|�t�g������Ƌ*�&p= e�7�>�v�խ\ë5�.�_��D8y��Q��qǍg�_�f���Ш�2�#��fM๣�n �4e�6��/{�s�֋*.OJyyQ�i����M}�j]
�UǗQ�q�!�ѩ�T��M��:�����u�/�g���Av�&������Lv�/v�܃�?�ޮ @�ǂ�+�b�w�\Q��M�c'AQ�/#9~�\�]_+gC��\�ؗ��K����R���;��]r4P\��N�EF�h����m�e���c.��)r٧H�HM�2>���JO��9��"�,>���B�]��[M�R�>��n���qCG�SU�\�����5�N��8K$�cWz�%��<�H�U�_�_���m$3�|)T9w�+b/e���#gyy����0I�I���i'Ǿ63��d
ר?Y��B�2��3�+���D�Q;�~�Λr.ZHN��7y`XE&����W]�s����	�~8�7;ݠ�=�p+����`�^����w��\�5�d.Q6�E����ysNt���|V��L����@�8�.���[����|��M��+0o�}90�P�A�1�/�Q3�i$�K�+��3��co� )�,���TZ84��[��Q���nX�]���y��Z֦q)v�m���p]��YU0��$����;i킿����#���o<?�l�;�z�Ѵ}D�F����`"3In� H[�qy�+��7`��!��ӆ����7>�܀v����8�fH;-�Һ�`�gchB�p�ԃ7n�-�'Fci܏��b{�}��<: D�橎�E!� Q@Ԯ���[�*�SA�b�2���ÕI L�`J�>�.��R�}¿�?��?�ｭ�����__�v���v�D#l�N���A�BǕe��{���<Jw�ÚE-pf�f���Ԛ@���u 癮�Y���yb�70=�JB���uq
UP�z�m��+���y-��p}����B��Zf����QJ��Q�#F�xJ�M��x��F�Iܺy�	�oh�Uh���\��X�P�,�h�'N�sCg>W�|f��h��"3�8}ۀ��YS���_�@��%������#6�f<d@�S�Jt���7�v�K_)y�/� 4��es��R�oOWjf�=�}2р��t���b{1�U&����C	�}�i�و�@ח��R� w�?ڰ��̡�m���;MU�6ą�x��K����c0"ͱ���ho� ,�%�
�k�D����/vc�P �좆r��\��c��;G�Sh���y�vE� �8Y��X���JҎ�'@�H9�rS<2�L�Q���	X�T��7���XѮ�!��R�*�eF���=�ܯ��suռ���I�q%z%j�E���D����E���=���7N��垪��Lb��-����:`����va�4�	씕�}a�E��r�)t�ʦTHl]]B~V�͢r5���t��k$=�@���E�K�8�P2Z����3&�_`����[�'�j�@
��R(ەNI�0�V��ߛ�-
UP���`�9��~��y!-,�g� �U����!BP�0���z�,&Z�i������(Y?Z�B���q�q�7��Ș^��]K�+$�#�Y���4��g�HX��Rb�|�3���t<��3G�����:��9�d�a�.dn���"�"��#+���;�W
�CS�y4���	����Ͼ�|�>�3-JX���E���r�4�אWN��FD´�cB2�]Ɋ'����}�n���U<� V(�(	�`��9�4�Nڧ�;�������� � ��m��?J+�L�emg��$��-��b$��:��
[���pE�}�G�f����\])(��@��.�d��j��u/��ӻ堲7�2����� �X�U�<9+��齯*�Wؖ��W̢���S���"�oȧ�����k����K}��
'�� ��2̣��v��i�`8�N����%sN�HoK�@����Y�Y�:*���À�>��~��*�0b���vE����G�OM�	sϦƪj0�W��d���.���'f�C���~��Fхv~��$J�����,�R<x����Nݢ�m�V!�=N{�V��X�a�-�nB�h�SIaI+�Hh�׳�$�Q�o������	�������)�ꎳ��U�4�"|���ӧ���Z��n��=�����a�{��<�g�8C�v���.�uş�_JB�7�M�A�����3沋�(�����;�J
�a�u��E���lXΪt�K�d�(D��'7J/CZ�^a�s���eF	?��'�!�6�eA���������&�YѫK��yz���A$\,]E����Kf[�6�{���t�"����G�B���}�ҞWYP��hZ�̼-��I��S[�l��*n���������3���%A �]s��r�'�)�CSɖ61���n�4'(o�O-��|�r�|xh�߷�n����E2�V��op�E��/ى\x~��CY�yؓq��	�v��&Ha��z���{��Ps�+�=��y�YwN4�)�����K����:8�Q�_dh"�w�����J��Ӧ�=��"��vAfu{R��(x�M�<�Q�5O���L|V�R�f�%+A7����ʞ���M[l:��s�jc�m��7��p��5����`��y�&��RmK7��&�Yyt��=�+�ܮ%l�! ���(��.^9�Ŕ�;Вq�U�#��IATJb n���eB���Qbq��*vW0>w�E���_ҡoa&����˕�1�ehD~�O�D��'�5Hu�m�j������B��1gv��y���C}yQ���id�X��C����8Nl�r�;���|l�)�~3��P�����䡓�k�f� ����m�ѱa�(�wy�����yU�M��t`\4W?���M�x�svN
wc�F���E�2�X�[�����p-���o9	+�^�Gޅ���"�JP1�q�����ro!�������ǜ=1��$z�YV�yi�>ȱ�Ԋ�6m��}gd�eW/g���sg���:^��5���M2c���,)k�b�����o�P��Z�g�ݣ��{����s��=4$��b��O#G�I��(�Э�L�w�+ŋ�����SV��zͿ"�5浤�����:���Ll���ڲc��N�k�k�7�>��1!|��_�_]�p<�,6�K��X��n3��puM��� ���G�@L��ŗ%"����eY����,��)��ڔ˜�m?eΌ��Kx_�*���Y�R���+�Pp�ǹg�r�&��И�2#�؝���;C�������>F�;�?�����іt�
C��R�2 ��0LSK�?]�1�Y�;Gt|��Y��1��o&�c
��c�ɔ�j9�Ҧ|-(ڳ�k�����Q����&��!n]�t[�A�s`��K�_y�R;�O0�2Q㷀���6�>L�)���}��)�ml���W��h 7�>a�]��k�K��؂ruw�(�)��J\��H�)�����J�X6���|��@�o^`���:��x�|���I�7@#e�9�������D%��S�"2�� ���x�z���{�^�`����E��(�z�
�8��}�������	���C�Q�1.��{[�ͭ�9��yY�g�w�7N����o����5$� ތШ~�H�j@%`�����cw�F�ODY�������[K��B�������Yv/�E5lz@��Kdj��=� N��"��Q��$����p�_���@��s/�;獟?�9��HQ����/Jd����ZIur�߄)�h�%�$�zyݫm�' r����P@�=��T�?,��C�:{������C��5H��,���8�.C�b�������XXkO��R項]�Q��n�\�9pne�'fY�}����5�
)8��l/�,�MiƮ��P���i��i*6&�3R�j��-�_8���`���TȾ��0'7 ^�0mGRZ[�����Z"sЦ�E����ɳ>}���V�]�b�e񹞯���o���yj�EP��͋ �r^�NF^H ��̂�-v$[�L/В(�* ]��^n�4�N4��q"8����l�!Ea0p�.��z����Q�w��q�sf�>�@9y���͜%һ��#hI�}�8��Ղ���fqO��o�p�e�D@��HA�+�1{�I�-�uA��G���?U9�3ců��+˧K��K.3r��Zx�~�������}!�g��o��[X*�|Õ�eY	�BKzy�5������c0�����a)�v$��w���Sc�-+/o�Ϟi��h떰�I�H}�d0��Y���-�|�W��|%�W�i��R:���PQ:1�C.��v $f��85�%np8\L��j�Uy�%It���0���3�H�8%�� �e��[��;�I�i}�$ǫG�Y��䯫��U7Z�&>�o��c�t8�z�Nz��-����a��x�?�G�x	Q��'(B!��k��w���U�RY*܆R����跷	E. n�6+H��$�M��":�ׅ+]6��C�g���L�;����	&�v�k4�f3�O�� �P� �(��,�(�X�E��}ʰ"���� C�X(���KG���4������b�"Y���P��ݷ�uꋄ�!���]m$�%t_V�S.hN�D�ݟ���q�s�Mހ��j���/�܊�=��ڏ3|��].+��f�UՃ���b<���8�h��mL4"'��`��E�8�S�tX�@}�*��n��7md�Ѻc�V��
o}��aZ���w#�9�i�7	Z1WUh�
3��I��B7����@<�>hY�(Ś8��\Eǹ\�CJ��[X~����>&aQ�;I���[c���n�C��COB�\o�T�)�U��!,�+y>ؠ�%9�I�G��R��&u��Z���(a/���,�a����N ʨ�f#����|�UW�F^d|z��XuL8\ڭG.��� �HTN5���6ʙ�v �]k�@:��}|�K�-(�G����j'	ka��B�q�\�6`��E����>
%ɋ��M=zgN�V/� �J��u�gQ)9EDDc�s ��<We5vn��,!��@b�9��꽹��9��J��{�d��}S���]d�E+�rl�H�?��G,���|���~zG�� �$��BB��Ӵ)
�� ��7��|�T��+ڐ�9>`���&���X��f�O��K�q��Y�Ҝ�B�n �<�h�6�\����a��Ü�
Ca{�p�� ��`���A��(}��\q���h*sL�{����ใ����3���='1=p�dcmnf=�ʃ�W�O��� @��3W!�m����U���DЧ��S�]($���88�+A6O{����/{���OFW�F��
��/�m+�4dM)�IN��L��;W�RR��t�f��6���`�o��{�Es,��17`�����mJ���{��k�g���΄��+�V1'�kc�<ѫ� �6������
?��{qA��Q@D+RM���%�F�UF��j��ېv"��D~A<�x�D��dH22rqf����-�z\1��a:�5�U��#)�k&"������Ƈɖ݃Txs�Պh�x*ˍ���K��|���� �'��HY=����U()��|���������-��q_7@�����9��O�Ҩ2�]L��§�L0�}�9�1��X(tK�}�}\��.����ږ�4�
k���o�!��!l]�׎�|�	z&'YP���F�|Bo$ϺI��M��!5��\���q�ws��g�b�Mb��{
w�������ۂ8�C�O�}b�޳	�OF�{�L��c��� E���h�s�j`��5ly._��A�ix㭤�i
����8#Z�s�Mj��<"O+�D�\����K�!&�6bAR�`����U[f��t�S��={��������ćx35�HsBaw��P��ghL��L :���g��j�"�J�YӁ$����7�����uh��\�l�?�f��S�Y��nvr5Wj	��}�˚�τr!+��
DB�ú6�[�dg�^�L�#�B����/�M�R�_ބVYP|{=��0����Y��!G/�X��,��-�'	.9�
)�|��E.~�����/~���l��&��6ɒ�(��2�OT�"�f6H�Fz���"����o ��]H̾2Rle^7@
lwel� ��&��	�~ؔT��݌�w�^�e��v���@ A����7�:���]�Ptk�I����J	�q����3��9;$��^\�������'���=��P*��adyJJ���S�iX��Ô��1
^i!h��S���6���$|������Ep�ĩoL�C�i#:_K$7i��#�_�8x��D��Ƹ��(��h�ȁO��M��5�7��Q4�r��}z��K�S-�V̬��kt+�FKK������p�Yajq���u���H��+�k6��"m�m\�J���fiOC���ZY���2�>���mٻ�<۽�?��ӽ]�]E։y�W%]ש�_��
�H^�ѓ����=�R��k�#�S;9E[��� �;Z�g����=}��i"�����Q��2��I�&�{����~�ˆR�e���p����P��f��$a�R"sn��DZKO7޺K���q���ei$&�[g��7�R?������1��l�{���3r�X%JW��;\
uz�����h�8o/Gje]��O����փ�b[�Z�濊:�DBT��Ŗk�C-�Y���+�՚��3�%���y�?i׶��\Q�KZ�TX~�����Y>�Ǎq�M&�KwK,aѻfҎ�r,���֣�1!g{���y���?�E9��Ú�g�eyRMAN��:�F-Q-{�s�r��@KL��'׈�����c)�u[(�H��!�*f���@"�s
�<���-�NT}�7�>�Q�(��RE���,�k$���;�뗉I��� ��!X�1p؃*��H0Jb9;�~�x��	q�/����"r��p�*����J�Y*е���8u�u�8Re'� �D�g��c��| .�檿Հ"��Qk��H?��v��#�/=��]���0)l� �I]��I�Z��&���'5&�,�$-�w��������o)$"'^G�%1�x�h�g�Y����HЭ�������p�D�G�����~�Il".���^Y�����Y�e�'��,���
_�>*�3��=�IP'P����%�vU:�A?�.w���5=j�0~If�Qz&�㶤���&�\V�g,�P|�����O_*��H��,�t>%s5��M�t���{�\� �s�:�j�[Ҏ������� p�h	���Ṳ*vN$��_��Y�m
SKۇ@�Is��
<t��P�y��e�Q���̓b�g�7�Yg�E���Ή�S��Z�x� &�����tђ�'����� H`�c�%b�q�ˏV`��y��i?���#��$.`��V�#�"�ﳻ����yn��E%d�nR�#�E�]��_�uk.b��(?�W��6#*��Ϡp�BA�U�*���74	��2����S��$�l�33W#a�耄b��8�G�z)�L�i���l���h�#~�����?��KKztQ���1�&�^ 8U�#���6B��{���`1���[Ș���Tsi��҈(Ͻ
[�9id��up���<v��규�
�<_���Y�&(`��'G�Z1����I�}��'������ ��
����}p�vָg}�4Z�E�0�42���剩-�郿y"0���!`�$�[��Aſ��׉�!x�M�PT&e���މ�"��<]M�]��n�Q��Z��e~���E4����X9+4�rkt
�
AA��m]v c�7uPE�g���h��D�ޔ�@���/V��
����'C�o<���oB���YIN��!f+ی�Z3����scpB-j��n�\�meZS�7���{��qLd]N����'�{k(Cn\�0��6���Ux�A��\d��auS���:0��{31C�(�r^�P�+��́2Ay{*��3���7�$`$��$ǳO`�}�U5,e|�$"s��3�E��A�@F`Z�s4����v}%D|K+n�O�Keg\�DӅ���yCF.KqC�y��҄��ꟼ�$4����/�S�,�,��]7k��]��7>L��C4��giψj_��W	�Q�L�O�C̤�Ҟ蚀�A^���3�2�Dh����A��G�{�Y~��m���7�_hu_��w��Ee��tHޒ�8�\���I���\��:�jb5���Iu��K��4��&��[+�9�&1��(��7[4{�Y@D�o�^ Xh���X-d�	>i��Rj�O�ac�ΞM�Y{�� ֟����E��A�B�<,�S���V� ��_���Vk쪫���\�j��.�`Fι8�x6h|Ъ\�/V�~`H�C��=K�SF����8G�mG�����J]��z��b�O<8?Pas{X��7yV��3q^	=*3!B���alq�N�U(9e�22�)4'����Hj�yؓ�b���-r��C4�0Ě*0!Zڪ�9�6A4��UHQ�|��ݴ��N���4����A*ę; p���&O��w-�6�Ek_��3��Ep��rm盘[�x��ˀPJ��������W$�la��(���<�h�Y. :��Z�fJC�+���*����D��������so#V��8Dpr@W:�ɛ�Ԣ�����ii:p��d����F�����q�Q:�ڱB����Z�[�F}qۮ,j��Rk��Y���_�U<dZ�G� i�-H���Ԇ���9N����/"�ƣ�]��+�
_*`�g�ɏ�vQ�IR��$�Y��uz���	�#HR��M��g��f�����x҆;�J_Ńr�r�")KCċX�*)�;0�x���h����1S�Wuε	ģ���/�#Ro��'�'W�]U�}�t�Hm�Â�g �g���mV��� *�E�m�mCP��[�m[0�{�V���%��88����K�
hl�[��FN�[��q�м����4��k�z��[������X�n|�
N��Ȯ����P����vy8� ��2�s�W~c��>�H���K�2c��������:S�WA���0�Jًl�]��ԃ���أ��5����	�4rQel�;���s�-�6��AD�3�g4�e2~����V�xG�}�y]�fۀ��m���,��+@����,;���i���G���*������0 㶣�q�Vҝ���?;�)Qt�YxgOb�6~��q��<6��5��>�sY��W���߈(������/��r"́qw��_��E1s����Qc�f3���D���t!�4���FEe&�zTO�pJ1���z�M��C+�^d#��Պ�J����P�he�_w�Q$�C���~�����DJ��&�U7�R.����y^�[/�3��p�P{�ʋv�����������"ŧ���+Նf�%���`��t	��.�Vv�LJa'��'��^Z��]>�qC/������/�(rP�j�(�6x�ϡ���"�?��Z����4q�zdY�,0tB���j�H�@���4:]��K,������.H�̑b�8�.��am�i`���܀H;;���}��	�jF��.q�ɽ�&y�g^=P.eb9�~�n�I. y�m)���M�]�1�y�����<�� 0
d\��-*��?��y
��+�m��H*��aʬ�  _c�p�K�mP�R�j7�.�~���>�8l,�TÒ.x#� ��#O��9`���������"��ϝ:�Y�]�?/O�s��9���/ ��]m5��6B�����:���+=�9\N��?H;yZ��9�����Q���`k�NB�^�`aЧl�����&ܝ��݌�$��#e��^�"L�C+jy�$�{�`�P-g�&s��9�����bT�/�p?�~"��~����������=#x'�ѥ�o���Ō����ͼR�g���kT�� �ٕ��	5��6]�D�![���|���@��a�;��'��q�9͚B{k`�b�p&�:D�Qs/��������)O
(q���@�3M��쿽�v���fp��p��حIYB�`�d6��8L4+�@�~������C�E,m��0�d??)�K�Q�ǈ�֬�O�up�Y���
�ԉyr/H�2rt��J����p��LF<w:͜�	ם�ghV�=V�ۊ��9P���~
�@?5/�Cm�u3��~,]���鰈
W���=_��%�H���:�9��F;W� Т�t�Y�ś�yr���m�u��t�$���k��+�{�Xf�B�){Z�kO�;o2���X���8{+B�ϋ�W�NeY�O�*��Ď��h���L%k֢����0_"���yݸB�#o *_�o底� >��f8�3��6,�j���(�)'��^��nt�^.�%���'A���!H3�m��8_V�6Mǋ��O<���L�帧��$�󑡯�T�~�{H��a� ��4��l��~�ʙ��5�%?��.Xy���;�.���U�iY���P�~�ym���:��䖦�?��֐�I��$F���U�|�_����W��&�����۶=a�����Q�=����&��\��0W҈����1-U�ru��:c�f.5=�_�8�J�,W���ro���ܫ�]$Oŀ�LrL@��nS���?�@1��*$����հ�l6RN���
�L0I��;�fx ��v+o@�u,�ycSz�E<���)�<���f8->!g�`�a�zI�/2�Kt"�jU�<�bx�L�a�>��P�3Z��'�����um���m44ʓ�DG���	�dŭD+��>kAcipS�����-��e���Ȭ�鱿���W�S菹�[-�(~])ح����~INB�5��:�I�&��m���h��f5�����#$���|��|\�u��x^��u٬s�·-���b�u]ż��V�s�6��5WZ�!�]3^��c&���'��d|\����bX����J�` �ڲ__n�+�d*[��0_�vk�����c�|r0�2W���:�;���u*�.ww�"�/8c��Lt|cMk���v�,e�U�QH�L��x	��޹]J���P�X�j�<M��Cd�մ�m�^���h=b�����7i :)�ĖSp�M��9���y�o�^xBcȅYA���U�]O�Z}���+[��?�>��ޮ$�S�9J�����;/�;��Z��qFKq�M/����/Y���8�><���%H�YT�9�;�����Z8�9<^��˛n�n��gy��!��X�y��4�k��\�b9�Oq�YU�^A}��6�	t�G���nxr���7��	�]�\ϭ�N��:"U_�� ���|��r�����9�|�&3+;?��Y	���.&�b�o�����'���S�VMQi:��0��_����B�~<�r����F����
�� ��:�kM�2��n8XAC�*�q�'������Mc<�)�m��B�Qh�pN�H9�b�}�ȣ�,J��#z��BA�ۊ���B&��L��cN��J22�d�������eG��z�����TQ����/�nC��	ő���`I��&uK�:�b3��f�[g�0bD4�4��[Uŕ�<�M�HN_������,ytނ�o�O��d༪�LG؄'��
R"x��D��,ܠ���*A��'�ow*oS@�돕Mm,��nޏ��=�,E�����Z�sd6�S8���ŧ���Z	ط�&�ֻ
%c`e��=�|��STM�'�h��n�0��KB�H�?�#Sb�L%�i���(���w~U����үP��F�0�X�r�:F#�WS��l6�w(d7w�H�z_ca�[�,����X�oG��Ƚ8x#!����Ef>�4X�H�����`>�=L�3�WE�5���Ü��{�+�q��&gr�OAY���d�n�u��_Ĝ��S.�� ��B�v+�6����V�,�r@�����j7-}����#1�<jc��2�BUX8B�u)(��'��!4v�y�S�-��	v��t}}.+McY�ܜl�<�lH���K���h�2p^ٴ9��Aς�X6���.#���G�Y�wٰo� ����.<�o�6õ�)�"�U�a%B�&Im�%�L�<��($J�(D�)6j��Ԟ~�:3G��r�h3��d��Z���}u���{!�F0��;�������JtJ�Λ|�:�3K��K.�'cS���t�]���fԹ�\�k@���g��s��Bp7P	v��$�R'z)e���b6� ����l�S�M���u"1ٻ���O#�E/��Myq��D�Nl#Z=��	,����kX�⧁�$\՜j�]�b�����}�x��Y���D��`�,�=���`]�NH	��n�&��<y�2)n,�nT�OJ����:l+���w9_J2��Ө�����/��i���^�hkS�-n�Xp��K�2���-��?�b��!�A��i%�W�;��}�2�C>kF���.f�fF{�#�)�T��<�]XE��9�ҍ�ҥ�͕�v�]R����j�,E���u<#�Ku�^�+ �5`���_��T��W�.�ApD�SK}�?���sAn�A�:w
�VW�T�~X �-�5>Y��#�INo;����7���g��iqU��?5�­�N��2\�?���CO��MD�)/�(=i��8bX���T�"��_(d�r*8��}&s�xhҐ�j���Py��n��nTƱ�/��>�cZ�L�Fȋa[�d��8���g!~|-aᩯ��;�F0mw}*�Ț��`����?�v{+��b>Vf��f����q�L.-�o���{d��5:�����P���?/�酢�䋞�]˴��ݪ���Z��T�lO�xg�[��9�h=�32��)@���+1s����\��]ӷ����;U���0��sJlbPS�w�~��>i+,O�,�5L=T��@�C�[`~$:Nes��I����h5���[�+O?�y�G�k���5c�����:(5w�0��e�e�i#O�y��Ž�{����lk�X�����T_�W"\!r�bۊX��Z�`C���>ߵ�,V��T���U/Nz���u�����
gb�݀q|)����o�ɻsU���\�Fqn#
N���S9a�a��s��Z���5�jw�#��Ի�uRg���p�ɐօA����دyl
��S�d�C�])D��xdU�'݅��@Q���j�Pؾ)�{���%�G���$�b����Gu�H��>��;;�q�K�<KU��`�&�N��Ϻ(������pFp������h����e\�j�3�X���r��-���,�ܡ���S=EL������4J[dJɇF.ȇfl�������YK%�ť��iOS���,�j�[[�3�bD��Cn�����;�"�!��t�]��a<R���]��Y!2�}Pu뺰���6�t�(�*O-`(RKö�͞�g�q�sV�)*q�('I�M�R]�� eU��^ �as�o�LW�&rz��=I[Ge=�K49�*��bn�5<{�䠆I�����˂����p8�קI_}�6L<q_��^�Tlu��#3���*�;m$rjW���
��I�Ă(��
�ӂ�D��A��>����,��Y|�IH��fN�r0j���|����c2��H_��`X��� �6#�裲)�]��Ұ)n��5�Pt���Ń�F]��d�����aJ��A0��K&-8�=O��_��f)+$�j�뢞ez�{�{p?�
JtZp�޿p���!�׋�H=�`ªg�L�m0��i�t��1W#mץ��(e�r2�źS��,���>�V���i �U����2yu9'�xUn/Y��]���[Y7�
l
3��:)z�R�wq�|B�㉲���>�N�@���c\nTU�$�+Ԃ�n%Q:ʺ`��ȅƵ"%�#�Wa.=�'��1��:���)C�s�7����d#>;�?���U����+����5���7�^!%��]'=!�-�$ �M�����Z�&�HCGt�_g��<S��O�tiYceXm2�Dp��^Sw<�+��J�_���
3�*���F�a�J�Y������]���^*��B�U�����b�f_^Q	|����L�G.��F�N�j]|�X=d:k4��6vbX��;���G�<��D��7?�0ɩ��j��C�޽��G������MYT|�}�~���M_Hz��"�}PA^��c9؇浑[�?B^��g}Z��^a0g�A���A:�k���PZ*��e�d�x�'�]W*F�%i�Yo���K�
W�4z1W�fM��S�&���w�	e+�ɉ}��|.�TII�Liэ@��N�Z��;�eO��J�
J���&n��΁�|��s,��n/5{ܬ2w�k���vd�E����Hu��Wr�q�?�3�C�D�����f$ugq�(�ی�c���0�&���`a�� ��.!�X��<��2ƚ�q��N���O��!a�SD#Xg6����4Q���k�\[�sk�]{�b;��@w?	�D���	h�@bJz��3K���ƴ���������>��������2E���*it��AFZ�!��sr�����D݄Ԉ���d����"8�����j���@��m���s���],�-��Z�H�z�W�5��t�e'�45�����ei�hߊ��x}u�S�D���Ft�lP�TX]�A���BGf �ڦ�2�h��2�]
3�v~�l��/0�MdW��At�#���
�+���Q�0�`�~x�#����6(NH��Xl��n�҆�k(B��ؤ���qhX�S]�TNM��a��K��{����O�V���o�40��"g`0�=|1m�P}^�uK���$ui'��H� �lhTX@�f��r�	$�I$�0�*)xJw�"5���Ư`�8l�R��I,��4�_&�~Ԣ�ІM3�U�� ���@&u=�՚�����8��+�t� ^�ǍzM�
��D�$y�����^gۤd'��s�+ުVՈ��G���~�$��]���#̷�P����H�[�p��(�����)6Y2��@<>˼�s�Hר������}����b")�R fe4�Kh�SR����[[���i�f��&�7��/�,��xW�Չm��`Z<	���X�!�:l�#o����Z�2��m�uz�v��L���ܓƭڦ/�<��}�/f/?d�m�)�ڟtT0�|���7�A۴>�J�4�Ƹ.`�,���fhȗX|� Eb�I$�YQ{��a��t�C!L^��*�Q��W�8pLCt�hS�R�Q�88�_n���ՙz��;l�%K��-�'k�bD��E�
l���_��z��oHX���`�<�I���^>����O�a��r��y��w������ߏVv<=#rň��l|��!s m ��������V�)�!ɾK}���3��)B:����F���}㲅�L����v��UNWx?��8�c�X����?[���0���2��kN�>��xz0z�Z8  �(���c��'�#;�NGB�*�|T��dI�0�b���uʜ_���&H�V(ʑ�Wqj��u���a ��$_�@�=��90u�2�dQS��% �?�8��h��������w�����*⯔F����qĆ��E6�c��n�����JTRnd���'M�?O/�F�5���r˻E���mS���+L@su�|,�p�˙�+��N(�'ΰ>'�-@�R���=��T�#�BZ��tme:���]��\x,�����6�=g��+�i�?���`��M�zN��T����#O�rGO��+<�B���ϪPJC5��k��F��嶻ס��Df��t�n3X�_&j�W���o	��u�Y0�d,L$��f��]zԡ�f`퇢��W!�M�#r�X�n@�����\���7�����s��y��|���#�H� �-:j�uS.���	�+�i?�wP��A��}~JtX�`̮�;,���`y��t ������j|N,X��mҽ�. &q`Y�x����6���虡q�[�W�J�!b)ţ/L����f�(����&)ߧ��*q�������O����O^k^F��a\��f�n�����)@ p�&g�[OK&��釫����Ac>�ʤS+�'�^P���p'	YK���@�
`	�#-��+�WG�����jlz��s��4�mXM�P��W�m����l&;��I<�|:˲:��4�ѫ�
��rūҾ�&�G��`�Pݳ��D��x��l��ٔ"9�}�jbVH �Gp�w�G�'��DC��q��$V�@����|�ŝ�_�dP*mcr[������u��l���3�0Ѥ~߂=�gД(S�O<�^����[�������D�ѐ�ߋ��R<�-T�.�>VWd�y�Q��:l�`E�esX�M	d��&DI+�qY����sQf:s�փ�<{e��`���̀�E&y�9����24*�7΂��:��%����eY�-�fk`)��)q���a1��*�[{��٢S{`�"�#�Y��Za�Q<����w%���>�0*q��rM����VCwW�Z<]c��i���J�'�b�jb��d�lп���\m �4A	�Ξ?�q��d�lP����4/Y<O��c
�פ(�uIM�FʧᥧyO�~�ã���]�O�%L[��_{�$�W��'�Ȇ��	����N�aNzR�����B�s�"5�}�ّj.�=�e�X2�0�����\������L�S��h��q\Q��m��z.5�8b��Z�����-�jD-�
�7�pp]�d���ߣ£��T�?1=��Z
9R�ϡ�|��U��:q*�� {'mmr��!h醔�/Z����Ѥ��l 6PYie�C�
v鈋�Z�P���%K�$�y4�2At�� �%V���06����갳"��#$ʑ���������}���|9�dy��Ppܓ9�nԉ0��I��i�NSHJg/9k*;!�J;��|�:4��\�Zu�<J��;����8sC]ko���S� ���n+�r���SN3��� �W��n�%�ln�J��Ӧ-MMHo����M�� ~TB�i�� ����'G�O!4N���!���"��؛ҬgH��\���e��S:����V�n��I�Vz͚����.(�ϣ%���H��^�?�ٚj�����S�B�#Ӭ�B��r9|e���|qE�^EAw!O��D"��"�z�<���2�}9�'	-�ydW�]f쒳	r7V��d�~.�.��Y�c]Q�FY�?��������V�`E�E�*~y����2Ky�Y�@}����]�Y���mr�N�[��Q`�	�
�0��G����o*	#����{WGʬ���ܨ%Q�-N_��Te*_>�n���s�\�:����z�F���1��F��S)op����w�Nw�X�w�:gX�̇:p��+�}��Bԣ�C�<0������yˁ�j��K��Y�3ߟ�A�,���ZP�3>��7<������F^s�"$�BD�Q�ϼ�/h�,)�1�~��R�yִ{QW��9�;j�H���=�"�f�D��H��9Ȍ<�U�v,�����gOC�&���sDxPi���A�y�z���5�)�|�ȱ&�f/ہ�D�������RP����ަ����S/��̍h޸�=m����<f��ذ��8�a���ɛ_Xx4g��TC�U(1F� f�jH�	�=p��2W%
.��	@��:��N�ɯ���s4$�d9>��(n#c�����E����lPm%�p��Hm_o&Jܝ��$h�4��l���b2����i��沖�j/^mh��nr��WdP>g��e��?I��ˀfA��X���e�=�����F�g�H��m�DY!�~N%�H��Z=��*��H�����ULW� �pP�M5;0X�!�Dc��z43�9Ұ�}�%4�%�$�orL�utwyv�`���*lVj�bz��4�sA{��T��cZ��,oߌ�K�eOY��7�t��@�>Ԁ� ��cU���������Czmz�E~]�%�&��345�8ޡ��w��M祣4I�֓���ႏ��~Q�@:mD�,tSM�O�����"�&�i��0��
�1=����/����+�Wo��v�ځ�(*#�#��$������괺{�����О��o.�w����SIʶgd {a�[�r��m
v]��D�Z�F���!h���Q�Bᴿ4���bu{n�L�1{3�Ο��۟���F:(�lZ\��X�F�>�QҤ4js�p>S	YѴQn�����':F�LeA�GqbPֲ'��#}'��_���Z�J@u�1�#0����U�]xk��-U@_��3�D�X.�N�""A"��7��5k�����D�@�;d���6��Q��d�_�1�ה�8|	蚩���]����3_��dOSTf�d�	Y4�t.΁6/`�L���'�D$���g������d�މ�I��k@��1*۽E9^ ��]������� �W��T��������E�z��g�ڦs�@ݲ�E���\��u�:�f��f-��\]υ��B}�S�u;&�W,�0��.i�D6�μ29����+[5T[pɒ�"�������֠)y���e͍��V�ΟN��j�՜������p}�5W�S3�i��R~�$���:t�)�r����=]r�u�QS�D��Ď�iR���o����i�bW�Bb$���r���*8w�&RUV.�l�&���?������}�a�/[�v�W�ub�Q5�ch�;{����ѱ^;u�Z＄y1*��[��n!B�tm���N���"�Ԡ1u	��������E��df���@W��V�!K�u����Ϧl�`�8��[���T/M�kֈ����a�;o4�N�}�`����>��X�����ٟ6��VH-;Z�7.�B�#>���Y�0@��s�8�n$��1�P޿�
��=-9�٨m�H�1��������!��f:�T|�>f��ae�n�lÙN��':V����o|�(>�%̫���0{�򔦎�����e�>�������9����~�.�lO��1k������}Zlp��T�{љV�:`�j�����P�)^?Q���[�,���r�y�9�q�X�E��\W�m�a�y�e��U#6���x�<Z�5�]���}���E����_(�묿:�6@E:���l��6�s�{�o)�)a $E����M�:5��k����C�B@���2�v`'��$.���E~����Yo,��?��G9�<��O9�%4��헓E�p�9ΠXg�>h�w�ܭ�4�1L4?�ƫ����0�%�w9�y�'��uҎ�|��h����Gm�ߺ��E�X�B���T'YP�e��F�>�^��>o/%&�4L	�u.�X��A;�;�%gCFj*�t����#���jB68'��D�/<l������QB����t&5У��[�z�/�nޒ1�C~�N������K1�`��(�j�2(�����߯o�VM4x�ȁ�W�Y�i��_�*�$fdŶ�֤���,u����!>�BG�l�0�!�U�h�]$���L�Fd�.�		!�C蕛Qk����9�k���!��|d`�˿�'%�;[���3��]N�%��H�C��}v�=H�����u1�0�S���'Oj�Z��g�v������V*�^G�A7��k�Ƃ�#M��<c�l�@��AY~�����@�#E�P�[1�SÅ����r�o�	��c�Yp9N��	ɔ���m����b�J��� � s]x��'(K%��ַj۬)�H�����q�H���P�:`�"TGp�a������BnΫG����¼�*��U�`�"e�XιC�1��eH>��^��IhM(�ʨ�V"�<X�D��;O}(����Lf�hWz�J����T�ngɭp����!���F.�q;�O4��շu�ތ�(�<"t!��
�K��ʩ�.6��`|R5�e �+�O���m�Ձ%���;]�)��1��<m3D�뽧��� }d�����0�E�bǲ2'c'ӥ�=i>�Հ~�*��X�
��c�P��ɂ�`�M�amE���ا;��^�˴	�iw!͘���
��ۙ����Q�\jg8�4�l������)���&�����p(wǃ��9i1��x�����rNl~Q���P�u#�����\P5��JE^�Hz8v���XX"^�ȓE������Ҋ+�Xmm�.��Ӝm��Y5J�;�x`{P��`��S�����DR�ҺC+��#�n�d�=�&������T췰Z_.x�o�6��|L����4@�����~���/�lu�P/�B�}�}��+}�m9䘌�<�X=��}nIa+')$`ߦ�7�d%$���Pv�q�frƐHGs,���1���������M
%�8T	lN�I�W.����"|����-e� �#��~�V^�?=��K�Jhq�s��A�()��R���\�+T��Tzi�2o?�]w��ݣ-`5o�z<2�>��v*��ec��H�ز��c�l����yAR��z��^\���И��s�UL&�)ٌ�v/n��ŸN�����U�m���<�.����9Wf 3�`���ě�>�0�N�:|���pg���@s�d��@�v땤-44>F�s��w�B�:`��޸g�r��Za{_��r���2�;F�x�棓���S�gO��|Oo5�CV ����OK�y% �U<�Nco�fg�G\Bn� �ID��QT���T���wF�0�/n��Dٳ�G���m��3.Hs��� ��p���*|D���=Z%B+�� H
�4����R).��?��\��S��Óe?�.� S!<n~�m��%-�F�S���I����HI0�)`�6s>Ү�G�=�ޢ�kB�$�͕��ȷ�×ܹtLS-N%�A�B����!�9g**`/_Z#���X������P�5���d�H�ŀ�=
M��i�9 ֢FlZB1x"�G�+�U{0x��.Mh^��K-)O��qS��{qm���ҡ�_��vu�3_{^ȉ\�&���\��EAM���/PJ%* ���+R�G��/������4#ַ��?5�� CE���/h4A1 �I��߈-��M�Ng������ �e09��S�Į,"�i�;��|��6{ہ�Ddeؤ{��z��V:���D����1߾��'�\`n^�w��`���}�h�y<��u�A㓙	�EP�Z/Ok�x����|���g�M�ĵ�f���um���5�2� ߶nȋ�x��:uG`�	�B����ס�6�wO��fB�J/��c���6��@m/���h���U��;�X�Ke���]&e�m��p�Xr Z�m;>��d������`y9w���	N�xeeS��B�s��	$��22���5N��e8p���="�X�3�+�@�x�ă:���Ҁ/�����(�g@L����F�G��3Q����
N�O9�X�!YJo&е��p��!���6���E��3���/�Ge@eQ�&��$�n[��O��L��k��Z�M�_\�I�54�7�<Ƕ���~�Zw0�4U7|�C$�7��s;.X�(���נ	�͚a�(���8��\�`����V�]���^a����|��j�}�(n���a�z���x��y�5x�,�Hn���{�P?)���r�2��T?������C<�x ���ͩ�MW�o����{�i#�1����z>�w��1f?�7����P�����|�-C�(h����Ap�.ft� ���D��y� J��X'�fKe}��u�a���u\�m�m���+S�+y��%��
�����3rE
ۋ��h����ԥfC��T6�}\�*�
�����z�:T��R�+�_�D-ң�����2d0i�Z��W�����Ŕ	pU���~�᡿@����qޜ׽�Z���&��
�\���<og�X�Y�I6m�$�����0��{�����'G����z:_��:��}��V8�.v�U�W��k�S,�z�!����LKȝʈ�����:���d�3�M_�fz,����F�\/#��ؽznC��~�Aa��7pR��V�h3���ہ\dWjqG�I�jF<Y���s�J��i+j�\,ēE��]G`�ƒ�qp�1�`�Ĝ�(��m�[D#�B���{�&ꒌ���Q�*��?�7�@��L1�dPk�d�����C���(\��p�-E�[�`o��� 0�Y����� >�U�䵴Z�,�p���������F��%#}�����Q�B���*��E�O���c�~&^��.��=av�D�5�	q�qw.�Z���Ԯк�����^���!��׻�p�w�A��f�a���]��@&�7���#<\@����O�K�XM�~e��5�]�����MSv��@y�Mw@6��a�n�ER4wM�{����k��Tw�G�d.�ʽG��]�
��S�|��(aOm|;�e�|��`=���4��9I���j(=��.���y�>y28�����T���H�)�Q���w;h��Br2Z�?�S�+�rX�Yӫ�s���$��G�mY�sq����=Q���x�1��B�A6� �o%���(��*.�7�e�=�=Ao"� o��e#)קvV(��S}tk�'���yD�619S��X�q�sqk��W�1����-F��j��җ'+� �\Y1��c�Rl`�ƣC���6?e��i��~��[y�y�;��gǻL�-�U�Mk��B��8-q��8�ij���U� �2�8z�� �_N��������I�=�Y��9�EwP���ơfP &��b%v�eu�(�Vh�����P\��-�L�:�k@��ɳB�&�=�m}����Q 𽷗kE�&8mX�y��O3 �2Pq��w3z�ZE�[�"�*���5[����v'O�W���!prs])��YB��2\�#7��2;ED_w39F�6uqy��6��zgM�gP����5���?t"����|��,���׮�U*�/��g��i�89I*�kdL�W�Ǖ�
��L�B��e�!@[wm1E�����!�����ë��_�'�v���:���q$}^�M���]w]+��$���9C1J�4X*d���56(88g.�4��FT2�U \3��_�U��@5�:i.�T�nW�|s�݆exRk8��HCxQۘߔ_�M��Sѱ��Zg ��!����m�M�DVO�͡[���]�����Nv�,��h���?��fv����9��pzt�2�N�UKv����I	�ھ#ɞZ�0�|��#}J����R@����|����+�c�>�U∾���~�xʂ�ޖGmS�V��@��a��у�r�6����#m;!Au���+R[.Hx-�՗!E�J??!,�s���������ౘ2���ٓ�r^xjp @]�0hW�d#�H��8���	kr��Td���\ ���W��)+�[�+<[����PY����y���3������|̪)���չ1�X>�h`��8%�n��lI�ac�����/��L�h�+���s�f)c�x�Dw�*-+���ϫA�ݛ;T���(3�sB���咅�5�+���u�(�y��`�/�fz�#<UH ��,�+�����,^��6�%�f�B��g:��g͘�7�~�g5�:�a��Uy���Xނe���(u��G�g��_#����j�[-�E��&B�G����p堦��
	0���6܂@�tU�nU�� �B�V�ºke"��~ƌ���L��"?�3�.�����4_~46����_u�I�ם��8�2�>��G�#����=�D ��f�Ә���ȴ���zG��b%�+T��"�壘 Z�]�8|8�(n�^f\�_���St�� `�Xk�+ve��)�gl�bJ�Ӄ;�>�8�������V�S�9E׿�ŖK|���A�Y�Ci L�{����NJ���̘@�:
ګ{Ƽ���nn5W�����q/#��l�c�cy�l��72�z��^JxD���G�Y���6�բ!��$��M�����)s:;�e_�x���)�/]`����c[6f�jr81P��{j��k�3����w�ͼ�l�F��/~ /M��U9��2������5�&���GZ�Qz�r٠���&��B;ˮ12�=���^f���k��`�L�G"$}`T�s,p��\���"Ls8���U��ɖ�jqf�=`$֝�RT�����_�Dh��|�$n����9*B4l�N��";�b��T�d0��\,�/�h<��n���<NW�<���ED��jRe��BNE/ K�msrI�-��2/�p��1a��� K�����?�_&�M��f��Z��Q��/ĞEQ�H{�: q��gT�z&��ϸj�5�ɽ�TVs4X���#�eJ}���о��n�U)*��jS��g�Z/8�f�H�]#�
��FIP��H��c��p�L��g�/��g��,'s���w�7�[xKNqb�!���j];j�s��Z��TY�P�7*;��m�lڧ.�����Z��eNg���+}�D�[/�><z[�,��B�Rp{W^�9����������8L���Cjr�01�;_iAu��-5��y�02
kZS,�t4�����U^ə���{=Ib�HC�@�{`���j��W��I�mm��E�h�F�/�x�.y��9:�5jL} ʣ��)m��&O՘5w�D`�1�~|3Ի�jO�Im{:tHs������%���po��ژ�ؘ�_�6�Zo��w���k�v�%�Y�8�ajJM��i1Ca��gd)�)�3КS�H#J��㼣�i$��n4FL��4�Z-C8e�%i�~�PsV9�u=T$�O�ZKq��ín@�K��}�l��9���¢���<0[TՈ��Oa�nő~��^�ωWD?��#e��fw
y�%*�q�-I�u�	솷>v�
8���U�R��]�-��%B��:��� ���6)�=��'�E��5��DF�ro�i�w��'���<2&�[CǢ������)��^���T���%�?�)R��O�K��S�����أ��ZǬ�f����BʧB���H����W�毉�%�ŠΔ�U���5q���H��e�N�j|R�1��)��@����9!�M���ĳ��]O�xSv���B�.���~�_�v(�zǌL���釾40�9�v�<'�w��+�g@�L*��$aƤq�"���	)�9���J%�կ�th�������#�1�fnx_�}$&{��y�����VD�@���x7�fn�
��=��P@z�����$�+���KZg�pjz����m��U�
��-������x���Sͦ5<�%[T:��.J�U����zk������Ѫ�3�8�F�-����:���#~.����[U���*J��;"�'�Lͺ��p��p|�6l"�����}���=�9���"�����a��J�&�BQv�>�wd6*H/��� 8����x�� �_��#��ҥ����{0Z�s�$>��+��l%ޘ�{ȵ�cҳ�捣��x̥�9��%Pw�]�)�����+�<��iS�9[�Fh�z�4��P���(�Ɵ�tX��1W6���T�d�=�� ��ƒ�E��rɪ�n�J��;'xE'�vT�B��23�����7��<1��ŉ�-͇j�j����{�ڻ��V�o�6��V�p���*�H$�GVV1���ۮ@)1�Ƣ�,���?uI�������[?жmc�֘;)�v�ǐ�q���F(��N�~��!ka��;��#?mk �=5�?}�b�YM3�9����"�h��b|�AIW`�sP��*.:8�a�7���Y��o��k���/��iAɃ�3X{��=#1W���S�+44M-�W	u�p�r-��ʻE�C�@�w#���SL��)��(��E�`J��q�����r��C3�׮����Z8�Aia4Ь��qK���<�Ħ�۝썽�MD�ԩ�oȾ��Ȩ��l?t���e�^馛��ۚ�(n���&�+�yO������:>�5����F�����Q|���>�f��L��;$qX����lDL���pc��J!���z�C�H<1M1��梉��LUM5�����	+�����.��B痉��G�E���Y�ߚc����dp������n�Vk)�\w���e��?}E���f�v��&P����Ǣ�v.S�&"B0�Y�Y��ë�����|��إ��'uQ��Fi7�!���������E�AW"�A����2Ttj�rEJ^,��~�0��n����e,�*���{b���δ
�eS��fl���e����ͦ!-)b�^�#@�ˎclW��ʠ��	6{%�4���MU�����\i �O��~�n��G,�\�)�"�>��wB��.S�;<���]��#�L�|�e��nx\��
w3Ӡ�߾G�E����A��lCdPZ@�I�Q�.�ʶV,,���x.�/?�pӖ�y��h�3Q^Z�����8�-$d��U�w�j�झ��/����(�����$�ɡ���Լ���fߡ{2�.r�x6���8U'G�����ʧ��`-�$��_�1DO1��{���4ۭ�D3�4�TZl�=�󛆃�Dؔ3��~�Y�H�k0�j�ҡBǘ����H ��}��Kc�ү����ap�&������ԅ�.{3�ZG7u4@f�B�}J� `<��wU{�_즖-�����Lfe��vwʓ	e~d�@Bפ�^��Zr�����4��U�*.hAIqW�{�X��^'�G�K�\��5 /���t�{_���&����=	�c)Y�}�N�)��f%b���|D�αX�˪��c5��K�j�,���'�
QƔ��Bp��p�Y׼��mD�0#�s?UiG�k��N��/!����j���K}��m:��'Y�)	2X�c*�|�tl6]R)w�]^�ЃP�o�+���2��̐�#�'�4Q��ј �$�J)�>RŦ�Aw��;?�\�H��V:�� c�&C���< �:}���ܿ�k�g8*�}�l���������c@/BP� ̊!e�՗�[PeI��Cϙ⊀1��#�X��u��v��X)�z�O�:���B��'�Bv�Y����=�����Ny�8ݙD�4���;̦c��]��	�&{�59�nMj����Ɛ�-$]0�h�����f��r�Wz�f�?pS�܂�a�*��h� 輯z��%%H��Ҁ�돔�ꏟ��RP[�ǻӸSW櫸�P>�?�\s:LWP��|��_����R���`t.�#5_K�U��(ˉ��(H/Ȋ	��wݍxs�r�'�Q�9����a*��� Qt� �,[��r~��	��(E�W�,��̩��B�U�э�����I����Q���A*��]В�.�ѓ���a6�@��^ω1z?�%u�� �g���O{���='�t�3�\Έ_���ém��ք�t�״N��rg�3z�E:��	��4p����?b�U�����q�h?8ǯW���1}���ΡO���/.X�a6�5��QRF������cP�>z���X+��nP�Ќ��6��,U��,����x�������yn��g�/��$.f��`dmx%�.�7>}�c��֋*�Y�,u{j�aR.�1���[�B����)���N�Z���ؖ��|J���QT�@��}5�2���N���4Ֆ(��q�K��k3(���o�GGd�s"_夣YH���m�E���!�*@@3����Py��_,��e�� ��#K�t�%IK��$������4g^�Vn4埥*Q۳ߊ�@!!��'rj�$�£��\��4x�\]Oj�xX��h��oƮ���Z���(�4S��ax��':b�8{�q4rZ��r���VV�Y�А�WVy��v����@�]� 0���o��$v�ϛ�>��%5�����N0���nӁ5w��|���S�����<f�D�T5m��8�1�ڡ_aW�,;^Fǳ����G?�uD��w׻�"I'��.l�	��?�4��2hs��fE CA��],��W&�ސ�ό�	Z�s?�A�}���b35=<�G{J���ÜA6�`v�:ZK 9X��"6��^��O�xV�I3��2�+��$AL��vjn�P7���� =�?�x��MXM�������D�k��O����R�a%]�3����2�4$́�S���M�>��Z�pK.|m��t	ŭ@y�Q�8V�HL%E˔<��>ȨE?�&�z|u�bϬL�M��������J.+R<2�Q�dZ�����6� �u4�pQ����d��y������|Bk�[�џ_6�O�S�VXP)9Z�_�,�U	a=�DѾ���~��q?ݜ�aG�V� ���?�*$&��q����|1<Z����c˞m�.�>3��O�+�8,��1(E�Q�?�gϫ�+��6WM�bw0sp*F�����h���	(|����m�T��Ab�xmz���}�It?����Գ�M8N�%X�����0���H$�f�>���穄���M�;��,g��\�ǅ���= ��'�%%ݽp�F�3E L��|I;==dH��X�dMZhZ����G6�"ƻ�s-VF�s�[
_��1U�XL�WH�@���|�偉Bѣr�9�S��|um���u��;Y1Dt��3���?�յ;�C���s�����<���^�H.�1>^R��G|&����	z�D&]=?���P�擩�L�/��%�����F��lD=��93T��[؀o����Igwq���s֙L�
�]��k�P�����5�	���{u�iب̀�U��9Nm���
<b�����O�F3�����D�q���Ƣ$*���:��3�'ܑ+���B�tL8[:�ךKx�$s6����W���f��BD繥�%*���}���?S~v5����)��a@&�!ackV\��ǅ�������Hd�^���e�V#��~��ԭ�M�D��6�ϥ����mf]�M&=�ީt�_@Y��G�:�g�+�dH�ZF��1?�.��F=�}`6�|�_+�!�u���-p*�|�vfȊ���T����}uGV��n�����:n�&�8-MP$�{Pj6����޵=C*̛�_=�nC�FGȴ�?Y�Ä���p�9�]m�H4J2֪\< �B�/mo�f���K,G����YǙ���1���iހx6W5�D�tt�l>��i�`�O��U�����T�����K�>G���� �̸S4$F��l�e�Wvl��G��OPwA�P"���-8ٗ�H5!7J}'+;rwb�7�-�^E�����tV�&�,fcI�3:9ԝ�P�&! ����7�u`�*�,\�_�΍����,z澝�{��p�=���gaM7t�a'�nz�eF$g�w���Ğ�E�cy�v�st���L����seh:t��9��H��qR���=zԉl9˒��e���Qg�:	����.+/�E:C�G���n<����i���Y=��d��>�w�4Lˎ��FH�QA���1;Lŀ����(F��B$\ȒJ%��!��
$�����!2���	�(b��u��cM�=9)�d��BA&6^BI��͌b�V�eX������NR�N�~�[0:�`��n
�s�;9�@���6XDc�N?ど�UiP:	 ǜ {��C=B�EzL��`�EZ�@~11����.��Ʋ���'���~�D'���Q��m��F�Ő�������z�!���w_PM�A���Ց�4�C�D�s��G#L_ӍH\J���ϢlBwo�7��ϰ�_��*Bh��*>WI�ףH�x�M����%�Ҭ*��:�i��"簴���{Wx�I|��̍�y4V�?|��hz� �_,�.OV�{�T�7���Q��֝Ԙ,��7K~Ɓ9A�rV�c���	�>As�˻��(���jg��M��7$���u������xV���y���t��UđNo�#�'�6V��;}��A���e����*�1���~�Ha������cK�?.�@$ذw"-�_�9:��S.r�OPӍøP�^E~+�<�h�.ӟs�$6��F�r��޲�����
*F?��s��D<)�X䔙�έK9�ߑs<�2pRi%�@ օ�P�{,hES�������d\m]��3~�0�b.�Pf��Z�'¶Δ[$j��9�[��i?$�'��[�ĬŁr�t]�v�]s��Mc�꫿�_8�x��i�A����A0�}=�2�s�b��u!;�֭w���sWKr�+�����+)�:�+����S2���o/z��4q1�m��T�)�7|��]v�{-�E1Z7@�'�sen��|CF]���
���;{�	q�̕���©��7<s�%�6� w����6.��(���ǔ�n���֌��-+V,�v�����z�w�43�n��u�m�� �h�@��;C���(<��>/��Td�����"�b1��ՍE�ʊ굻�r�4CWȀ]�Uxۉ%���w�:�]��w~&3|�V:�m�[�)���J."��˼vJ��i���B�u=]�Fo���g�P�Nɾ0��WW\͒A]o��4~�"JģBEm�$_�E1����:x�q��_�(��ǯ��;��(��Id�zq��ݬ�3���Y��1�*6���"$�ob���~�\T+LCǁ��5c�.cJӸ��\�޻�b 2R�FY�J��#�l�`������44�	M!�������l�E��A���w�W4��:0ߒl2����+ެ%Bc��ڧ��`�]�M���X��b<�g�n�i�5`�c�S���N�,�̹��g��~�Jt�V�F�\�_҆���y�Cp%��?�&�9�K��� �;G"�� t��O}2�\�c4@���"S���ZਹW��,�k�+k,���%#@�άQ�D�(,ߢ�8�ms��t�J=��
�#�#��b�l8�4����$�'ue{��7q� K�v�7C�`X��A��Y�(��DwBӇo��%����V�>TB�>�	��|��Rl �U�)��c�n=xb*W~Q'i[����a0���5&�ԋ��x��ƀ-�\�A��N�=HE-��/%$	�*^��P�6_(��v���j�=n2BvΞ/�T��۳��+�n�������᩵B�<���y��<��L�
���
�bVzbJ#9�r>�A�=��_��-3&��w4dX�y�Df�8���:�@�Y^��~���gTJG[�W���3�����UwB?Ǖ�s�W�{�WH�uv713�(��I�wp�4_󹻈՘�D=[���E4m�@�?�� ��#,�D�;�ZW�^��m_�G��~�R�����0A~�qp�9��������k�N#�]�����	C�M��Wx�5��]E�����U�'ie�>�D�c�Na�k�n=�KDy�7��t��v�����T.FR��.�a�tgRF��4a*�,��ŉ� D�B��qX9.�3�jQ��:g��K��[u���l쓯~�}��Z(�8ч��m/ݾ�<�����Z���������Ƭ�ڸ�l� �G���o�Ǉ����dHN��$^�K'F	�����;8Ͷ�V[n�(cĊ�}�ص6�W�}'�9�".QL��un�9i��/��>J��Y�X0�K�"]� ��2&_��Y���;�&Y�RX~爺�>�r�V�����d����6�T�r���2-8��r̋��&JM,l��J���[�{���U��/~f�,����ş�#)�1㎴�����P�{F"7����m����8�˞1+,b#X�N�,辍Ĳq�,d?�Zꕜ5.�xG�,a��
�*s�<X������p��O������W)����u�����'���� �i��������I�c���S)&������jb��2e��gXwC�$蚷#+���)�������F�2L)}�&�d���d��I2[��q1>��H������6�2����k{4y�~��&,��4-n���$���`
ö�^�pY����������w��1i�m��l��ث�5�`b3�=0�(?�*�0�h��ts�)y�ʡ��|o�Vt�y�(�����`r�xR�J��D~v}\2�x�T}��X%�D��9��HtJ�͐W{�x��=ޤ�UŲ�`�z��6L���V��[C���f<8�E�9�l;�c��Mt\"�@w�����w�e�HM��x�ikj��Ѹ��k�y���Ԧ��vM�v|z��9�nM��Ӝ��h����B ��G�`�0�ɦ$:�Ly]6!�pG/������t�o�Vh	��?�Ж��{jC��ʼEm�`f�zD����n��+�n�����V�[��f�#����,iН��$a6Z
�-�F�Q^�#v���n���@�^�#	�W�Y�1��ϥ�MS���n�X�F�쏡��g�8��/e��bc��:l9:i3��ǘ# �JP�{lᯍp�����}�w���#��D����g�#4�;3�blAOk	��r�k�Y��b�$V9���������v�3.�(,�z��W���8�����a��[2V{�b	�ܵ�=G�۞�*(,%R�t�L����pq.������c(	��_� �V�_������e-S(G��B1�bQ�Ě�`8��:_	����A��ʖ��[� >V.-����V�׌f�_<G�x�zF�}S�����P�V�������M�)W�_0F���a�U�Z������/�QQnG�1ɆU�m�*F@ի��_�Țˣ�!�6J�<N}���'� 

m-AÏ�5�Ę��{^#�ϟ+$z	PP�䑏�/3�/�x�AW��WlR�05y�1=�U�Ԩg����J��=I^��U�x�A!x�P���Wj��<����Hi.Iu	?@nL��`�.gz��OK�8��$���K�u�'���oT�l\ݸ��E�X����I²�#Ƌ!��
�ܯ�5E#�\�\���[i��3m����9ρ�:�/��!]*��O�}��xq)X�B^Z��u]��c�U�D�̔t >�� :��{X?�q�~hN�ζ;�N����h����l�yr	l_<��{�MqK��0��.�zB�����fʝ��x�"�j�?�()2G�3og؃w�(�z}�&�~��H����gX�d_��?n�2@i�����ZZF==�"\�ul�U��VJAS2D��|F���Iٶ�5���$�G��M22(ꢞ@�X�p����e��$l�R;%7>G��V�<t��^j,)3F�L�]X��!F�N.\���ϋ�jȌ`��*��.����V�!�<l�P�1�!r���I���O�^��,�&}���x�<&h�gܚ��T�[:<�{~C"��/����"Vo��H�����Qd�;(M#]�!SZ�ң�b���p�=h�|�V`��f"X�xPQG<�T+��:�������Z�=���d�5\H���ؔ��ǋ���ͻ�\��lI?UK���������AXf����Ag��j�h@+O��Ȏ�Y����nzt[1D
�D��������_���'�������#Oы`�ėl��Q�6�!����%�SN2v.eFt8�
��Ҡۋ���ٳ�߃���\�d*�5�*�eb�a.���SO㰐�U�9�1�4ۋ�ԧ牟�"}��� ݼ[��ԧ�┚ۏ�΄���bx��[�"����5Oף�̹%G������#�,kW��`^��^��P��jN/�6J�M��p��=ׯe�s��.ş�qZ$W�F&�wa��𵲦fx`K@��W����y���ڱV`u�O��ѭ�hߛ�͚��Ј�@�̳�*��N��:üFp~��*>g��U�8����kz�Q~ҧ��}�B\��nVu������`�6�U��TZ����uK�%}"���N�#�O�<��H'Tw籂�k�`TY�;[X�Gb��w��PcU�A �IW�԰? �Wx6`zx�m�e\��%"?e������y�3���P)���(���M�E�5o?H/o��v�j�ͨ����yv����F��.��}dl��N�\#=i�����C�[��Nނ����қGc��@ѵ�"�A���J���v�n�r�9/��"*�5L�xN�-�%�tו��-���9B:��$���1pHlv]���d��!���IdL3��;�S^V��\����}����*&M�<u�Yvq��[����Z�G�b$9l5�<���+�P���睾yJp�:6�q>BZvu�`�xW�`fD�Y����6z����U�3��&��+�Ӥ����[���f^�"�f^n��������y���{�'L�n(Q�@]���הѢ˾�շ��(����R�2����y^U�7:+�~dG���n�Q%�e��V�d��\��$�G��(�հ����+ٔi^l �8{H��CJ~.�.����X�8��8i�P�R�\�$pLPVY�4�~����"�<eW�n���O����Q��y*�3ly�fU��#V@ix����UV���0���gH��i^���K���O�!�"���X�۲i��%	��R4��"�C<uO�G�YO��� �ΆZ�vS��~�`��vѲ�?�Ώ��
ROd���K�2]Tn(1=2b�4	��`"�[�μg�}�>Y��'�L�u�Fi*(��l��6�����Q<�}�u���%F|.U���KaG���k��>e�6�Ȃ�6�l̩9�<%tB�l�(=��~�c��l�D�:>��FP^"������P�C*Põmi�Q��e۫�k?Јo��)�9�G3 >���%�~A�Rͯ�;VHob�Y��_Ԃ3�I�cj�c� ϙU	�n�K��t$>P%Àh�S1(�X�����j߰./t�҇ �9A�%8,S:tt�yS�#�8�j��)�O^9O\�#���#y�i|�����Ȣzx
�+���4��I����bX��^��E����ý�ūLw9e�)���d��h r�P^ܐ�=bg[4��LWO�h���k�+eӃ!�u��:e�����ב��D2��ZKO�1>9<�g�Yꂪ��Ar�=�s�&8����I���JRO=l�X>��T��8Y�������0�+��ߨBZ�!l��^��RhH8��J ����-/,#��귲D�@�5�J��"��ќ�����x�/�C�����`�i�N~�|�Oh�D�����l�U9����!�ڙ�Z�wDp3��沐�������I�nV�I��_IE����P
�V���j�V�]\4�m�7�����~C�`W��UZ:�Ԡ r%�u?|0�P��K��&s����q��˞�8Xr�;K�mߢK)"�f��m�,�i�b&���V�8&^?�u�h�)���OA�B��zWP���f�,x『��7��iU<�|�D��A��hA���� /1 ��< �h�32RњW?�����8����>L已�w%��B�7~���m����a�öh�OKOy��L$O8�J�`����O��NN� r�w���7;n����d�):�p�YWo*�v����z( -_2;%앨j�6f+�?��6��l����ʧԵ��2�}A�X�ؚ͂i�Q�����Է2%��O,�(�H�8M_�v4�j���|:��i�ǽD�1+3�׋,:��@f���ws��(�����*���o�ǹ�6sj�l�S!�q��
��*>1\] n!k�k��1�|�E�A�"�h�r��^�_^[
��N��q8�ߘ��[�A�_���C�\<Ϥ�I� �����۰{yS��\��7�v�ԣ�"
�qr��(H��7 =����J*.X\&�]�?�j�X(���ń�@G��P�F�~���Q�#\��`�08���F[P�B*��v�͔ I�Uoˊ��ݽf)���� &���q?���Tx$���>i�[�B�j))!^��W`��cNg-�0MN�'ca�߰�1'�QK�g��ґ�q�;�t��S&xMEX�`ʉY�ֆCf7r�ِd��+�i)�����'^0H<�����9"���.��Qӳ�2I��Z�A8����Z�ޟ!��ߋ�F���kH���o��Zi_��mGhmJN �4>Da�?l�݋H�T�����c����[[� a�ר�A�01u�x�<:Alb.��AcH
�W�>M�CX=O�}f�z�hV�X���_%e(��X!3�L����6�CB�2�t}�B d��@+𶼐s��`�3��d�deH~jG��v�ő~g�2�&l���3��_O���oAѢ]>+^��WmSƵ2��AO����Fg�{�#J�
���	%��儨��Nl@�l�\JMV���E�`C�yJ9�A���)_�4�:Lp�ݸ� C(Σ���(�@2p_ᮎ�f���ȁi�����,��O���k�)M�X����od3'z�P=o�1��>]�a!t�B0����k:���*��)�\�e�éW��"1���,|w��Jǵ�3������n1p?oT,�UF6cA���I���}����s�9��o��U�8}|������:}K�Q��/�0�O8�kR��|�\6���.E�T�����o�HwB��o�a`D�XO,+��L���+���qh�_��w���*0��+lBLzu��2�Z�/����,k���e���NmJ�j@T�,(]�ap-�	`oP��׫�X\��:ˉL%�Y;+^�~�LC��¾�&1q�a���L���w�
ďu(,.ȥ��cz�0ͱ�uZ&�H+��(�a���)��i]�_+����m��)X9c���~��5�|̽*���U��t,jBy��p:Q#�BS�Y��:Qvȕd�=l/���pG�w�
#�|C��v��D�-Ft�UŶw�fuz�O�x��č%�2U��8�
7�k<��g�7�
-������ϲ#�B$������8�n2��f�w��	��q��M������f@O�Y	�a;�V�U' f��:��i8B�Inee���ۤ�x��.r,K&�d�=f/���]�S�V]��^�Z�zt�v���@�F�IC76T�M;5�j��=���
c�u��
�b�,�uG��~�.����hF��˅�]�pca-SX5�f1�9�r',MCE�Kb�%�!۞Se�֓��ŹN��l�����ʈ�K�v�緥2�����ֶ9�Z�ﱸc�!S(����[����'�
j^�F�x�%�W`�F��{k�BT?����f-8m�+�X��)x*!�zq�b6.�L?&���6�#sI���Ra������p�|����] V ��N5�g锠�*Ib�L�ƛW��M4�D����)M����������|�?"�őq��bs�b�Z&1O/��<qĕR����o^ymS�ͬ����-I��'x�vS~�_�*BW	6�q�_ia�र�o��r����?��?qL.K��'2M�����䆆O�#A�H�{d���Ս�W��z���8̤���P:N��MaRI�I�x��6��\�ky�:��Gq"�1E[�î:��p\������i-ʞ�3N���Oɠt�U��JW*����� 
=�`���gƗ�Y�x��W�s�1c�l��^��jl~4�O7��!*\��Y�4�~�MY�i�s�h�����y���NO|���� �ww3���=��>��+`cB���E��#L��eKI��3-Ȼ�~�{Ϊ����
�-�e�C��+��Vi�V	X�i��[>T<��-X��c�n��c���<�8�JY���f0��x���.�u{�g��M�F�$z �V�Y��Ks?��ؼ��8����l�py������=,�m�.l�j�0��53��4^/�!��^�&J�]��mer�k��hԃ��ν�����D@��B����f���-����&�[|śz�
��b4�d�]�ۋy�|��ͣ u�����N5��E����Q<D��z���8$󂕸�����|aֻ�R+ZS/�C�Ch��鑦�ex/��Ce&��}ͅlD��T��8ѿu�33�V$�?��l��pC��-�s|�o�f1�=���>A��z�Z���{�C�$���+4�⇏�N`�a4	e��~n��E���S��Ҟ��`��mR�dn�^����!�!���첂������SYeaI�)�p3Mڃ���α>�.5V~�T˰�jS�7k�ρ+���`�+դU��?vx���C���U����*�(pOl�	Qd�ET6�^{9�k��gic<Ư(���6_m�_�NI[��J����:y��J@�o]�6^��R�%��B�[h�D��FB���׽�d|�r�;0�J�iy�.�'a^+"��*�e��<hl��Jj�����>ӗ��1��Z\�Koq�=[�ҦO��ff+k����$�"
AW�^���_��ڇ�����h3l�<&�np��:�J?�[.��F�5I��K������,����ʀ͖�=��	CK����ݕ��$��O/�id}RQ����ŦSu����p�{gi�М��	W�jxj9�1pAc:%�7l1�Pn��/�yȻA��%��� :p�G�Qw�W�\`��dZ��1�{n�-HL��&ߴj�J�WF��^7�I"��Fc[2f���@�܇���P����LV�1b�2y�m�8�l�V�������M'����$ZK �'� �	g�wD'5����|<'
�_���K��d@������єz�"��0��?��r��z�m�����yJ�+[���眾�e�ԇ��*�Wf��"�
u���ٟ�Dba��̛���G~"�E�%�F���~@����y�U�C���G�
&e�s���wI{_emV\S	��D�n��rzMtr�!K���vL�:�J��<	r��c+2zW��ctn�?腁�(C��G, �	�7��v���j�W+$#7�f	+U�R<ƨ_E�/@̪��j�8;�b�	=Q1�0&��,�&�5-Ζ���	�xZ�T߿E�j3��g@!�P�����9bo1�w�^\iۯ�u�GDU���q*{,=���ރ��B�cN��!����lݞi->á�
� !4��t��[ڋ4��̚��5�\��%��Mr{% ��X0K�bK�.E�%(x�nY�V�t�}��(�r9�;�?\������+��nI�wiv6�$�ʉ��7��K�Y���h�Ȝ�WtΩ��e &J�?(�b��tb
D����3-��8��8	'�L����۲1���q�%M�����t�⹔L]���������	u�ߡd�^uz��2��.�!f�"��ն��`)ȼ��={ �sG���ޏ$h	���mÞ/m�t$���/H��D���m2�X-gl�Q�{ȱ�C�gR�c��&��1+���[;$d+hO��}v��m���������|}f��SSu>^����x{*�o�6�8T#e"%�FGl�g���h ���y���` �?�m��f\������,0g�q�	Q�M������^�Ⳝ/��:�W?Q_o�ͣ���L).��A`!vJ�ق���}�`�~�P^��5��I��Y&ax*?mī�u�����8���m̓�s�[��@�B�UI$�d�$W:�T0=ӌ��ْ������_�� �)�߇�wޠ���'h�m�AC6�j��@�X�A�l<��������}b�
�0�	��;�ӓԙ%MM��O·��IMے�k�#"px~ȅ6�`'J�h�m,��5��	`��`�u8���9Z�85Op����f$ J�ᓙi(��w�9*9D�CY��!+u�N�{A�������\�-QR��FP��頡M�O�"ͺ���������ٝ�*Wv�I��:u#�g;�Y��/���\'�,CF��@��J�H,�@��t�r�)�Cf��s�R �C�w�>L�
T�Ww��z���2������F�ʥ0�v� �ey�e���;`Ok�K-'�2�������� � BC��ʣ蘷�&���E�-��.���	\�V���/�/�0M[~i7L`?���Y(<��*4��6uИ�=�*�¦�^<L>�n�Ի��-(��O�o@muuj�}ʚ
�`^G1(��w�9S��נ��0�Z�n`9$w�F��*�+T���������X=�i�A��Ӌ�Ҿ�LZ���CrB���
GMLg�.z��]���]�n!�a�9��T���{��;�����lєE�9O�a6�ӵ5X�G(S���$��Ir��f��IB;�9�tj~�`�E�oڐ8�#�*RF���p� �}	
I��U��s9F逪�M��]��{F_'�������e�\�|�W[��-�Fe����?���ND�o)�[��|_���>�m ��b�9d����CT���Ͷf�I{7/�a�;&�\Ix��{��t�b�	���ҿ�<z�f�~��\�����޾�u+�����/���
7���c��m��\il�(�Jo^��\;YTEmQ���y���cڂp���%��Ay<��xT�Ӈpot�0�>��mp�Sy��/P)���JuFRS�>�$�7����O�XdMi�h�������G�6K�}J����.��2�����[�\g,L4{8�ې�g&�C��ɨ�l�)q��}Z�ꓤt�[1�__HWB^���Q�@H7��EY�2�C(@o�)�$Ȣ�jxjGA�:s$�M�#�P��c���/�����mE����}�%aW	�<[��:�"^�����1މy����D���`��`��ĴE��Y�fH���Ǚu}�]N'�=����]�8�,F�P	�`l�+s�Q+��y_�OZ⯸�͕��h=�o�z�/@I���C�t�;J����z����4�n�a�o�{����S'C�5�1NNP �e��3�=���'JTs�^��&�9j��mgt��p3;=�u�N�'����P�� w��!#ˇ���[�,^Y�aD����dí^�Ȭ��D�~�ڗ/1�O������1/?5�R�+=)l��`Z�����*�{ dv)���ǧ��С[|��x`늶a��/E��SSʰ��D �O�I�[6��Ԯ �N՝�<��Y��5F'��:�ۇl����\��_:o��E�����.���ߕs�Ly�Ȝ��D$����βt���,���2JL�G���fwI��iE;���m�Si:�@ҎoubB[Vw(� ����6oR���@h:Q��h��S������H�Z�v�R�Ѝ#��\�=Ly��w�U�u�	���r��U/��ߕ��:�ׯ����ˋ:S�7���hY��_#�S�G�(�8|�!ݍؼ�nIlFą�d��'�W)�,�?��0�ο��q_k����hg������1��M��U�]K%�fu�8h���׀M�"�3=5Ka�Y���m��Ԙ��	#:�ճW����`�!��=c��������xS��:�����A����«�4��"���R�r�N�UA�U҅
�b�qqPFj�r�9�*Ϧ�Rb�ո�{!����ײH�r)���`�%�у-����U[Һ}��:��:��G>�|{��i6��2�1�,/l��HS���Zb?�NC���@B=U���#��*�����ǋbޙ�N�h�������gURN�l.ou8��<�iy�wE�qב��+�8'�ǕU�����A���#_�u� g;"��W̮*��pUont��7��R/�����2�s��	oݕn��f(��HI��sx~��7i)��ޮ��W��N�����$�k�:�3�Nm*�ԗӇA���I�볅�=ϒ,��U��QTh^	��w����]��[8��AU�,X>~�AR��tlFuh��~�y��Q	unA�pY ��I�Nrg=�pd��s��H�y��g�idN}�@ڣ�fE��Y��5V�M��B��5(��+̉K;��%f��{�"��s�?�`_=]<9�;��о�Dֱ�!�!/b�'��@�G���V���lbw�r��|�������HyL�25S���0�A�ʖ����۠lM3�H�!T]�}���[�X�v���J-?�$t�ᬐ(F��9��X6�wO'�,%LO۔�Z.�άn�k[����D��`Ma��gqt?c���Z��$d��b��*�և�6)Y�]˔�T�wk�p�U����Y;D�Pc�f���Wϴ�;�<ϵ��*���)ϛ5��Ƣȇ8���wK��.xG�C	��~w2�g��d�c���z��4�,�
U�	lc�A�a}�.��������SL
3\X��qL̽G�	_k�ꂉS����ڈ�ޱ��uF8������_i��Ϥ�28�1�Ӷeĕ�|;�<�ZDx҄�����2矽����x���SGP�,V��}���CJ��C���ڌ�m�v!�����ǌ�YM�ߊ��-�N`1c,H���=��Q��L�ʅ'S8�r��aS�R�*��n����lg�cc����>��:>���1�j�`��)T���8z'���mt�?MP�%��V�QJf���K���:��l���#�k�K��d̐%��gӱ��b%��s�NR�s�a��@�F����uU�eڦ7[R��
g�V���Qe �ΰ�U����~����@y9����s���65����CS
��3o��{~KLl�6d �; '����4�;��N��^
J�q�����p�z���B/V���<�H�tM㤈O#
�ثiQ2w�	k��e��T']�u}��E���b~q�#F�nz��lY�No�r��Oa�^;�aP��N�����Z���u��ȗ��Ց8��p����}�r��3��v����i�Z��G�c�F��N�0z2D沦���i�FD�u����hw�kH�N���a����5��ii�("�:?P�t#�
:��OC�*;4KO��A?�`HE?h���]d3KA@�Il����'=פ~�� �.#�v2��ocuAۜ���6����	� C牪�TM�����x��i�d�m1�����>���Q�P"A���m��dD�rbR��6fG��ZNm�����yrD��0 �(��T�>uHvǭ�r|�X/Oj�j�޹�[>(����,�M�G�X��l۩0l�-�� ����yܐ����d��}nDZeB\U�ȯ��;�c�)1N�s��D.�������߀X�VQ	�z��8�ֲ ��;G�����	��8���~�CI�����<3�?B������sWFs�%�%��^�k5��͂�e.N�b�]�� Z���9�tH!��C�=�A�����Q�/)�q�pf"�}V��tQ�;��(zVυ�y���"�i��N�O2Ai4�RxT�S�>A��m��P��ք����PT1F���o���8a�_�Wd3�NQ1i�\&������K�Z�>��� Vb�?�gZJ�B�����|bF�`��9�B�|��o�J�uLY�N"�/��Y�MU��|{�5)�0^�e�/�&Y=��݂!�rp��#Yf����;�c��)�� �������M�=������.*~�7��YXL�:���B�O\���D�o,�1�D�<��:������v�4����,6$I�����z��l�MH�?���uU��y���b�"��0��j�����lK�����Y�B9�iՏ�+ @$u��۔'�~v?�z-�5\����V�ī����{��Ն\*�-<º2�F�C���HG��Q�e��UZ#����A;�g:����YPtv�W�W=R�8�z��&��ȣ��w�溛�RS�8�(Яs���}rE͠0���*���'��S�_���ִDo�J���G$��u>�ϊFv,rl&	�%�y�B���w�b���Am���|����"\<��c�n.`��k���r6k�5Λ}��[��~����rFF
��p�O=���� �Zko�����y�T#J�13���4��@��^B��u����ɸ�}~I�m�)]
g�5���5h��f������R��;��k|��e9B�ަ�u��O���(y^7/^p����7:�lR��2wֻ�΋�ƸP���e�[��c��,8�������1çգ�j�6/j�@�ZML���5a�n�+�s��	���G�&�:��.�d��(��OϿ��gvg�Y��tC��x-� �s�۰�`J:$#9)Z��SD"�7���j�;�	�Iݐ�m������ְ����&r�2T5��Y�Ay����j�<��V'��R_d��!��nF�-��9�t	��g��uA��QyY�n�"�K�T']����'����K���J�$�Si����)�evװ��=D��PN,�&#A��?L�W�+�s?E�a������?h��{4'd��ߕ�<JR�d�I9�r��?�
����FD�~j�p����Ŷ����$�9l/U��h��:P������b��$J,ft/�
Ֆ�h��Ip�OG�����H�X��NDc�eY�F1�pA}k	)Z@��8��>_�rÍ�(}Y���37�-��A��6{���d��@���.%׭���_}�H���pu`X�}�=�v��A�����% k��,� ۵�|�K��^Jȸ�으A��hU-��t�	�����:��� �npL
r�M�t��������,�	P`H��,׭_W��>3 >�ME���B��ڀD���+R���bp9�y��::p
��9I�	��y�)���ؖQ�6f�y�նp\b���JZ�7���f��g�w�H��>���r��1��Y[���*_]�4�1�=�G{e��A��W�T�u�2��_j�i{2t�Sۚɮ�%O�V2��{��e��<_�8�m�\��ӫ����)���W��S[���To�\�j�V멋/T�9gD,����<y�}���cS#��{[MT�*�t�� ���'5�����
���:�N�W�~�]j��K�@��y��u9�X��^�%pJ��I�Q�;ڐ$D��
� k��@YʶX4[�Ӷ2�/p��Gw��vWh����[
4���O��հ�&���������,$�r�_�D{v㟫;�~p��aa�w]�ԇ>�-+�����/�&��73\C�܌� �95lc��p�w�gD�rs&~�8:���f'���!��� H6��n|��u�9m��t`����a$����Ss��Z/�Y�.o	��?xsB��X�{����R^�J���O9猿Q�Rǰ[Ѡ7�[�����C���%�vbž�	��0��	���70�K�𗾘�_�5�N�U�"x��ڣ��_/���@��j��雈�֥�^�C��/�zL7\|Њ���P<Q��D�ChN����n���U��}m�Z\j �i��Q{�%$@ߍ.,��49�,n�AV�숀t�倖*��T4�t��������S��][��!<�Rs2[�zc�sԤs������Ч�=�m���W���n�3�3^�oF:�/I
�ҽ�z__iE�ߤ��.�1��3*r��o�&CT����ܛ�p��{'sjxGIMY�#C@U�q�G�R�L�ʣ�O�#�q�g��D��	��m���I�k̰���3��s�[����P�hˊQ �I�$��`#���u]��!�U���PD��}-P^#��%N�m�E�t�@ի��Tړ���(��ߊ��QQR��ۊ�mG�J��A?!�*.�Z�4�ș�=��\�..�XP�aE�G<=�i������g��$�+5%f:J�bt^�"��M��m��t3|���^kA����/�fg%�S��Kҳ�+���:7�P����?5���B*��d6�(Ќ���|�@2�
yi���]��}���!�-�uݵ_?Nk-�s�$d"�9�,���18wr|��,�.�B����o�|�3*��?��2��T�"L�u�O<�.�ay�1��(��U5�������t��oM�r,̚j6��j�C?�C���:y�k)�AK��6s��o���2+$�1a�7�ޕ�̧�l��|�TGf�w3�����@� 
.�5\?�]A��gYe�[D���5���}KT���p\�딡�T{�:�'#��`��/�s�r�',�^�R�L��4q�����@ɎĪT���Ӎ�_|
jz�H� o���Y�ģB�WA#��o�؃ǜ�y��+��76\0m���Q�+�E3_�B��(^�;���2�1�	��Kᦽޗ-Q�9�W�T�͗�r; �4ݎz�����J¬(��f�$��:KŹ�8�kvg�h��N�Κ9���X�:�=>�^����_��#��~BE6�v\���`HAR�K��o&�;�܉�-d8'39��4������S�l�m��J�S\��G�p.ˊ���Y,6Ȟ���WQ��P�8��EtS}o��C�O��' s��zZͭ�O����%��~נK�r�����-\��^����������6F�Fjv�g�pq���E���a�p�U����m�g�� /Ǩ��n�J`�>���7� ��u4����K[���Z�I���D�J���W�/9g��>6_�2T�Uo[ƸD��Φ��n�\r n�s؄n̖�%�В*Z�6�B�2��F�õ�l�bܱ����w��d7\Ͽ�>�p�����ٴg�v���;���j�Χ�}ɴؕ�9AC���Pe(�������r�pw��9=���L���S��T�,��T6u�h�`/���3����C_G��`yS��M�q���/5�n�@��"��U�]�?3zs�����7�h�[K=��ȿ?�Ა�Z|��%�\
v L�&��a��d���S|�j(�(�k �YU�|���&(xzdv/M�w�~,�*ā��x'
Pt�� ^Y��7�i���H��45��F`������'�XfH��
�ZHYs�J^O�rYfkq��ڏ�q�䋠�c~n�i�� &l�#���om��>r �U�C<i,�jᥠ�:=
U���th'�9ED�m�WqCyu�K�b�j��49�F����d��?�b�,@0vp��0p糆_�I�-U���������+�i;����[���9G#�of��	�qF�	]b)}�W�=4���џunx�S]:�W/�ـ�FW�3�=��rƯ������cP����vD�z��#���;KRP.�d�!|��\d3��Q_rܣ��j=ʻ�`�J�?�c0�F��`ީ��b�������Sf4�vX�{zV^=��S:Ǡ�{�H/u�����G{�-j� ��|�����n�X.I���i4x �t���Bn��k,�"�V���e4?{0s����ߤ *�x��y�ޏL僞�����X�٭qIrxq��ƕ,Q@a���N�}��7�<�H1VLh�5�i�V��z#�ud�K���{>r?g'�3�{8�ȱZ#��C����⺩�3�9{�W�􄶛�O�C2J�I�k��@H�,��'�.��ٛ��M(�<\�����V�"�ƌ��Wmd�B	�)Y�/5}T��_	�q$JxJ��>��8�����Ò�3���㣠�^q[��A�>m���B4�aL�İq��}*$.I���M:�3T����J�*7t� ����M:�P%�&�Bީ)�%D�S��Z�p|�jqhe@\����7��O��e4�~_6�׾�v�LE?�����ǣ(�7����Qwb���b�%gy�j�r�>
LAȲ�5o!@��29��I�g���^�HH�!~Pø��7'v 	�*�t_�<�)���4����Փ)��j�I��	�7�_0$�s���M�A���A���N����k쀣�m/Q0�Z�93��BA�ܺ�ڼ���'W�caH=5tE0Ui� q����=\�<�u��0=���*v����I���E|�?��U��Y�X�s��W�����ؙc���ɷ����k���}�jm�����-���4&w8
��e�r�_��7\��ε �;OIc�����c���Ii,��Nn�K(]�iO���&ʘ�g�v0=C1��6f�g y�Q����8��?$0�V۝�<�k9�
�S�	�>�����3pP|��h�N�Jڞ��͢	F/��hK� �;�4 ��F�͋2a}���eQ믹6$0���7{��t.��;�a�T��T��wj�H�����p��wu��7@��~����U������G^Ԯc��<�2�LNp*dş�� ��H�QEo�',p:���AJDh�͇�����̗;2�ia���۴�We�^�D�ޢ�AMH�Pْ�e��#!�A𧎝��:��*��8��R֪ ��A <�����񔪭��=~��C�P45��x� �����\�_�_�]hK��6Y8>W*�
l�^�k�>\�P�>�M`���̤�*��WM�r���+��=~�p�_�s}��k�݇WK{�Y�e�8ZO�9��N���U3)��S켨�a
Tc�xy�(��޷��އ}-��GB��-����q4�tA�?��������\��kg�����h�7� K��t�E�����b�r���-�Ck��%�}���M��A?��zv��钿�d�(�Q_�;��N�B���Etjv5!ԧI��7����Mj�9�ҙ��҅(�%=�����V`y�㪨�T�n_���QK5:?�-�֬��3�~}`=�­�G��}}�='QO�k��E��A�i-�%�Bt�[��D;8uÖ���N�N���{��7�k_ه���4*��.����mF+���lDI5x�����2�ٯ��\Ȣ~#ٮ_bO��(�Z:��Β��o�r�~�A�v�<����Q��\��@��[���w�����=K���@G'���f+w<i�g��Ⱃt�[���	����-L��jդ#�
�V^fV���~�2��7�S�X����崣7:���,��/'�q-�B#	�����<Pic>y�S1ܝ�YF���*��A#��#�L�������XF�_}74|���'"EV��u������ƫ�R���9Έ�:� ��B�v�T.���F������Dq�"u���ʝg���p�4�����t�U�X�$�8�����;ېaH�h��,��ォ�`��I��ӗ��~|�>�"����6[�n�ϐ~ʏ�.��"P�㚗jo�ӭǲy
��3�"W�B�uWb+�� ���$�� ����]o�bI��O�O�c�)�az}�S3.4����L�͘���f��C��	V�Ƒ�~�/��>>�0�,��V�9�*z3�;����]��1c��>�#>�"4i����o󗛣)�A��bRr��ʛ������ƣ��(H�ĭ�Y�[=ƶ�;�����h���q7�F\#9u��KK�^�զ�IG��t&'�3���iOӄ����/�kwh$EJn�_��Hؾ����v%��/���	�r����50 ��>ON�	�T?:'�v�ڌ�n���+�=eD�>��9-*%QEDզ�B�V����!%�h�'�����W�܍w�"֋`����2 �����y�<�m�uϦ�f
��p��x	5>��8h:���-UnI74:l����NFйT(i�$?�k(�+�M�?̷��\�k(ުJ�A�V�"2�`���g\�A�8����^�n�Z�����pXm��>A��9���l? rLp��d'�-�Ztؾ^8�����a���.�f����̇Q���h��R�E��#�k�Q'�����Oe��?�����H3�׵N �3�ko�6:���aR�Ūԏ��6�R?�F��E!� ��]m �ۭw���GbP�""%Y������̨H!��i8�����61g*;d�v{��y,���^
��F��0�^K51iݮq�f������(�%�j?��T'�0/�~*/AR�����M����=~;E�3�ߚ�5`j�T4��Bi]W%�����Ʉ�G ���?�����ԃ�*]�����FڷD!_,w؛j�r��η�B4`�nl�d��"��Hؔ0v�����#Dj�:N�x���T� ȅs:"N�)/�$��KK�Њ�R��T��vrk.u��f`}MEGj���ꎏT���h�%���=�Քv]�%*��%8�B����XF1߅��8P�e3�8>�f���ژC4���2"O��V�l��-��$��W��8f�Fc��$.-�!Y
C/~(� ��9�P�1,�,�|q���牁yX!Y1�n�ϫ�c(�uD0I�/$�CK���G�PN���1��}�N����?�(�N��%M��wY��Ϊ�Ih�x���XFo���M�:���5؞�fD�@�L�[�sڄrk��~m���V���wTu;R��P�Va#
�׸S#��K���I	�"�$땋@N�ɷ��f�S镅4��a���'N����'-⼝���ؿ6��˧��W&��#�]OdY���h2K��{�{n���qI�6�J�OC��:��6:��5��ˣ�4!4L���@��)����W?��ң�r	�~*:5���m!:��ʹ¬��� J�4.�nM+`�${.?�.�9scK� ~�~E1�-�v3'��2�hVΔDD�m	��2��E��db 6��y�$�C�P�e!@X�m��xAK.�pb|E���v�����Ԭԗ���O��� r����H-���[�Ja���y3-q�I�?���@ �;İ�r�r9,i�0�\Q����I��(�y2���0�nЊ�&]w֗j���H+�n�4���r�6����R��֐F�e*8��6��f�0�0�8�?��
d��'�b�'���-�c5S����M�Y���s�oc�̖�Ӛl9����N=B�_�Hٖ�]��h��K��X�=��I\��t-e�d��sw$EX�-9�r�/�]���I�0tyr�������
N�7��	�b�﯅kC8���DT��4�ݶ�L[�R 7ڭoLE�H��C&\������)ֹ�FQe�����8.t�s�^V��E<�,c�����:��X���2�����i3[w��q��)����-��,���	m�*2�W�L`4�
�T���8�ZC@�o��cJ��	,Q3���w�#\.p�T�ȯ�XS�>��mg��^բ/5F.A�	D�" i�Q  |� �l�x���*:I���R�i_�0�ar�E ���i��S�͙����������0�_�U^Y��[��v}���t�)�Z������<��n�=���Ûl�H���eG�%��بhܳdZ5�Q��^�҄��Ƅ�̇�]@�CV�eݖ @Y�b���ϲ�>�Gx���w@ֳ�q��>�Q�>$O�(zNӲ'.N{��`9\/��2H�w���μ�w���ٵ;�R��a��GY�5/�L���U��@��M%�WOB�M��-��{P�J4�~ &K�E9@���a�l�^|uj./?�C4OB}�V/�VE@X�3��� s��o���`����~Ik&���U-Oŭ��A`����o/1+�B��O"��>��,D_�ö6�Z���~ih��a��s��3E��{&!�����1V hx�저��)'?��� ڡ�k�$�c/��]�����rH_� �nx��润���Y���X��L�R�ex%m6��k3H����b����a_�}|�83#I�l1�[?��~�n˟
��J��rl,I�D�:x;��� �!�2B����&�s���^a��D��7������/���2��9���(F&�ʱ/P�R��PFbY�(�Fy7ʁ� �_y1�8�}��*Tw��4��y�jc�����]���N���r��\ˀl�P'�q�)Qs$p�2]?ؼW������Dh��UvR�n�Γ����(���M��"��n�W�X5�Bi��Q	C���M��KJ�na����Y?�Wr���pﭑ)l��k��|�`E�n�#�]79`��u��F&ٖ��lN�s�\���6����4�?�{z��6Y�!�G��b,�F9�NU[\��V�MlX1ZQ��f�I��eW�E�����&WP�?[��SxT�:h�����'8V�PݰJ-��08��~®�d��� �Zv�Ҙ�ϊ�K�ޕ�|�q�����)~�e�PN΀�^����!��ऄF�%��x�ы�^�`/�+o)g�O�=�2]��(���"Ó�m��%'?��F��HT�	CzV��tH���˺�e��`�y�I�SXE����O5P~Q�� }`hH�N��$τ3�1�B6sT�R����iY��a;PF&K�),-l++�}䒷Ga��_��H��dŸ媴���'|�o�{3�'����K~�UT�Wi��)��ގ>Uʹ+�FT�+�H��\���N䷅�x�H���11?}��V?�b�{B�;ש(�sR{&h���?��e]1�������VƳ�����'H�CL8
A����b��v^�	����|B�|�(F/��BCt6_�d�#�h�}����&6h5�e�
>v������/D���KQb�q�>��'����T�L�vf�s��4����I���-��#"a7?�*��?vg�F@Ⱦ}v���<L"j决�y��Ǯq�N�l�����N�1X�uI�Ŀ	N���7~���8Wɋ|���3�tM�)�>����u�U�+���
�S�y�1<P���1*�/�G
݆�w�Ben2>�?��l����lOT�>��6�iJ��4��r+f�@#����:���\ꊘ�d/C�����8�&����n6�g�	QїS���r�&؎4r��h�x#;o��H��V̓��9����>Z�|RY��I���)���>p�r�Ǖ���%�*�l�(� �O��puy[1Ly'�a���\�(u�B^!v7������q�_CK=�ۭ�r�e��e��}�ex�j,�P���i�Dw���ʰ}�\#AfȄ�Jb����l���a��S��saޘ"���m��'�=�JS��o�3#��`������0� TBV�ʗ)��s�M-�40�vU5�j[��n�Tg��J���o[ڝ�	ފ��P�<��C�r�$��Vf=�x�=2���/3�ي�3C�1��~n����e�1@Ȱ��ℯ�dZ��>�޳w�hR�?KRV�Q��@{�+��8b�@
������/�F�ix��'RZ`���i�|?�7��׃� H{�	������. M���_��#�cr,��⡕���떿z�>�Y����'�}�/����|�5�����,@[�^��/�������C�$�d ɉ������
��cg����g~���2�j�l7�
�h�`��
7��l��
��3kE���_ӑo
ʗ�wpn[�HS�yTEI��/:uu�fi� ��_T-�S�Y��N���`�t�<�Լƚ�1,!B��Z:�iN�{-�+h�� R�eW�ڪ%�l�����(�=*w(�э`�#���i�/(~k��K�@2��ȴ�E�ky�I��6�X�I��h$_��}#����j�.��.�I~� ��M4�C'�M��Q&�����B����{����&��0�'d���Y���gP��s���)��˧})�H���;N5�M�i�Ʀp`�
67S��K4kk�]��Ջt�\�>D\|c�ͼg�8O�d��x�#pf`�	��0��O�6ͬZ��6q�����&��b�?���bM8��><��r�y߯���ʩ���4x?���d��R?�8��5��:��l��rV��36���/���A?k�D���~C%��%�3m�������Q���a��k7ؑ����F��T����ا������u?#Է��(a{p��FD�"Q����x�R������Ҟ�^|�R@��`S.���h�pi*J�B����V�D����Q}�ğw�<O�N�?	ˠjE��\&����O���A���wvQV��bL �W�=�+��E"�G��އG M��-�	��(�D�u��`�Y�u�8��_���1.u,�n���?��"��n����������#�`�kJuU�Je�S]�qx���V���KkEʯՏN���������Bk���$m����.4~�9�U}P���� w�a٣���x�?�զ��n`�K����Iܙ�,��dzLA�7cm���$�K�T��������3��׆[b�q��p=�˻Vi�Z�m@������N�#��T��k�>D?����O��p�o.+Q�%��UE�_c��R2��i T7�N�hШ���1Br�w1�_��������_��$Mv�T����Ƕ[�wf��I`����f���W����?��z�X���ׄ�	6[)<������CZ��9=;��I�E<�R+=��GQx=������	��y.A���{��m&�Q�'x��v{3�0��
����|�O���?��?X�fU�V��j��]^9�|,�f�,�N�U��?����3� �ٍ�uԕ^S���ʐ?��|)��0��c��C&��%��Ѣ�5����`Rϝ�Aꢫ���?�Q�ӳ��!�����a`�^�����O�y �[��g�a�v����*������v�IY��}��U߭��0���R},� 汿E��z)<����d�3s�J�^q!<�_3x�5~I�L�	��m����������)�=����(�m��42r�ղ�j�d&�kA}�	oT�v��d��i�}7hc�T�r&3_�CѾ��{�:2X{ZO�>0���^�o�Y�����Y9q��J  t*O5���ʙ�b��hhr�DH�5�90̩��Ö�y�.<O��@ݠ�&��Ѽچ�H�kT�/	>�ڋ:%7H���h��*�}Z�����@=U�a�' ���۱t���/��	0�u�m�����%L�`76�� 6(�L��Oը��T}c��Dޢ�߼p�'�F�S0�g�+U<r��=�x��7ͣ��������R4�[�~
c�R�;����I��}�%�ݼ��gc����Nb��rb��%u�%�M��yɱ"��z2��ay{G�q.�7 ��X����4f����PץuP0}6k��=�. ��=d����m=U�-mD28�]k��冄�'% ���>t,�W<�Sh{ʪ��͚ki��};�cFӪ�!�d�k(!�AHnF?4�9P1�Iz\�?��A���)��u1�C(���(��I�šc?�l�djS�5�	C��L)���K�����B��p��P&Э#H'�x�A�	n[�I��P���8`ɼJ�|�|�n�=6��)L���o���c���Y�u��Ws��#瘯/i�H���x.�7�*c3�ؾ���.�(y�4�a���Ȍ������w)�;��
�a�$��K��X��M�49=����5�q�\K�]��u&&����f|5ʲ	��9dr�X���ZAgHp�|��op�G�������Q���N�-rH�.�=	X�����dt{Ji��`�G6���	�����C���P1����{�X�ݞ=G�z�Q}0�n剾�6ZL
A���\���Hh�{W����>�1-���NHjڰMO��D���C��E�Q��i=�=^���	Q���.��) �rb�ۦ9�`�,{r�Ț=Et�ڻ;a�s�mhi��,o�A��O/�.�a�#�k�RYN���JX�֡�Y$�����l��^��.��%�u��ǺOZ�@��E:�Z���/{׹�w!��T��ƿ��χ&\b�t|��o�j���=�=4R��Y^��]�خ0~���ЁK�<�vBK�_���OO ��n�,�O$x(���J=
N7z��S�tiV�ʲ�[&��ynŤ��b�5e6z�@FjCG�h�|Pg<�yU|)ae^MVepU�,R)�=��p�"���E�����2�94�J���~i�?bR6���J����]��B c@��l��]Y�[En��K�P����95P�z �{�Ӊm�>��&pFr8����0S7�z 0�dѭ�ƏB��R�.1E�CD���0[��3S#��o�FnrT�U-�ϵ��
� �K ���8���@%!s�*�8�4iԋm��HD��սw$s]�D�2���[S��=�7�f��$����Ѥ���Q��&�^OR)6�����ۋT�oL	J��`�L7`�J+\r�\a"���;�m������c��m.~'��v���t[�1��G��]8�bIEhp������.+z��k�t�ݚGxA��"��Č��ymMd>f�����y��E^����9�h����V>�e�U�#����	Z�6+c<��K�F�^i���O�Q�e�	�(_w�,�2�9 [�ݥy�x�H�1(���ƣ��[�@�Ք@c����7�z1<�e�oI���_�{r��d�\%��@��t�Z	���QX�\����^���12c�Δ�JjF�Q�-�S��ԻX�I��^�g�W��}d
F*x���W�a���YT�� ���,	ݯ�~e���4N��a��@ 4Be2v�qd-��	��Q���w��%�����V�I�nY"ڵ/�&P�Nо�j��j&d�2F���%�e��<�A��*�#�d�=uNgH�G�AP�g�z��<(P�.�hc�5Mic@���q����tQ�j��V�>�k{�S�\;4�P;��G{��'E;A`�TVs�7��5߳Odw1����bt��P�s��ȝ=*��%��c�c�G�L�L�6I"�);�J����Y�n�'G� � |U7�ŵ��	���OM6B�I���'��@{V��I�7xq>�rg^����w��[����D���Z�[o�7�C?M�`=4��?MQ֤-�sԇ���7�K\�c���!�Aљ�_MhV�}�^�9zU{jϪ��_���@O�q�~&$�s@{ES��R������U�}ZJ� 
Q����`�w���(r��\b����i��� {�޸�����}ĵ֏�YOQ!O�#��!��L�5A�I�_|���;����(�4ъٝ.�=c*�,�x��ʒlcl7����n�*B�)(6�	�f+�v|�ǒ��������@��l��N�T� ݍ;F������$q0�*c� ��K�����=���*�*>���IώS2MU��5���9r9���Y�bN��6+�\�1J�|�_�gDZ��`9�\TN3AcM��Xs��&)��zdi��w�!�,"x�Qx����#0g:g�{���%=%lZ�S�	
U��U�r	�B!��em��2��z�\ЭF��v,�eU�UM���6(��(Jw/��!φ�q;_w� �X����m�4�#�~�6�����?��ݙ$�lTn���w^�g�]\��4���(/"c�/ c���4�����l���Sq�4ρ]F?�!�I����+qD�0�SP���.y)ժ�����7����2T�"ٿFo'�O4��� ��:�Ւ^���5f����ԛ�X�Rj�,#����J�uY���lB1v0��2����ǉӴ��^{�d���;��r�S�#���露!�Rd�%���?�?D���ge�����G,��������`��쇿ltw���<"��̫�����[gjJ�Yjz�	�d1-�
d��GS,7��덷ס�!�JARrF���N�\�i�)v2�NgO�9ނ?�m�Q0hm��P�	���$��x��;�s�M����4(��|\Uxu��lCy�3�����"Y�j�4�qc�4�j���؏�O�� �|o���U�`��6/5�����_�}�L��J5��,0IX��}����c�^�"�w�Z�F��4�!�.[&��5�c�����_�����0���60U�G%�L����#jLu�{&L�P���Z���٥<u����㢄�a7�����X���}�H��-���-�(I��~�4[Q�g���`x�m�ߣ��K\.L��5Q!l=���E�Z"+�T^��67j0�x�R�/��4���(���M�����e�ċ����/����D~�)�}�^���<���|N�_#��M��#iU		� ~<d>�%���7���2}E�P���
#�c��Ҟ�g�����8(j���Zd��Ѿ>�����pU�����x��	95�S�;f�3U���Ù��$�S_�5vWgsY��@�{�<��!���q�ە@��.��b,�}g�P�S��`˅��q$���ߧ�sg�Ns�c�m��̍��&۴פs3�dR׾ex�n�H(���B��A���K�[�Ρ�Q,�u*�sn��b��K�?	�҆����p���Qon_��� ��:h"�}�޻M��>#t:p6�z��YA݀��e�]G���SKW
��&�~B:���Fh̨c-����Ѻ+���ob.��xKDC��Q��Z��|���!)y���$K��lm
�q���?�|�y�=���n��SSԧچL7Ԋ�+���9db���3���E;�`l�z"��'m�mgJ��5����`�<���;�����"���<�a� �o�ܺ�1�����R#���O���nj�n���u�݀b	�%�n�\�2�0�E2B�0U*N"YdYA�Tê�.�q�5wvB��6nX�3�^,x��ű���]���+y�1O���6�:���{�=������5�D� ϥ7��U�.F�k[Y��A�>��%SS\�6�]^#b�B����AF�1?���Z4���[I�Qc^Pf�,)%�n��ɹ���s�N261p�{/�
���-�������֣��"f�|�6{�oB>=�cz$]���}\c�s��*Y����Y�\�	=�(�0>�E�[���,k��պ��w�����P|�lˇ��vQ�I���!1pr�L�� �Yl���v�	`0kQ=�ӵ��e��>	�x@�ձF��/�y�n�o�YsӸ!�[��f�fڔ��g���>L*��]Bel)�X�7�b�4�(�T��d��<w��e���n�')�o�\҂ʗH���j�@��j��$Q�[/G��$Al���<�𹜧e�_!���dSy(`V<m�1���h84ӻD�@ܷ伔g��"R�=qVn�[�<@W���I�rBe���w cS��RD��";;�R�hE�;�f{�������d��v(4��I $3 +I�����Y�e<�{GT�&��f���S˴��u)z8S��S�:�1U��Ι�~�C��Pʎǌ��$��a�s�&<E�'���ub���C� 
��r��hv�J��2�nP����ETNEȵ��F0����g���r����Xk�LBfc"�ʟ�c!�˙@���۷t
J�#�����a�
R��r������cs<��8P�PD�� ���}ٚ@�������ܩi�+p���L%��m�`���r�~�J���I��>c��>4���s<����,��7�����B�J��߇�`k��K�-4�q(�xu��n�¨�S�
/�;#����Ӗ(CbC\�����؝ɯ�P�%��N�gk����i�5������h�C�'��H��X����Y$mP$���=j83��9���2, %�ޮћ����|"s�hc��S��K��p���?x�u����oI�_�e	���Q^7�<�ݗ$���O��B���d1����F�O����eI��%�*b�Z/�?rŃې�[t_{$M���l�]�J9�!h�[о�b��c�y��tM䘯��HjI�W�xe�ʉse�#4bޙ��I�U޳
Ȁ��	O��j<%��o1����O�~~�:8���3��LӲt^K8��	@�#xH� _�ʕ.�y^��?�3���[_�¹Om��n�.�?���*炙��!VF��b/��-�p\3��u���I�7f!^!(0�h�!�߮�GA[�B_��)U4��e���i�
�K\��f�:�1���w!0eH�vBEx-&&2�.@�p"��Y�&��g��@�B޾l݃\��	�g�#���*���5�8�X��j%e��ו���U-9�Xmv�>��hfH�h����r�-V��50h ���9:�=�Kܥ9���C����Cg��Z/R1y��b��q����]�$�?[s����h�Q�#��P�_3׷���ĸ�7��g]=|�|Ћ�ê�X�E�Q��}�G�r��!H�]�< �ҟu=��=��f��
���_��t֟����ԫ� �V$�&����ۊ7���<7���W_O�'���0��Eb|�����4�a�
�`m�*�­x��Vȣ�KO�_N�H;|�_B��he���Q4���|�T ~��L>��VTbf�3k�����sBaI�윒�s��3�է�����M<[:��c�^U8pJ��� `����Ƃ� ]F�q�:���h���3��Y����~g�2z�^��@�	4w���f���X9(�!B����4��`�.��ͨ4�D����s����)�ƉEc=q�6;!��}[3l�K~D�a��h~���X;|f�`#���E�a/
��nP�x����/)�4�&���n� �P��N��1�M�ǻ�K5�K^���x[ �RͷY�6.�>dR�2��_�.�����*�x��"�rf5��X6���$�v�!r���_7`�+����[|�$���F>��7]��0�F��S/7��]x��m�ӟ��H|�@s��.���\��ro�,⺟w��ߺ�zX;{~���*���׼?�z�������؊��R�4�׃�_h�6��� �L�zh�s���q��Z`9�J�ʫ���6���z������T̏����uڦ5��u��]���Ϧ8f��'%�,� &��oϭF\���v�:��~�͵R�?�0�q��F�e�����c��g����G�|�#��e�XoP��R����Eq����,_�k�Q�K�?�6b����u^���U��p\��3�/�#��HW�W����Gw�:Ze�Z����׾P>K/|�3n�Z����)����>Z�_�*AV�Ԧ��	�j/0��0�Rn��ǫ2m/pU�O[��F�W����]폍��Na{�j�V�ӹ�*`1�������W�ۡ�:�P"G��8$h����%�q�����<P.!�$p<A��
YB3�$]k����I�o��x�q����d�^w�Y����*�]_7�c󦇫�DIV>�նٓ�9���3�1�NyY�����8��|&��d7g�'��aP~��~ۍ���"�Q9EF&��k��ި�֏�|0]����tf`�-�쉺�@A�gh+�'��!�*C}9k�T�	z��I�2mU^M]��,�#uA{
=��������R�1az�`01$͓���-��V��B��AI��P�
޲S���{�,{h��WW�p��/�]7�	[C�MD.�G= ���b>ڨ��S�`�D4C3���!�d<��%�1���@'GDy$`I��ܵ#X=��#i�'�z�7?� r4 91�ǫ�
�~^A@�]�bO�r�[U�f ep��9���p�'p�s�M��ծ�1�8��b:�]43?�g�t�$Xm!��)e4'�o���M�d�5�M��;RBg���95I�����FF�4�o4X��'{��m��\6Z�|��2΅V�7*׆Ӯ��赸_�:���bG�p�@��0�8�J^��o-�K�۹���q|�w9&	�ަ�K�a6��nŅ��c�+8��y�Z8��~�z�H��as:� #���+�4E�2f4݉&��|��P�+X���Me�a	�bB=����$Bmshɵ+Ewrs%G��~�M72[{����4P:�d�x�6�����i}�+����`�\�fS�*��d�n����[Ų�d�s�[��d�Px����m�uMفk�1mD�	�Y+����m�csZ���S�E<��%ݠe��U�V�H��2����_h}e����c�n{���AÝ�1�_l�ղ�$m�7��L���EԤ¬��_�n:y�=���vL������u��n,���0�y_�3���R,��3��tQ.q7<�+����	µO��z�Q�Q&�ǚPng���u64��TY����ҍ�­@����,;y��f̓��x�9�i�� ��e,u��{=��6lp�x�I�W�n��3{���gp���'�(t�P��Q�}V�2���P���'�C�eB)�w���{�d�������� ��CT8�D3H��"���XS0W��UjO$�� ��yr��v���@������(�x}X�>0m�2��W[}�݇P��
%_0�2-T'h4
rMɱb��s\���=���i�2��h̤�^�3�U�g+����c�dyr�B��CЮ��b�{���׵��9[M�+��R�<G9��©;�ҿ�
�Ř��ʬ�*(��,(�eS]�%i�dV��m{ٰ���B�?1Ԓ�h�Z<�8Î�~%���_D��{:ҿ���G@���%e3�6n�}n�~ܯoZ�P������Z�Ŕ�W7�n�Lw������}�C�8`��>�f^�~g�8�+L�|�"4}�+g�:{�?|����d�#�D>���^v�YY��,�x�G�nPR+���MPW�.u��JJ�����|��eϘ�/�E���6� 	7�~Ԅ|�*��=�d�=��>	�q���dfḴ�͒&� e�t����	�9d�	��|��j���7Ǥy�U=�BLD�������9��ռ�2/ri����+0`��i+����@�^bn�V׀��$���#�;TG��]��m�Ve�'UW�vp/-T�F����¦W��E���8gKҥQ)t����2��G"�q*_�J��>+R�=�/���*3��ȔR���*�����#����޲������a��ܪ1QT'w=�*Tiss	��S`�p N����eڢ��d�\�T[M�\MǬ����RG�~�vO�N��}����y h��h^��Y���*( pI�����Vo�ג��-����

��_䩤�6 �C}U@�:��"���Md9��zCz� !Ҥ��ʳ%��� ���;�@י��X�2=TrZ��GP����%a���v�������]�����P����9����%�p�x����)z��&Avi��;0�	��G�����8�$��>�x���7Y��	���'}y8���^�9_n+�:q'�7�8M�gz#m�-2G��I�0\�j%��F��"N�	:=�$�k�|3���Xtu�;�D��%-�"�v�,Z�,�sǉάH!�~�kټ�p���=lH�y��Bf��BC���Oi(K=��Ȫ�����f#����4�Hb:�r_&
�*�jmH��[G��^*J$�!���qQċ�G'��c�|�7��<1�U�֌l\�Ju�_��/I���/	/��_�
�W�7VW����k�2���쨩��#Ϙc~�F��Q扤\�b4M�>�0`��`�(!��`"�7��������g��'/�߇�H�������/�m@��m:,��5���g���7����.��F��ݻ5H��;>7��%�nY���m�hnY$��S
����1A9�]�!���ŧ�X����6�+����U���N  ��rK̗��3��&}3���HD�����c�Be���s��"���O��4��1�����M���w�Y��ڴ.�W��ɜJD�B��)�A&|)D;'��J�����-��-Wz
Sn���C�e'E�Z����G\�!X�g>��XjkV�*h��R��I �+lְ^H ��s�r�?����2��f�� w�	i��7��^���J��'y�d�|�H�E�g�Ey��k#)�-U$����`y뵹O�l���CkL������`p�Ӽ*��M]��".A��o�9��'^��H_<��L>!����Z��>.P2	,%qEw|ȷ�/�~�c�?��f��k�A����`z/i�<�y��g�[���ӛ�6�=��f�on긊�d��L��4�ox�NͻW�e(��*���0��]�L��0�k���Mh��F��]�QAK)����(@�_aɄ� O�
��������������0#:�æG���)��ڨt��:[�W��hʘ��zd�eC4��4�0��#88�FC���>�ԍ-$
��_)�Ξ' �LM��8��T�lKx��8�:�WR��{M�2[�n���	f��*U��C�U��U8�Dw�6G��~���P��R��yDb�F'���;�*Otc�|�����V*��M�P��p��e]&�5IQ.�lO瀈����b�)l�s'̤Q�q5�&�J���O�xo|��^�ȃݖu��5)�jG0�2��ig<�X�|F1S�6>Bm�m������}��.�hH=�"��qgZ������JNE�g�#v���'���r��yN+�M�3�	�X����.��D]J��X�]ϐ̦㙚@y�C��1��S�	@ǜ�� �#���27yC���BX���<��A`�1�P�e}41X�6�ŞnX<ֽG}<&L\�-��c��u��#.{�
Vf��g�;J>��q;�ELmV��4f�Y�HhN3"��N�>��\��>�k�^����P��(�L�P�b�� w˥a@����Hh]Ö�uy�)���{�p�X툕~�$_�A�$��Wo��6�:�a6����=й��9��[2�6��x�4��|~/mG�|�-\R{���5� .p�J�iG�=F&�濃c�n.Q��-Y��D�ST<#����slw*c���L$���F�#�!��;��<L�Ҳ���a%vn�o]J֨���h��:���5q��=�p(����wG��\!���}���ߖ���b�g�ͣ��� ґ�Ȧ]0^��W���F���)��k�=P��Mr��=�-�"p���m:Z+�FR�6l���' �ք"=˪<A�!aWڵkU�]��\�N��.��Ss��v��P��t{��>�38�h��S	d�:Ċ:t[�9ĎQ�o'7mZ�<��9߉v��zHI�:Ԥ���%��@Zw���>�����_����;O��'�4L�jJȣ�)�o$�lV���J�������:- 7���d�0B�f�:�9Dz(�	�7�d	q �cA 98`e�v�q>�>E���:y�@b9���"u�A��f=���.8U��N˦��w�N��������sbS�d_ Nď9��[��|����BE��᮹����;�G���Z_-`䓱�K��,��t�oԗ�E_n=K�l09�^�M���gy�CT �i���(;�ܘ����7����e+�`���	��o�����n�t�m�W�$Ţ\}�W�y~.&���̭�.%.�D_��D���b����ݺ�����mN<q�����q
p�l/b���c�9+��HD�3h��Ez����[Kϻ��Z�#���C;��l��ߋ�k�S�����h��=�N�_o���R��������;u$O����fw7y�S�V��Է��(GPrMJO?��U�۾���d���e��q��k*uu_�`-�N��%@�q�p��M��}�iP�Mf�1~s$�A�F��S;['q[�"�|����M�_eEV���u��-�{�����a�Ӱ2m��M���K%�D���űGN��ɱv?,+q����.�d�V�U4!�fe���)g`��mX-���/K�#�m�6�4#�7+iOz�� ����G%�:�)�ˈg��_�y��{���D��8��s�|L�a�I��ͬ�m}�l%��)S=�<������P9�:�\�4� ?yI���uS�����]��+JhPQ#��|�y]_�}�:Q�7
��MP�_ p�:$@��ĸZ�K�Ɣ��.�`p�7R֮$�e���o݂����bF�0~{��u(�mɒyu_��x�8�l�OV���:�M"��p�:��v�chT�ѴYO5�b�� fo﫡�ٖ{g�)����Ra>���o�+������GC1�֊O�o����{��唛��ŧE�6"��bäI�w?/ո���{�AFnx�)�t,�*�t
b��pP�E�g�to\t}�t���۳�!b������W>YPh�C�������Y̌��%@��o+��kQ��u��fQh����p_RC��|Y����S1����seI�D1?�J��z���h�o�T�a���<��+Oa���d7���[71��'�|~�E�0`��s���/�½�Qxe�d*,�z��d��4&\>��"�r���ͰZ�"sV,���H�L=�A�At,h�e�A�g 纋����@A~lS`��-�ԛ�25�\�C2G���h��s۴|�"瞨��~79��H�/���
g�
%��{��V���PG
��š��4�&͌�k���0N?��[0�pJ�AdDܨ�Bf/��*��IXXZ�_Uz�M_q#c�%YO������9�웤�>�f�//7j�	��P��!Fhc�E��
_��Q�v9��XYu��Ha���_���#��7��'��4�
X�?����ڇ�yrv�!�M��s��y7wN�Ͽ��2�{�u��׹��H�a^ڪi<tDݓgk������0��;���=J�i�Ȍ+�CK��,�+IQ�j���a{�|
<4�V���z�[-̀�NTҬ�gЌ�����N�ǰ��d��nf���Y\i{d��r�W�j���RTm4}�;�W�h���_;��κҫ�H�]JQ�,�h�	��=e+IU�t�����XB���(����]GF�0��f�?����Z��̼{-�8z���f�EqQ0�P*����2xM^pe�h鎊��B2��2�jx�¼'�m��T�t%���q쀓*a��e0x�vm�p��]u�U���T�j�#��W����|���"��^zW��f�	��E�� �#׋Y�G�'S�.�zFuX��;�R�hÛ�X�U�;�3S��yC�9�Hv����8��|�U��q_�W*��q'�6�b;����I��a�E�o����v��w�7r���N�ngz�5���)+O��H�|�EX�`
Qz@��� �f�>>{a���S��+bD�WR}�h�_��&ҕ�2\!@�]��i����E��(wE��oȎ�-�{���+���뷀�]kJ?�/�ih��E&t��Dz��;0����o�P)�y6Ɉ�9A�
�� �?���B��UV��,֎1C�W���W�SL;�4Q�2��y�z	)�#K`aC�H� `�'եk�.a�f1��q�g�9��S	ᴙ�w�D����ȉ�S�#��Cn�f�E]�Q؍��M
�����o]����Q0�&���`�L9�$�cө��n����j�Kp�\�s?���0t��a�n1?Z��\_A�� ���F�O263�	b%�}=7��*S�ѻ�e.^�"��fe�H>�����J��	���I��)v	��Q}��揯���R����;O��l������ӣ�{\E62$��j�|D��*>i�Pp����ۉE�c`-䵯u��@�}�O�M�dF`�O}�I0���cL���8��y��6�P�J:}��L�c�W�[+�[^�y~�X祡����^�<P�悕��{)J��G!��
�i�A�TQa�D��C�!�eJ�{Lx�<�ԅ�@x0��3�za���*x���|B��M s�i��z�������,@����#�Pz[/&��������&P!m�/��Īlg���5����7X�������>p� �=���~5�O�Ҡ��~���P%�
VÚ���q,vU���
_�ݙ�9�����+��8]�R�X�1d������f{&����5V����Iй~+�)�W�_0�[�P6�S�ӿ�.�-�]Y)�� ��y_�O�絥�U����l�*o�gJQ�yMS��?�uT��f�DgrKs���ӢK��yA�C ������?v���Y�L��k����8���7��l���Ψ3���z��H�xj�-�V$%b<�``�	?|w|���p�v���+t�25�`zZO��3����ͅ�ܫܶ��L�d���W5:~pu�j�ј�Hb��)�0��<p��D��p��ק�,���'��T�G�]��J�t�5�P�YV��Q@�u�$״�@�%0�ؕ��)�%�~��ӿ&gRl��֬R��ŉM�]���Wn|�`9��#P�!-��I��S�_V�N!I%�'��,�(���N7㨛t�mt�b��a�7��aP$'W��[Gv�r8����j����/���{�7bj�����]�W��u06A+U
��
�V��׹VL��k��x,ۥF�NhY�q�-':E�5۠k{4��!P�y�z8���y�w�m��u;�qa��r>�l�h1/��
��[#g�=����� ��~�51��î�j��Յ��Lp��B�'�/:���8�&�Y���^�[��=���+��q�F�ٕwG����o�2��E��P1�A��'���Y��[��@�R���de���c$����6�v�GY�-;���?�z���a]���'��d�L���?��?������<1�G���t1�k�4�a7�c����+�"�T��Z*$�.��bqY$C��8}�T����|��ҙ��;�ƮFO�v�����r�-/���Z��Z�Y5�Ŏe�r���W">r���$�?���)��Ѐ�*� �"Vz�&�Vh��6?�bM�D�)d��y|��������Pj�h���s���}�����j��-�{��O/10_�M��e-r#��_݈*�E.��Q�f�r�f�Q�MT?F����K[�l�jW�D�	+�'�RHW�SB���f�7g�
�E�:�\��k|`7�+�stR�A�*��ַ;B�U~����_�R�3�l̆2e�@q��L����Gc�_��|n�I�\k2�b�E�����d|���NR����ރ	u�w���!���xۃ[eu�E1��v��q�D��p��:Y�	������fr�S$�ڼJV��ѻl��&��w���wóO@,�a��3ζJ���a	?�*w��%�J�#|��Z)�	O^�0��C���W7dd3Y�Bߘ���i�Q*.�_G�5=Th�0�eK{UL]�G�p�:`,�׈"!U��^��ە�]����Q��R!~�����?L��R���2z�!!�����7�ǉb��K� ��R�J2c���懪��6-��C���!�+_�WAK��k,�NY�\�"��0� ��}Y��� V��9�c#L|����?����WJ�"�@E������AP���>�S��*�t�(F�������J�eFS��e���8��ُ!���Hm\�4��Fs)�cc��H\�qkDR��r��4w���;�Ɗ{Sn�]�ө��S��Y���VS�����M�H݂X�*�^V�m�h����:�u��<TD[<�%�,�Q��@��\a�<_d����]g�1�2�lH����'����m��,_l�T
�)GWh�i��������9��1OdRB��T%-�p�������/3�l���{��"4��wp ��0�뼚x�:�J��rep~+KΝS7��
��$)��t£.E��2����F���3�nB9�rW�.l8Af,�oB��i�v��vV�������9]4��F[0ь5�1+Z�1z#���	rP ƨ��lz�?Q,a�iOϴY3��Lct�K���ׂ�	�CR�Ux�{��a(=!�*��K)fM�
�G�F�L�^�J�]��+�b�r �ӋY+��=�u�m/��^�V��=J�sו�+@��b�I�;��㞎 ��Ј�����#�No�V4xӠnY��$3}h	��p�y��zo�����
�j�~)O�-<�DZ�yG��cл��R��,^�{l77}��Id"�?�1�E�k!U��~�����8�'@�'�޶����}�։��\`��oG�� ��bI{1�b^��y�� ]5�?�?o;��e�vy/�����Kƣ�b�Y�R_`7{�R�P�{��	�ߝO�P��#��:இ���B�Qm�Ck��y�CFt��.�ԗ���2s�ʏi��(]��&�Z'�&����{;�_V�Ʉ�����8�@���5�'���0Ç�B��.�����|�����.���WNrHPi��lU:�p�~B/C�/�����t�y�y��V����͊�����*b��R�>,*�}��^h����8�3c�7U�hj�/��}ȾH��k��g�b��#]S6g��
�R:�����
�K�i��P��X�
+Nߤ��Q�DhI�t�w��c��HΔP�t��۹�ց �M����[�|i뜨FDޜ㴡�h����9���VLšB$`q�|�-��z�x.<W������L1q�-��ܮC���J4��k�S6l:\�a!8���ޤ)���g�Ʀ��_�[D=���nb��罵؆|�`Q���zg��F(=y�g�m���@�	�G��C4�;䪘}�Ij�n���[���
:ՄQcܿ�Oj)3@�@��\��F��qv랶��AȈ��5�����e��!U�*YI'�N���0̀id^�l[S�l�zpj/p�#0,��َ��*J<=��c��BI�iAS�1*g�*����!rOB�67w��-�\�����QY��L�Q�	D�p�e��M?���Cs���9���
�]m�Y4[��MDIln���z����a���V6�����?sʶ��s p�Q��� ��Z�8[�g�*.֊�n�R���#s��jc񀗞���bX�K&��$\�����Ռ�6��m�L��I��y�B�I���b�W�^}���
���o�����(�쇼&݅��Fy�e�K�٦a�&.!�f�����ʜ}�x�ߞw!��B��f��;m��2��n�Z�%*��{gv	���ݨwv��%�Q.ά�O�Un��c�ڹ��kDB�y��E�Z>�B�1Kd�|�o�^��K�����s��j~��U����H����������1HX:<��R#���E9`J]��׽�C���&����gJF#u���U"�I�֋��!�������.�z��=OG=u��0��2dn�M�1w��/F�q�H����;c��3ɽ�^�*�_����	���*��,N���&ꆬ��}j�Q)�"B�9�쟅0�������`r�_�:<�F�<f�9'u�1�G����I��B`6
BE�CM�K���:q��&f��9Fc��,��t$�sN@�G�p��WG4%m��F
���
@B�p�����V1��D�a)�o����.�3޷RӖ(���ϩ��j��8��Qk�I��NTE������m?_�w��ٿ��>��'��P�^�H�':3ݯ&��,ٹB�̶6��{&�>����ރpql���ƻך���ƌL��[�ܷ�$i�7b�.��<�	?�|ξ����h'�>/��w��+<D�D�5W�k"��9E�	�r弮���Us.��)x�o���T&P7�����/P�;����Җ0�G��c�z	� zWȁ�[����I��Yl3�j�Fq�񪌭�"O���
`�������v��CO�`�!�|������;��I�FV:���_��PR��?���s�Z��$��F��GV'��������T��w���\mK� �tH�I����OKui�G���x���NѦAn+�^��q���g2���V��"r{�ȑ&�H���o#,'��yu!�RԚ�e盇AJ�`�����t�ԁC�2L4�t�@6r��/��W���%���j�S��M�4��5��Pq�a��|�`��~�M��4Wm��!��N�:�#��o�Eu'��׏�h�C�@���9��F��)?��[� �lVM��m8!�����e���V�oa5���t����q�*%� ��O�dub���X��T����yk���iYcX,�˛18�N�� ~��^�ڮ3�ɖ����#�TG���R�p5����d��	!�q%u��v��y�p0�4�ȅ$�j�x��v<��>��t�����"�����{~����{���c-��(Ճ�n�P���`�5�fD��F �Ga9�JH�G���6�il�H�6�9~ǒ��Z�����Wzlf{�)Q��+��J����E%��O�qX�js�p~���"Ö�Y�	�wR�{m�ɮɻ��>$�Z�$N��O��ѓ�O� %1��u$�#�S#w}�EU�����Y�oel9rW���L٬���`��-c���'/�X�����D�t�)L1�I��� ����_��0�yDD��z��H��lS+�G,!�Dk�`.#��[�Ipd������"~����lȃ�B�h�%�!���ߛjT��e'��Rj����x�2QZ�n��2���(�2MOk�&,���w6�vG���B.����v� ��UP�e��&�ߘ�!�3/���4���߾���#jGg��}�_$=��A��_�N�5tW�}8yqN�m�3�s&���<h
#6�<�5hy���'G���z �$Z�j�����YYP�&�G��:�5�������%�%_�c�^��O_M��%i�)�8��]�Q�v�i#�rp��l�u{н�u���7GC�jbr�@�|ωeS�b�Nn$��H*l�0�Rkc�N�1�\�_�GW������Īy��_@C���)��u�o����6���K���T�蓿?A�v�e�u cU�g{���I�󎟐T�/Ͱ�죿��saW.ӓ㸚�a'���8AJ��� ��5�=�G��MLhCM�lJ�}��4��էkzl�wSKo�I���_�,��?�v��T�
Y>2��O�4,���� S�J""xg��׹�\�Ja�J*����B�1"��U�s0�Ľ�$؀3*�е�0���g]�F)Ҷ������:�������;)�_|a��?�|hIp�j@VN�7j�e/��4���	����#B�O��o��S2�&
����&�� ���|�A����k��S��w����ʶ!>Gz�����ոjv�d?��'N�W2|'D�׶��ԵX�L�bs�r+������D�#\���+\��T���r�Qܸ�$u^���/ӕ�Ŗ`v,��쇃�5�!Đp�Lpзak�[��+���y[�����٫��=��kO9�0,{;�4���˞�|���?p)�dTo������-S��b���T��3I�,$9�p� �����l��,�%����摿(�CCLĻ���'���dG!]�>�.8�{8%KhQ�S���ȟ���j\,�5ￏT>cg#�򍸒b�a���O�8�	N�N䞢�VS��"�;GK������N�Ǹ��k�0(���ʊ���"���U���|�0�QG(2�_�zL�7Խ".`g=�\���NkeC��k5K2++�Ec��Ks����Z��Dne������m�R�e�yȒ�cN|�2Ä*���RN��� w�K�P.����*q��C���[�pp�}�����վ���ާ������UC��0�R[1S����
e�[�@/���$pŻ��4d��I��":. M�˚�zY���gRM�5�����_�6ޅk����r���ߏ��b�i��R���7Uaf�	��mI7�3��%�+>�7/�����Iߗ0��NP�?h/D�ֻ�e@���YW�>Q4���n2�B�0z�]���1����{�����eW�ߋ�g�����]�e�2y�?�Wẽ՗o����\�A�<�n��[���
<f9�)�xҎ�>F�O>I�c-�3ޢ�%t�͈�ID(j����6��f���dZFz-K���c�������y�j�Z������@_�72�r��C$i�Nw	�8��
���F}:� ��z���(��R�:�}R}�Em��W�p[ 덪�	D\5%(�<�Ս�_��x��o%�EId���`�l�"=�5Xrm�Ŭu��M|~&��e�'Җ6���w۾�FG�lR qA�X;dj����O�V4�Z����;@����Ȯ2g`��{g�/�~5���}���L1��bي�^��4ӯM큺�I�LR�Bs6N���Dw��d[�};YxSy���SeP�2z��="
�j�u�2��C��ͫ�.��KlQ����9�m�ĄPw��6(7g*L�R�P��P��lT^�L6�W�mw�da����N�^��z2��� �)�8`�
�k�ȁ2�)'���c=�͛8��BG�ȴ�q�i�~���f�D)��s����	x[-;�FRW��R[��͆!�tk-g��uއ��,@pH�Ъ8���VU�=�1fN��*@�2!�M�6tߒm���<��K8=X�h�3?��w����ʡΛ�y��������� �/�ɠ˲`���{QHf�Þ�_A�GITt��lg'r�Q������@��	�	G0�=�E���;FV��F�z5�f����ϴj�f\�%�S�(�$Dg�S�Ah�����>O��ȇ��*cH�xZ�`��SO(A�z�U;���.�RT���`O��T+�V�K��x3���Nv~�͝�G���D���b;+��ɧ�I���%�kt���6�95���t�/���5�[�ٕZ.k����B���Y���N��y�<���6�F��N��Ӟ#�*h2)�9�����2M�a��c��n/�� j͝V��7�0j���\k���̢h�Z3�4�;G;l�k�pR�o�*1)o�ZfpA>�葈U�N�	�`K�Y��@�c,ڱɳw�T{�)r�]�W)��'m�J�ނ�I!���A�L�d�]��?��7]�4�!E�е��M���2\3,��KV�x�t�!{]�/��v��N��T��ǘ��/(�vpY�w�
��U�[�cNx��	*���N���4�tJO��)��2�E�[B�d��s�E�F� �Bk�Q�d.b���即��,Q�%�0��Ë*Y"Ր�R�zSR�E���M�^�j�n0�F��>^�M -ALp�e�{�2��0�5/b�Yo�0����/~PJ��PG�G���`S`�L�J:��yr��
^ݡ��yoīzB��/�˙�ŞvT�TA�mn(İ�k?;^T�|��&��SA.�&Ҏ�RrV���Ω�/�,��8���@�o�ͿB�u>l��#W��ϰߥ��F"�	d;h��J�b$un�/��Y�˚�K�ҭԎ2�Ś���G0n�m΋W�N�"�J�gP���]�bp/5i�/��Ny�m]�]�����v#��{dT���)��Bۮ��4i2�������:tO��x x��~F��'�L��h�8:���>?�����5L�� >3�C3*�\�-��l��q��ՀK��!J$����?�o�ڲ��$Gp )Aŗ��o�K�MYT ܃��{k2BMy Q5�֭X���kHL�A�6/Io=�f�O&������0�Ok�g����#Qql�\�<'{(������~P ؉F���N��^��"�҉��k��y��ǐD0� ],쵏�Lt^�G䪟K�"��w掷|%l�BG:�ܝ�#��LU�"�� \��zKC)��H�P������n��{J���A�-�z���}f���m�i}��_A��r�?�a�!q@�[����A��͕r]�"�i�Mqѻ�y���ME�]7zp�[��5�k�E�ߝ���;�=��9RV�A�)��Ek*��	dl���*������m����I[�8�mЍ3ǧ@�4`�����g�d�Q��� �����TtO�0���F���*b�\�b���I�%�f�6-3l�+�E�Ax��/ot�+�l��@�����$�~w�u�ڟ�Fs�����k�[�ϵ�B��6�� ?Y
,0�q��;�1C�d)(L�aX��wiaEC[�(��M�D���W2a4�������&��Y����QW�}��K��`��@��ѲF�������V��[�`���4�������w��i:O|�3#pv�X�|2�B���
��B#��E����a�iC]vxr��}`+��Bz:�_oZ�d�d�|���Jd,��Tc��!#�n�°ڊ�����ӰBMLc��v[Cz"U'`|\�H�ؖ�J�iW�VH��ӈ./
���u�����>8T�K��
�Q=~[4#���j��`�s��ƿ78<sL�������0ܓ�\p_#ؗ|��w�VM?�M�����Nv1E2w��ܱ�|SWPLl�﨣h� O����Hw2��L��L$1�A�����*mW�	^7�|t��&�Ă#{��|[�H�S
Z\/Nɝ.�2��:�jˡ�,��� ,r� x�)�L�U\|�����}�Uވ5w�7�;��g����~���(Z��m�B�,�)ɖ�%S�9��q9�k��h�V�x|"�n�h�_�z���wg�ý�@{)��@�$Q����x�����m�8(��H@>x�4m<�
�Ki���"��������-rg�*�oKF+=;�R�ؗ��� ͮ���}�"��4�R����<�}c�c�؀���.Ra�Ǆ�sp��aK9�� m$ &ѣc��])	\QP�a��#������x�ީ�@�=T�A@��!_�������$L��f�!��:Y��(���+����tɓ�M<>�+�M�;���ys�?S	��+�Gf��7�1o���2/ʷ~���f��S\f���]��'�=��"���'U��f!���>bљ
��D�X��
����C��S�;Y�
���N�ȥcR;�l�n6��b�wԴ�>q8"�߄�.Y�QH�F�u8݉mo�����k�����/���?D<}k3&����M�z>�U(ɬ�9�jD�?�G�z#x(�^�������Yr<�����j�bK�S����@u�F��'�%%n�"4	*@٫�P�XPM�yM�J�9ͭ��ƢG�'�]͆G^�d\*7>�EQ����Ӆ���ӋȮӊ_�֙oo2m����3f�ZK���Y�=�l����ɯ�ʞՖ/ۻ�I�}epU(E�X��������[\̓�����AԾM�o�^M��P�����,,~�����������|_P]��RD���>*If��cG�Ꮦ8���ۅ��(�X��oփ�|�Z��Og�M�ت�a�sWB��>�U��xRj:) 9�<��@j:z�F�K�I�!3ʝJw�e9\�_"kh�P���3:�I�S����܅����(e_BD���n�f�"�LS�F�Dq�19*�FK�wO�F��o�n�$	ی$�:ݠ�+�B�GH)ˡ�zq[v��9HKŶ>�{��
�|�$�"�dj��dOC&W"j����N�08����-�}o��9bVE� �����,w��&ٸ��2�ꞙ7 ��d�T�� �eJ����'v ~�l��l��Z���h�v!Z6�Ɏ̩�\`�3���3ؿ���,�3����{�Jzwٽ���+�:�ǋ�/;�md ����gkW;�|��*�3�S�S"��!��v��k�˞,�g�`��-���3p�����!�qp���H�`R��.�`�A�Y��I���7:�ι�V��e��ݞ
_�d݋Q;rA띶p�&�� �E����6(��>��C��c�:ErS��f)�`Kp�{�l�3�ךd���܆Wz\,z���m�41XX��1�>���k�-M��� �H�0�R�?\6�ea �<,J:!����9MiҔ�މV�1K�,���oȄV�x^��E=�PaR�2��f��;�r��-�y>U�N�$N�w�	������D�)�J(�bbKlx��вD���]=�y�����ލ5i�>u���j��XerM�h'�تw<)o�L�C\7V��W�N�:`��9P#���V���)uh߳�S���=�C��$H��PݣwSO�ag���%�>f�-lBIL���7�Vy��m�V��9��;���m?���|��ҵ#:�t�h�x��xB_��koǉ��?�!1		`g/�x�5j�!�x�9r�:���{v�>z�	FX n����t���Q���@!*��}g\��>8le��/¡�0��������+%��V�  �Z��Q|�`����R� Z���nL�?�.Nw�'�-u�l��;r�Y�9�H�@����%vx�F��mX =@%p�b�5�OM�?���K����/lV�lra&_�\��g� pi��"�I�VW����4E�Lj�m�����^}T�Ͼ�v��Z/!cG�GZhK��ᡊ�u�����sU��� ����S9�%���.q�r�;��;0v��| ��#�Du��\f�n�1�Z�
�n��x&^�]�Vm?���~��4�j�HV;�̭��J�A��¤,L쨬p�ʅ�)��(�9%�\��'I�E	㶻�T���+�_y����𚰿n�h�)^m�L`p�WĐ�쨬>zI�7�9ݖ���y�i�R)��A"��bl����u��C��^���0�E��(O��+�LUe�w��vRY�3�W�pf�zb�ܜVَ�s:���K;H��݊LF�	�⇐;u
��������I��*�F/���\���F���UY7�1�9is	���w#I܇��T�V�d�X��� ]2�mv�^��eiV�Z�x�f���N�j(Y��#�%�&{ԘrX�'L�b&ȴ��MI!-ڂ��E�sp��c���Љ�q(�@b��J_�u��^aQݡ��ZBz�V���ztq����8,�G��@[<Uq�bC�{��3�;�B��}Z�ސ��	�uƋ����n�VQQ_�\�n�K��O����a��2�v>6��J]�5Z���pcWH��^����9Yz��[w^eU����� G!g����ʏ�Sk�+9�V���L�)�� ￪��x#��*pm�\���� �������J�Dʅ��a$P.���E�������.��!�:RN��LBY��<4m`��v�?�%�K�bIL�[�ߡ8n�z�Ɇ	��$�y�?Q)�?�/�dO^�c��0�-��:��}��M:�`�r8�P.��"�_�(8�����e��e^/�T�~�y^C#�?ύ�*�n���Z�,�}�r0�X<J|��P�K���Lԓ��p$ݞ?@l�R\$���8 �����?����Ӊd�_[�0��}�T�`���Z�۶0�������ь��'�	�7�DZ����i� ;S�7z�r㊀^�Mɟ�Ỳ^�\�ȗ��M�7�L|u]`�@��o`��2զ�4a�q�������	��i�g���4-ٿ�<��d�Y忨zYEi +�E�_�rA���t1tEU�E}�"�3���ߞU����j5�Lf���=kxD��!�0�ۊE��BY�1���[nz}ҢQ�I|��7�Վm�h*MPB{�ݑz�&, |��O�f�����Gb�.����C�a�8���7�m})��,2���Z#����)'Ux�p���pPɢ�%2*/3f�e�r������0��U:Q�F�T�?P�%št�Ѻ��C��(��)������I#�T�����Δ@A��d~�$��
7�tՉp�؇�&�|pn�6�q�����K/�=GDa�qk�����Y��[ݬ�e�X���Q��X�96����U�n���da疞Σb�p��`�b�W�N��QѺ5�zW�&�'B��P����V[�� �D7@y���/��̤�>�QR��`���0M���(cc�#.�*�ms2�p���^�e'!��[� w����	}F��A��}@|tΎ�(ou�YR˝B1�j���Ձ��>ۍ�QiKwzpb
m��A˝�����kb�@h�gw��*�Uh�){����0A��^�N�P�,`��0�����i]6W#+��H�Cw�s�\�|#��Ѳ-������Q�|"FhXV���v7��f����5N��ٚq� ެ�4�M^c�.W��v�0�Je
�����[>33K���L����y�$�T�2�GAn,��Ƣ����V�( A���A��F�d���8(�"e� ps��q�J���]�I��2�uK�C{���D=�Ո�ܱ�K]�y�E@�v���勜w[���`y�Q��6��ȬXpU����6Gɝ�@��,ɐ^���� 98Ym�V ,�+�"'�����C=�7��P�Z!�U�r���.`��Ǟ2���E�������j�/�]��I��h��A��6e̜�e�ߢ��6���9��v�A:;^h�-�3%D��U�Q�@C$e�jK��q�x�38�`���<�������2�4��֋C�J�@��k���![��:�*aoB�[?��8� 9�}�	�P�$���M0��1
R�9k�c�o\J��p)�9y��G�:��8V�� �����j�
-����1:S�K��$��a�L�	�7c3c�Z�&#7?��7�Gxs������i��}�\;,e���~��>���o� %^���)�V�!��_�;#�5y�(�8ǅ���&A��ro�����Dw:  \�>�@N-���U�Bd�y��
�|o���/�oJ���y"��e0`����v(R�]�K��X��T��G>�0�Τ�:��޷5��:Hא�r����A}eY~�+�z�^���	�Lj�PܘO��18Kf]ݴW��|���y�>�j� ���V���6KA������B������lp;���.����1�<�a	/��a<�@c��k�-�y.XKԙ�Z�5�@tSW$z#�:�K��b�O��X�Zl2T�Ἶ��3��R�q���o;�?���CE�@�.��|��~�*�*>�a��^�s<)J�{��2�0�(��[v�\��V�"+ϟpŏ�t
�˃���S	WC90���f��:�m��ۢ��,8.����Z���i������;�o(�.A�W`��k�d<�ϊ�FF�JG[��%��yR�����:;+U'i�1���c�@}�����7�&Vc��݀�x̋-s����K�Mx�U{x������+=2e�8�d}�*T�y��4��QD1C��h��I��dp��5����18̾=C����ܒ�Bst�9�����m�qh��cDL���:��/���~�Dæ�����+p��b�2��#��gV.�+�:^\v���DJd�+�@���>nקi�騿�0WӒ�[�$�:[�:� ~x��MSԁ�u��f��L��'��u��kp٣�4�6��4=-5�Q�� �Cu4����A�t���1��k��\��x������$n`���ѭ0���S����3���p�G.Y�*[�,<-�R���ٳ;��ח�O�k��_6Fu�O�.�6	���l�
aNP$���	��??/J^��Q=@{E�C�ɕ?�$6��$�T��Id�MJ��qut�<�L����;!�1�V.ɄD�l���&��v�%p��찲�Z��س(kv�D���t?���/��f��hij'9�U=���_����C����<���nk� �c�5*K��Q��n?��B�I��F��P�ec���-���Ѡ���ˊ�d[&t��\s�a��4X
z,}�2�/5�9pX���"Pfi&�ڞ�ۮmr��`+���'�ʀ��a�$��C��`p�l{�&hi�fk�� ��\�
V��|#�D������L*�K=�ԥMg8�����p>0�A:��ah���G�Bϗ���f##�ޯ����s��CDw�8�����J�S�N��Q��jtC�5�t��(������}����w���8�OӰh�`&��Mp[G�.o�}gx�,7���)��{9Uw��X�Xrx�Sev� K��|��&	�����7�[q���s8��a��TID���D�7yl'iNH ��.�_ɠ�؉��U�X
�d/=E�B7v�,�Z9d} [���@��|��=�$��YD9÷ǒ��B�������;���G�[b�ER�t�B�.]6U��qUL�X^u�4�F���!x��i�%�D�!�0>�i⒚��T5�<#5����E
k͖z�rp��X�Ot㡯��1��*ޟh��;���p&FpU3c�
��l-Y�T����9�F�tp}.Y��J�񺴟�����\e��3�=� �@��Lv:����=���R��oKv�A�W�N�8S�� &�/P�B���VeCl�ֈ��	����;�^ÑG�AHds�T?��63���֦w��b�?�<�h��+�����I^���7`����3��1/a�I���B�9K�vS��c����3�h����N.��̣���.�ˤM o�[͛���	�����`IkOI�b#�~��B��A��ݏ,WM�x�V��JG��9�
�Ԃ/!�o#_}�aך8�����%�ĽOO��+ZPwU�o���� Ƽ.GH^GpcS�Bf\e�K�&~z�↘��NuN)t@s�
�������.m��=�)�<�{�����JW-�⺀?[�RmO�0/�rL5�V9�k\�e���gs��F���!�۹T����~�oUv��4-�i�v�L�&%*:4ƐS�81��R��kZ�'�~ -�13q\��`~�5�0����жC��������'���d�U��U 
6xlb>�bgZR��s�J�I׹��&��~��-W��q1��6�
R����9�b�$�z��	��C�]���j7jg9���^�s���Q2�.��U���f�}��	Q�k�	
4���h�6M�n{�U���y�A2���7`�?=�hm&�5�z��UJJW�\���D�_�9 �}� Q��w_(�(��	���`���3���P�
T��pY
�Z�C�ӌ�j:[�-00���(�׀o�K�l$L�t_��{Cc����H�ژ�6rf)%Q%QY�����pv��Ԥ�<�}f�'�?YZPX�/y`6����k��b��-�z�͐��t�"?�����y�9�5�PU!�g��~�ћ(1��k�k���OȨ��].޼X�˫K@t�Ğ��@�y��k����qgVܺ����5��Tb:H+������Iȶ��2^�n00�5�a��n��u���Vـ�`��BK�^)a��.�t�	��V�yM��C�4�~�Ʉe�T=^{c�-�|&A��,��k[b��F�4U��Z>����P?Ľ�b����]gB>��x̜��p��0<�	E�\�Od��Q��ٚ��9��u�;Ѯs�A[�2Gs)x7�S��ʬ���PKh�>x�W��CI�0��0e��i�#�"ᛐ�+Bp‵�(�8�����iI������Vl�4P�_H����L�u�&�y}���VA����K�6�M��Q�I��>y�	+��9	�Z#���٣yh�v�z�Y��񁷳�t�p�+V���;�S���Tn��8&Jx����d�0����
#�l�eJ�P#3�(���	gz�|�9bki�x*�/�x�ɀ� �������ۢJkF���Ν�7�E�y%C�n]���d��Vq=�����Z��կ�����oy=	!|������<�j���y%ϒ��~�^8��b��as	�:�6��]qd."�V3,W��>PS��o�~��U6���Ԟ���rz�[5��W��!�,���qj�������s	�%YtL�y�>j�x�D3��,�3
й��dȽ�L��� � �/�7Bɍ�'���1����V�s��.2�}_TS�AЛ8����Gn��~��4պx5үe}��[���٨#�P����@6wü��P�Q��!��Y�Ƈ��q����H�#�K(K�
7^���~�ٴ�SKƫF�,�M�ďv��ny��1�y��VN��3h�esg��B͝���~����:{d��M��fJ�te�ϫ���,gV�8WӍ(?�Gx������s�J0G4��&�C*��BLJ�z�<�=�1���9ګ��ԏM����%�W�.���TC���|�?�VJ�N�p��iac˂0�j�<e����{�3������İ�Ʃ�����o�%F�O�=�g���PA�۾�0Q��ӑ�[1�ƛ�~W}TddѴ��'O����8�˩g˓U3�CL�l�%ZF�,	��+/����ѡd!��xS�u͇W���??��5	3�&�և�fk�ӂ��X-��hܿ�G�9G�Z��\�Y����a=&��#���5)��]/AEK�V�G���Hj��{��!�%i���0�K�MO��3��׵>!�)�]�]p��9g0�!�@K��a�=+��(��}�%p��"#��؀H�t\���Hz�����d�=�R����aʚI�ٌ��uR�Tץگ^
\���Cq��9;��2�ed��hT��8��QQ�ρ��C�B��7��m�[��;Oc.� �����Y���f�Dv�6��V����ݢ��<�U��#ԶpU�Y�ͼ��L�xb���Ѥ��G6X�+��Wԭ���	<� �WU�ֽ�X�����2��d����ܿ������L%�!_btml3���E�KU&�h�ƽA I2��!��h&���tp�mK"�:l2�)IR`����x
pl�K��ͨ�E%�䄹�����Q��e]����@����L�{���B��(�P�}
@�T蜋�YG�P�^�~� ��C�"�� �P�S��V��X�� �Yɫ��z�u�]��`������e2����g�q��%�v����V�S��5 �=5V��3�Gy~dJ���C�ZpbY�J9��(t������}�S˔(!˪�F�uh����6v3����wwA���J�,{�nؿmr�+��%:�����]�v�P--іo���Ce�c����u�M,6��q$���u2>!G�u�kf��z*J�d�6B�9_s~_�"Ӕ���N�@V��>���E��?j�NS_qx��+�2�������������%�W�SP� ����&X��	(�����qe5ܡ���#�g�-4�('~d�O����۪���
���N`�?mv"����'��F:�I< ���p��բl!���N�_R�9�D
��Cw�Ȭ���g@�/�d�-&�xD�i2[�mo��m,w.)O8�"����I-�����F!oi��i����^m9��^>���B;�k�h �H���to+m.s�1.Zٵ9�th����fe{�ݎ��4� $s�0rm��J�|aE2���-65�"�S|��KAA�WN7�i�jq�D�ՙ[з�G_��[����)��u���A>tJ�Ň�G�J�V
�,�����09C��hC�i��,����v<�,1)h�	�ڀ�3x]V��hj�i?���Xo=E��u��24Xz�{\�~��ێs"!����vh�C����g6��~�8�P�$���P� ͡G� ��fh�6,N�����5V�9�9��A��N�m�Q����Qb��d��v~8����\ί����T���^�P�(d�B3��J�8�%O^a�����?\j/������w����Z��ǫ`� ������=)k:�Z�$%� �=�����,g[Y��9qgKe @�'aY��{9�c�ӛ��Hm�Xt�x���bK`@�r]C*#<9r;�����4"����f,L���9?<٦�/�$$��,B�|�z���;�����"QP|��c�S4'3�,%�IQ�]�wF�Fg���A�C(��c�W+aA���(b�����w�Ly��kj�V�,q��]Nֈ���7]�����~�	�n�)��/\���\��RKz��@�SyEZ9���U�_8ߤ#�]?����T��Xx"�m��r4өj�^�X����3Nc�F��`B՜S+��,������p���~ "�Rx�ֳ�j� EH�v�;Z�lӟ�)�&�*��E�� w8i��eR�E�&"����4{eé3�������"�@\H��NC3��������p��.���P4j{K�K*y�.��d��d&���.��@�U��7��N�}��F���l���n-'�q�6}}�C������K������F2�ߒ�"��ޑ�9HKk_��
�U>W#�{ˠH�>-<��ςu#N
F���D���1����TT�:e�?	��ΰu�@3�GC+^HI���	�t%����PWT�}l>��^����YѴ����A�UU�6H͹hz4�!Bㅢh ���ӽ9��4+ޮ��2"V�FN��A���B�oD��95FLvY���@�lO�G�P�����
]�f�O{��d���`f`�=�`��R���g0+|�9/�g���j��$޵BJ(+�ȅ�5w�F	d��ґ��?jY�;� ͵_l^��MWn\�̠ƓP�l�-YZ�K�st-�áP}���T{��8ps�P�#YJ������*i5�0ɫՕ��|�R�lǅP	�a���X�_zv�E�P\�z�ɲX����Qq�NW�g�f���k�ēHvWY~P6�N�	M����D����L�#mP����m��6�q�UT��n��'~a����
�P �F@�U;�\o���G�<p���b\�"
�Z��J�b�����Ԓ	�B��������jC�]@�s���^�k�	���њ"\�μ+#���5Q+��)~���A�GB�F�����P#lotW�
�R����O�H �[�8N6	�~((3��8�����B|�� L������G?��TF`�r�3t[ֻè�M`����
|<��ʜ�Ƃ���}n�^�
�����/K�7����ը��F�
F��<*��C.�Ss`ѷ?Nk(�~��]��fb�_�{��ىdѶ�H�~��
V�� VS�H�(-�r؈'�����_C���D�@-��)ǗA%Cz���D��l?ص����F�s�B�����k�5Sy~v��&�뤭�0��X���v�'�_(�ڠ1���"mNW��sz��Ӝ\��s+i`��mN��b����S��Z���<.�~�����s���#�X�a��Ԛ�J�o[�Y�`����P���'ڶ�j��������y���u�=�X4�b*�Ҷ�:�RR#���ɽ�?B�V���1��K��Q�U<�"���=ƉIx���u`,^[��/7V�ac��S���1��*G1�:|4P~~�|�.����ͪ�����=�~�ټ�H��5�Q@��t|S֑�J4B$�p��;|L��r�z��e����s�p@����;ף�.L�w��M̴,~11�cjd�v�-��I,*Q�*��!o�!c�����M���X�n���{7&�J�l�����n댒�)�,����SZ�L�f��k�̘�����?�gc���̧��(�i����|&�<�����m/.o����<�����\��oגU+��P��xZ_��iW�Z����'��0\��{�M���,����̬uHT�Lg��]'!Dj�@�L;�[~E}q��e�T��_�	�]��X�k���>��X��6�с�\gO�1A5�r&)�B�:[6j����2:}w�4�Vb
��N��*�oӠ�GJV��T��f�
-��ռ���mxM
����J���HI<;��"p{{m��@�:S���
�!�3HvS���ݷ����)Mx��N鬈���U$�'�Lw]�Sd�',NZ�֮��G�z�t��- �OW�����v�D,���~�[�T#r��ڀs����������M�Kq��κج|�,���P�Ҩq�	ZVq��]iŋ���bC,�d��[(ĥ<LJ8#�-h�0\�̵��(�	|���e]�P���+_d����]
N,��,S��qz��ȑ���Ɠ�a��&"-8����p���gƌ͓�t��zz��@�@�9�΍��SA�Bq�^�n^$�8J��s���[\1Z,eiW�M�{�i��Ԧ����g5�L����H�<@t��x��T�s��Ju$�xqI�l��*���b�-����6�5'�'�̒�(=��ֹ�uwuS�II>���O���\�`\�t��I��.�C�s��Lo0���|��N�Nm���6�j�˭$�ZPq>�G�0N3�ń؎���l���U�J�T����ֱ��l�8Vf�L�'�<�>밎x����.I��^&�>����.��������j! �l�t��6Qy��j��B�{�d;&�Ĉ�^����f]���/�G�-�AL��+�FGͷh�Y�ِ<���,`�pn�A�S�Y\3�o��}R<��p(?��H��1�j��Y��jJ��HPM(8�-�4s\\���Ly-ʷ��I�);��Q�)M(J����X���v�C>�q����GW*���;Ě1�	ǚ��Ae�\�T�>�J�mK�u@�-���Ci&n[��/�\�_�j���/u�-�՝�R�q�dĥX5���P�Z������[����\ؤD���KI�.Z4�)!��:�62/��Օ���w�=@�&Bq�a#;1�Y�l{X����
pi\��cqZDp�^�;���~y�@gu����D��$���ks�AKҐr 	��iNe��C�2�J�FF��x��oWU�fk��	̘�s����ݾ��; 5�z1�إ}!�Ɋ>j���Oy�l(����	��� ��n:��3�<>����DY�eSi!��9�Ҙ:�礼a�J��5�I������m�IZ�V��o��d���ùY��1|��0#�`Q��G�s��%kT��P�Zk��U�v�̑�F�oT2O�r��Bh4��D��V2J�k����ZY`HZ[wS?/������e�yyi��cź�Ή��iBUfQ��"L)ۻؐ��q�Z�˵��s�?�fV�O��2Pj�b��V�Ֆ�P"z)�X�umz�)������A���~b>��Bgpm<�Sq��RP�)s�Gi>95�jJ�uU���oVe�4�v��U)��q�oa�A�6>Ė�J�ա.���w�'�8ܭEE���&h}�"�����3�P�*m\6��F��Z����D��L+�A�Ґ)���"��|%���>@}-N�q�Q�o��f ���'���+�R��R�1��d/�!?qS�Hq���,q��ƭ$B�m�F8��8��)�8��V��~�
Ɖ<$�P�<�w���Ug#Ax��M�p�%Q� "J>��ǯ~�}kՔ��q�zfT%�h���&xP��Φ�/�v$�7�����S�5�z�Ÿ�~L,�ķ}d�N��I�d���j��O��cඡ���(�����!�K>	�{q��3S��WF�	��&ذ-��S�$ ����L�����=&`��s�w�ƧB��gF1�O�/�����|���x����~�G4����c≄�}�2\NM,��f$5Kl�ZZ�����YdK�zn�z��QcA����L����Đ��I�R�΄V��G�0���xY�������%z֥��'74CQ8�ɖ�!k�cY<o��\{%�@����WcS��%��*n??���+��+ �aHMx�-ֱ�R��d,�>FB�lg��{��ۡJ DH��bGq�x3�s�@�q�J%�����=H����J��'���n'd	 #����Z�����4��B�anC,����9DՎ�l�(C����b�Xq���<����9���+n�6IÃ����Fr�I�.�:��*B5-�8M!]���	^kA�&�ҫ]}�D��A��*�Q27RB�z����3�Nsl\z��0�LTz~kqH-o�*jh�Y�)b��ֲ}1�ĵ�}�U-�iV��-��c�8�^Rv��t8%XZ<����U��q�� 1���A�oK":��ĥbb�a�p���S"p����I��k+���u��c��HA8u�~Cvdtu~���`��=wl��&�޼N�:� D���@/%��ꋳM8=�??�o�qe���d+~� ��B�_��� ?���@\���p�������T:�a �^�殺�G=6	���e0�(Ml���=	+����W������ �^"����t��02u\��p��}����k��\�1{R>��<RR?��=��좰k�iڐԈ��4x���T8n��%��Ea P�evq;�D���gO�+>ݺ��r7B�;�n�55��:C�?�� }�@��[�^ȝ�G!J�[�rh���{�ɫ"�U@.���̲�h�3( H�
[f݅���0
�E���
!٣~�rXh�`X�_�!��~���բ����R9Ϗ�[9	�>��7�we��J���mm>ZlP�+d^o���a������w���3�X+�h���m��
we�Q�R��e��H����ǌ���;tI��A��/��J�M�(�g&�='��Iw8%��Y"��@WK�1�Š��M%PݹfĜh-�����.�,�� `u^��ٱ.��F �w�2%	{��͡y�Wh�5~z�e��.�%O��y�<��o��lT��4&�grɾ�o}�/C�C\ T��]2e�ѯ�g���6iz��ugȜ@ڹ�[���B[~��>��>a��zr+L���[�o	�Nlb:HGHϹ<����o^�!W��(AI��{��~�mBX�EGkE'W�]��޲����y���Kۜ#����=��"y�p��Mؼ�;�{y���7z�մ�syv��k��	�%�H���s�sU��ah)"��*��Si�o಩�2��%�w
ec�"��GN�5�����{��؉�I�4����Kuۡ���1_N�I�&;�v� '�4ַMa���	�n>���p�� �P�F����F�%U�bj~��T�H��6Z��E�p��˸wb	6E/4\��s�ɧ�&��k$��'/����{Ѫ���|�1)���/V<���6�����4�;V1w׃�	�씫��VSj����+X���^�砓��4 �
%��T���Lb
����,���Rus�Ζ(c��0[�A�i�P�>PP��D�k�g	h��<�a�c�E(��4dom�o�GK˓i."zL�X^lEN�H�� ���zG��̎���[O��R �DXO����FA��$���U���}�a�k��Ǒ�&q��영L��T�����iF�r��|��zn��5���>׾?��p���;�J�I��TfZ'���F�R�"�Z��;_�� {UpGB8?�<w2��b�c�CI=�Y���{m�{
�i���pز��O-R��v��W@U��'�MQ�fAF+���P�	�����"�k
.8�a��j�S9,�����OG�})�b�x �B������`�
��`6p��ѯѨ��}K�X���L{}K����e�	"���Ŧ����J��:N�$���"��$�L�wN�Nu��$��hf��K�鮵 !&`���`ׅ��uR��!ҁ�Z4�y�I�`��X4�ܾ��I�5"�o�3<�P��p��Xn�wK�\Ϫ2w�(�!��j��]�MOG�y�+sr�- �_��FMܕ�x�|����'N���ĭwq�eW�
��1�xe	�q���>�	��n7�no�경J����)-�w5�"m��-̿wz�'ç�:S�����'Z1=p>КM�R'1�O�`�d���U���_�ש2���3��������&越���{��8�]�>AS�a��ͽO!����6",�qnY�0>hp!�U\-��@n��TtǗ�9SH2�h���9g� z��!�8�&���d����J<G�iL/@G߇A���� q��"\K���M����L�-�֮ү�Jۍ.�Z�W��h��*B?%����4�҂�w�#W/�8���sSZG/���b���$�mz\Ns�~+��=�����ˤײ'��(�"�˧V`n%���Q�
��"�-0󆐀]�3���R�-��a�k��Q����=����U,@����j�s?`�w6.YU�v=�^���||�>�UO~?Тl�(�91�G�'�SQ���6��?QB`nCw���C�Jđ���`y����Wn^��R2�!����ғ��W�u͑�+n�|w�Yp���h��2ף�/#�����(Jz�q�-��b��A�"{�ڰ�W(U��Nc��@+�Ϊχ]m��n�^�߳^'r��@�w�^PA0� �œe򷕜�EsX@LqqU���D1����)`��EG^d��^�����G��YS�9���ؙ�ziw�T�ߓ��1
��Gb}�k�"s~�swؿ]XMkzw�[��q�*]�_C��*\�N���:���M��y�H�e�;^����6��a�b�+3�_.��'�e§���%�[�	�*�{FAc����+���Eu�:ƃ����B`K����B�8��>���[@~̉2��P�\o�0(���Tڃ���/�
ĺ�C����P�;��֝V�����zk	x/f}�]e��W{��|sy�|u�K�1Q���EpQ�;�4��#�G��|�I�(�<��Q49�['Z���G9���x����*j��v0^L%�e����f�X	R=�DB�t�Ɲ����T��I��}�)������ƻڛX(�䨞v����o�Py](��&'�}������^��؟%!�|��"����x,��Yy�>[���*���+�&�<.�'/UCQ�.H.F�W(���PDh�(�{E#����I��J|�s�M��8������{̳o����z�x���댩��9o�O���wY�#�[Zͷ9�Ec&����PB����9��U��f3�5��|��e/e�z� @t��JP�b��p\M+Z��z:��ܩ��2]z�J�խ���(�Bt��������9J���Nc�1�)J\�ҵDCˍΫ�v�&����>���Ŧ�y3}I_m#R�4S/��}�jؙ��;o9�wB�..��n�T�V�Wξ�?�E�d��Jz�:�>���`pĊ���N�d�U��̒�nxJ%�A����fYl��q�}��
	�z3�|��ރh�@h�Lj��0����uѕ&&9�#y�H'����S�3s%����:��'�&��H�p�4���k�Lס�if����l���1�@Z�]!��c�hyI �5�HE�5x��m �[6�Qb�.(�1z봴[t+�*R�@5R`�8�CLw������VT^8�J�rIL�l���[�87*[I�ˌ��LM6�"l���> ;�����]��(*�x���2����j���)��<���66d5�A�s�|G�͕�g��?�ʙ��ҾE?�u$��-�;t�ܑS�Kx���ԗʺ!/a�C5��9^�Jm�|o���;	3_�h�J/�B>n����瀦��֦�q%A)�u%�eӞdM<Z�4�¡�j��}GPo��A�H�d��*ا���RRM�K�𖶏��	FED��cܓ`|i)�M^�	��J�ae����d �c�CL�+綡�(��t���������\܊��8��J�xO������^�.%3���ɨWI�����F�=6�NÔU��H;����f^�am�b'o�uv<�RRp/�R���T��N�s�r����>�y!,��JE��ܣ�E�3��~��\c��4�ݖ犬���J�	x��V�)x���M�j�n���	|�q6�dg
�q k�J�5�/�E�!�˥lG7���6k��A���BRH:�9帀#wlrջ*>�CX
SoY;��2�io���V*#������:�h�+p��ŉ�.�g
ׁv�W�]��v˺ޮ�mn�����s)��T�`~Y����i��.*SbX���|'�;�=�����F}�����cY�6�'�j6+Q�+����=��&}hf5����}����b�3q:�x[	>�}�X�	����N��=�QM�x���dw/q��
�pLm�[(�Y��B�;X���<�Z�7u��R�JĚ�?{I��w�z�*][{'F������B=���c�rL��hW/��6�l3�1��M)�3�=�/��9����O'B��\��Y�θMX�q��oP�9'c�pz>:�Mn�+���hF0zIO������^�oy�ݴI���v�.��]r�݌l;ݖR��(���|5q��kCٌU�ª����W�O��b�<6r�;�Vp�3���?q�s%�)��\����S�<���F2[m?�"�#�1_2���v��0Ʌ=wM���?,�P�Mf��o|���I��+��en޵��g��-�k|QYt�PN`4,/��0/�, ){�)�Y�st���wp�_γ욼"�:�Z�}�a�T�Q̎QL_��1���_����mϢ��m����mȉ+C�d�pd-�_�Ғ��:����-����ͼʽ���&�����&*�y
:kW$��k�ć��rV��gA{�@JF?�*
���/+�����M�?,!��3��3��:9",��f�_HD��?/�lƭv��JK�'�Wk�s+C�ذV��!��뙎� � n�]y^��8+��

Rf@(w���[%�p`�-�LkW�F6�j1��<��ejo�>(�ёvB������*~×k��Kq��JU%�㲵O�Z���� vD�LY�W�"lg . Ѐӵ=_�B�F��H�*�UK*�HM[iѼ��,��BͭC7�������]�N(�rp���#����QVXH���o�H�^���e�E����oN�T�Ծ◞��-�'V�U�
蟇U�K0����O��}'JipdV������4�7��:{ ��� "�E����n�L%9�b;�SoB;���m��A/�}�<��[B-o���" ��1cI&��i��\m<��C�����c�^��-��9�6�m=�X| 3�#�w�����䠌�3W)z����&8(Y�ڌd���]����Y�%��&t�i_ 	$�2����->j����X��!�8@����F�,��L��M	<eIu��Mi���@N����#rPVGb�����Đ�;�	#3�]V��t��,%Uԍ�1�i��SϕKIE��A�	>ގ��cͤo�<��x-�-���,�>,�Ho�!�05n�]ܡN+MQ�Кc�87�ˑޅ{�Cb��{����HXx+�-tהOVm���Yσ+e�J�����鄢�:��-��`��R��爝�U��k8��nNs�^�	wV�[&�Y7W�˕)��c�$1\����Ə���{c�f�)�GB�� !A@���a{7�e�9�V�"IJ�ti�N}o��U�!��&�݄���9���y�Ȗ��a�!��Vp`�V
�:tfv$�C�n˵���u�_'/��֧����*@Д���i�D��h�M��=\�k���s�[��:}�[,8Qǿ��H�����>�P���sD�eM*��A�2�G�4iN��������e��W��z3,nV�'��G�t+更�=�?��YN�nǡ�y�'��
]�8�q0?	a(�G��;q,۩��t�-�1��7k{\�_���MM`��P��5BA��ƻ�-O3)~�-���zne�A���\�,��
��J\�j2�*�GN��NA����|*z�3IZ�B��z����w�DZ�������; cE ��!�b+6���g@9c~�[C��;�T����%.�cL�2L�@t�������T�`��a����İt�a�S�$�5�h�\�����'� R]�x�O�#�T��q$7z`Znvk��l���&��v���u�E{�B�DӄOP\�տcZ�o�r6��w�+ &�@�/N�6�`ۏ�����Y_M��̥��&�a-����[��L=P��V?��Q��]k�V1�����=J�����=�B)	�`���k?�6j�I�H7��=��\���n$�m�/���	���"?'>zZ�i�@��ū�>3݄��	(�*w�O+ﲈ�懢�z���0�b:\I�MTK���ܱ���`ؒ�87�X�v�����J�՜U��I���83��J�j;ˮ��[���[\/�h��k��9�ê�\��Ym���gW~C�H�{��9K��}q{%�Vx�*ػ�(��uvt'�9�$���f�X��<]N�c�]�0	F%�vՔ�<�U��,л���'dQ��+T*��Z6[l�����b7�rG��`=�L��MgV�A|�x]��|1=CU�k��"�	�aЧ�c���}�RJ/Yv��
��.��/M���;�	�����8������ڦ x�!~Ű�dO.�Y��R��/���y(:(\����oRg����*h.�D[l^[�*��RrGxSٺ���%:ӡczt�|��D}�Zٞ�Rw�;xd�k�+�ph�Y^F�V����Y;+�w�����9��ۚ&�U�\�Bi2�5��O:�x9y�/VƢq�A0���ߥph���DC0Ϯ}ǅ+8�0�3&J�&!�8'XP�������.���p}�B�M��-�9m���&�4�rS����oN�U�s!��
�C�7L��k=�e�b#��&>�f�)D-)�ׄ&i;}'�5��k����U��O�1�X�� ��]*�^��Uc,���)���r��N�������my������&\i�����π��M2Z�����SX�v� 0ҁ'�ks�ύ�0'�b\Nd��̤fI1À����ڃ��s��ڇ�>��j��VQM#ـ�&)Ţ=�18�x��-_���}_0�9�$�oxr҇A���� b͆}���C��R�V{d\�Ůc���>�P�����D$ɤR�VDY�9j'NF�m�~�d��-�$�&��
tk�s��g��AK�S,�s���Ϭ���T���0���~��+a#���t���3�Y\�{���'?Lf9��'^�l��Z�g���}��l{�-��mvN'�ͪ��Ҝ�a�, av:;!�R�����jO��E�xC}�h]^KC�6{ڂt7q����9���C���982�oSV��7��I���^8���a5��O���r咇͝c�f�����X���h$"?��ɠ[C^����<X��HÜ��w�&D�>c�3��)=��iR(eV��6����&$~c�������@�'{*g\N��F�)�����c�*Z���a7�n!�,H�z}�H?/hztRw5��5�U@�7b��g㹅� Is�-����,W%�@���U0򲓅�5��;�$)��ښ�]�)�5�nM<�Ukr��#��ss��Y��%z�Qz0Q���^(\��N���y�Pъjr"�*��!�nE�$���'��hH�*��Q̟`z��Y؛�J���}��N�/-�W��{`�����ۻ;���F����'�:�B��P���4�M@|H�����$�k���Q���־��D5��&~�7
)�"z]�F�EI�^�"�;Y	V�qc:�h��+�_�E�L��C�o���mfIr�\�9.�J��/������ߋ�B�YQ*�X��0��/��2���`�ϼ,��Һ�g��%�q�p�ӔJ�(X=���Z|��6.�Gw�s�;
E!�lj�Q~���y�1ȴ�j�1���|+?��}bש�n=u���T4P0����v�i�jqH����ˌ�˽F_E�������d����&�0���:\P���ϩZ�0��.�O�����Q��NDЛ`+��s���Ƣ����pL~�I���Ol�j%���&^
{�2�..Ӕ�������p悓U{�>�yo�P"�t<\��+�Q�G��	Y0��/q`�FƱ!�m2Ĕ�$�~�r�J����2:��v�~�̧�����n��}�4PnOf"C8�'��< ǹB�8V��Ay51Z�ˣ��l�ّ�w,��p�*e{ț8�1�H����?�#����z;���^A���y�ɘ4]��v����\��y���9�2}�mc�`�Ah��Wl�f. h	��?I�\���8�=��с֟2�腺�{�,b�A���ȏR,��]�%�!�@ʬ�8�hʡ$J��S홀�53Bu�E:���d���1����^V:���h�ğ�xE�g�$���O�>K����1��G�/
T�6	�n����F���L��y1@ܳ��r%a��'��y䭻��ا�2[X��H}+� y�u\��o�;��O���׶N�6&�C_WQ2�V��"��Ĺu�*@�pfb��� 8TX〱��AH@Z�cW����^�vu�@{��t���j�r��C§��KE5���b��q��Mb���˅*�5w���"8�kF��t_���q�tj�wB��i�R��*��(Y��6W~�l=�Yj�J�$^o�p����4�X�
�)ʆ��=��,n�"�{p={��H,����64��i�E����dW����H%�I����vm�B'�v��r���	i�+b� ���s��h���I[K!A�� py�f�$vF_K� ��FMܡ�նp&����>W�L����(1�����#���6TOT=t:pΖ��>݌��В�����`�?RUΩE��^�K�Z�e)29�b0D$�?�'�L�W$�B⤼��t}�N�?͋�#��+�&�/'��H�<G����W�Q��4d9��ؤ6���}N=�����0Uۖ,�f4�{A�l�^ x(�/�P�m?���
�ٛ�,�q�g�s_!['<��:XI����@c(��|��ŧ&��������i�5�`��������oAuN�p�np����$���qӪ=�R�-aC3� }j*p���]�*��#kep��7/9��&M���e�KbD�r�f�@����1�aJ��F�ý;������h�pW�n�p�_�������z�NQ9-1-z��o]Ծ;O�2���I�לݥ�k��%<2�h��J��,t�RS ��O��5�cWtWE"��X2��r!~�$-Y��57��y�p�ZS��t�G����XՔ��!�Bt� _��w�F;�fg�k���5I�*�v����v��Tm0��Κ:�~��	��)�/$L��RpK8��m;r���y7!�Q:q�l��e�\�M�|,�����H�`�B�T}3�k�mk;�*����Z���
c�^��H}�3�Y���t��ǂ#H0o��."���za�6R�w!��2�\���IR�z�s��5 L���Bi�[���ҷT|�r�	�R<xʎ���v2����7SP��>��ei��κ�F��-%u(_�8�����+��$<t��-T��n�����=�����;`:w]��SDH���w����Ӷ?�'���lu�fC��u�o>Gk��7�zqj|� �%
�L�Ĕ�q�Kg�����#L�<��*0�򘺂�y�	�͜vf)�ΐ���&3iܳ�=�{�DL�v�Y������S�nV�*l��(�S�3�E*�����8 �Ş"�ʹ@�¿�1u�rG�����Ҩ~��h/��;���k��>T�މ��W�kwv|���ƚB�-[\�q_���zt�a�%mf������#Ia����F}7��]L_cd����X-���V6�m %k��S��r�����
�`)���e/[�ͅAЎ*ʏ�r����U
�_�O�%a/�KӍ��5N�_7F�Պ��� ��6�բQ�e)���R*���wçK�زf�"�f�)3u��&G��g�n����܌�;�Ŕ_����c��n���|=Z�n�;��#h+8d+��cS��������H��`�/��v�	�9$��Rp��C~(Z�2p�ڏ����Ԩbxe���H	�:I@�?��{ѐ#K#�U#�����\�

�/[����;�)���wbg�)i�g`�n<���C�P��9� &f�Ǳ���5��N�A�����;΄�B���jX���R!R5N�(���.��)�;�� �z����P)��T�����#X�`nm�T��#���S2c5�"ϛ�~,9 ���z�`+���!gV#�U�W�_��OB�Qe?J:�����}X=|����Ѭ~�Tա��L��k�Ow����f��;���\�T�\�H(w��r|���3"{���(��OW%lΪ]P-N���Dɘ38��g(F�	#�<�	�&l븲e��S���sλ�L
b�U�f�T���lzWȥ��mw��fz��:ድ���F9�&�ީ/Eo&��&�5{��2���k���׹��`�s�뾅����8���/�?�AM��果#o�U����,P:�T��0�Lɩ�9ܪ��F��G��h�I��d�{Cv��`�V�7�q�$ܻ���:h"�o�X�l��G�os�r���k��/��!vg�@x�~/��OG��jS����V��]u��H�#���>@�E9Z5h�G��^�[[B��+�U���c�$�o�;�W���q��*GMN#E
~Dsa�/s�l*{J_K3*^�X�acG�C�A1��-K��E�*�*1���
E7|���_0�3�;�.�O"��6����}��Sk�م�-HQ�s���`����"�$$
�:D��%$waҿ����g.K3Q���������ҥ�Y���ZFܜ/�����U�-�4~l�}g7<>�)CvVֵ�Di���L=�=��j{F^�"V��y�׾�`��U(�rh<x�����j�~��cAf3mJ	�5�^m,��9k_~q۫=�N�L�A�Blٜ�&K�c+��WA玊8��NA���w9�B��Y>n����	��S��M?�Q�٧�]	.���~���
i��Ѕ��{˴j�-��1����]���K_1g�^�cLt�b�����Y���-�`F>�E2��2aS\�.(��X�}�9	_'qn�N��K��@��2\���&������q��i��'�]����Dؿ\��}r X9�/�ܡ��"X����(-æc�;e��=>�=&H24xx��K�5f�C�G<�K�P7p������0E���UM!����<��T��4@L,ڐ���	��O��b۱��G:�b1�>d�ޕP ns��X�5	;���TbE�|N�`�*�$�s&�:&���H��{�fbk)����l����p�*�!� h����'s�,�mԶ[�2�E�'��X��$7|!u���M�t|�%cܫ���ߧ�V�����ER����ܑa�j��'LA�S�A�i:�^RqT�
*H�"s2��M�����t:*��E�����#<Su��
Y>յ�~�xO�U��
��XC�Z`k@K�$;F(����WC2�R�����~�S4��e�6$�9�ܳ!���Ja���3��M�6���P_�~��[��+E�V~D��+]h��R��O�߆E�Lg��-�<�]T(��S���^k��Q���S�����8	v�
[V��̎Q�L!��������.3����W��.~X�*%�d�����QZ�y�sTMU��蘭U�@d�ң�;>!�*'����|�5����w/H�y���yuӡ�Tg,;��݂Am0�Y"{?�&�8h<(
L@�pȖ�=���^��O�/xo����~YB��_�W��ݬ��Q���Y�Ug6Z�G��6�7��Y���ζ�qӹ�h�ٓKz�� ��� ��PM��a�'��|������4)��f�$B��!?!z�z�u���Ɖ��s�Θ�%03�-MdYBc����"�%(B���Lh8�A-�A�֝�T��dfy�G�T����Z?���0D�i� ������ �V�P}���Bݧ��j�AQ�%\���:� Oe�y�>��_K���}$��q)tT�接��9��2���6Z�Q=}T4�KQW���S��݋H@B[����Uj�n��O������_����3X��<c�Dz��[>���*��i��8�LR跫n�+S~5�KI��f���b���V�O��⺘C���le�MM��G& �eVY�-�d��Z���n���S�1$V��p,�`�Z�͓
��*��e�j�[�7-m=���m脢f�ϼ?.B��Ԯ�,n�<�8��y�e��EE��"�c���K2�r�U��]�0G���/����ΆC.�Ζ� kZf�W)ݐ�>hd/ܘ~�!�``ч@���&;��ܟ?�4Ϩ��v�*b���(b���k"��55ՠ=DD7b��X!�(�Б�!p�+�ﲃ�.]q~����e�J/�nlh�{P��P�e��(��cP�SdK����������L�φ
�d>Ԩ׊J�5�>��y��b�������c�B�O��o���:ey��Tl�����"v���U������$���	~�U�?�9��A�Q�r}0 (!�U�1sh䅀���~�*F��5��Q��M���c�$K���w���9��.�4r��)�Af�5Jg j[�H�f�i�(C�]g��ɱ��$4�i���X(~Y4A����^��_F�pxV�m[�)�X�nxǸu��#�]�F.�bJ�7����MG�kW��fD}sx�G��Y��0�
N\�x6,S���@�:�Iۇ��z����.N!
o�3�����<���fė=݅ھl�+��NN��{ߗ�4�5j[���&���N-t��{}*f��1���P�x�O�X	���F�a�2<3���X�t�ڑ���v<�"\��%��8oO�Ѱ�)տ[G��(�/�	ǢД(� �yI�zBn���R�b�:[��}��Fu�_�����M�����jXk���v�Z.k��`��Uu�x�ʅ��~���9s8R* 7Z�&��F��#\�Ji��,~�@�oN��'�`R�6�����lm{����78 �e���UW!���G���G�ةI�R��4�����TL��`tW�g�?ȏ��WXVy�T*��&�:�0d�2UN�9�\�|юa���?��b��ϥ��Bs|"��f�m�xw��X���.σ3�O������_�H�S/o�J[�wC��^�;���+E�5�X�&����z�d���PI�Op�.zxT�p��U��7�j�}�T�8�$�\%�@ޚ^�Mt�]�9�� �qrX��|o���(��:��̾�������%]Td\�o7p[ ��{���[��k��0����FS֖b6vy��we\­��Zc���6�q��:#%d� y��O�X�d1�o�?ď`k�Ż���|#�s��4t!&����W��Eyx��2̪/_sM�B�s����.)zE�m@�$����u��}$�"�'ng�;'ol��R�j��,Ԣ��gj��0"�ݲoq�8�Uu+ldNy�+]}ρ�m��z���lSK[��S�Qic��
I,M�uGW��� � <ӸZDD/y��$Yl�fD(u½DZz���I�r�b��mm��/Q���M�X�k��pF���E�5�a՝*HEh�@a�:,���.y�oE)������3/ڄ��.P�ԛVԢ�=S��Q�d�C,�yr rS�;��u0�3��6P�fa�D܍I<�h��8#h�x;<�:��99�P�yҪ�hc�:_����tv>��#�q�qz6�����C���AХ�6�m	L瑆fޫ���r�sv�!QV��N�#����NFr���kT/�1�Ċ� �A0nu_�'ȸ�[��Y�.���ru�F��_N�z2��i�c�_��ƭ��/�Êu�xb�0� F�=խQ�Z�$��y��1���4tXE�ۚ	�M�Xw|a�M�.�<���K猷m�"�􄙺j��C��.HI�,��>c5*r�p<���W���11�|	7(�� �
�W0;r�����q�<뵠������U��b�����C��G>Swa9��[:��d���>|�lW�ؤ6��\Z��t��^;��Nm1����?'�]Tr������Qˈ�����q�q_���[��W���bA:���QÏJ����"�����ߞ]��8o��g��i_��s�'
���!�\D� T�-�:T6�@��߁QKɢ�I�hl
�NKw��!�!�ͣ�����]-�S[�f���o��:w`!H�����2Ȭ�Ȓ���i�]ͯW8�`J��_���Ș��>���ᬾg���BZݣ�s���z�"N��F�)��/XE]D�u9�
��P<8��jc"��v�T0U����?�|�J��Kw
�p���AfD��7N72���O�!�&�׃�~����R�a�uk�EC�۹={8�ϭ_��e��u��K���$�'��*H��D���VV�G�o��:o3m4���xit�`��(E��q?�`����Tl�c%0��C@��jC�CʔK�~�� �gw� �6�Y�p1��ǮM,�~!uYk�h/�H�a!�Gj"�R�( �ў���1�[�!VK/0�[~>WK��� t� ���i���C2V"���oҼ���O!9�s�� #���N�C>���oP�'�㣿?����@i��þO�n��������K����������sޑGA�8��ڋ��U�;]��.�,�s�ZT��k1z86r�}�%y�0�
� F�����݌��ነ�BDba�e�O	~J1RIٸd^�i����	pE���	�d!�Zy9��+X�Il�#�*�,�i�]ȡ]�_���$���%�#z]��]lU��
�N-0>ج���%��*�=�p�C�6�.���5=�����wXv`���n�y�5�h�~������;Ȅ��S�ޗ��YJ�N�;>uh��l�ñ��p�`�jΛ6��Ԭ���A���N*F���覙�#�|-�{��
L��8�2�xY
dE��Đ.�nhۨ�֓���L`���� 8��ݖc���z��z�Cc�pR�]