��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]Zɬf(�'4�o^d5��o5�V+�����YE�٘tv~ұNVz��!#I�PWa���T!fj�T�(�Q�P�=�׭�[W������L�9��0E�K�M����C�N���K��N+����@9��x��ѠB��yPI�v���#l� ���F���aK�:���$l���X�2O^�lA�sQ#��ϊ,�5it��TƗ��$��ȯ���-<���+p5O�RD���<���bz��~\w�rOdp��>�W���?wȎ7����,�T �ras�2�IcE��#L{9���ȟXjI���`�62�Ѐ�||J�:ySq��!( ¯�O��ξ-qm��ҧ�rmC�<��f��UGW��R�f��~��B���3�i$Z:�s���w�v7E|y�Jc�x�X�㦇�Vi��K�g1��S��F��n$�_l@�L*�؀ri�a���O����\d��~��񟬰l۶�� ��v�������S��\�;-����@8r�3��aT���a/ɒ&H�P6آ����~����-5~�z�UDgb�a\ܯ�R�b��z�|2�Z4V��Ƅ��_�\r�`�I
e����b�|,絳��Y8�
9��XO�cUn��:��%�qN�1�P@#��� �Kd���R�9p5�����E��ꎏ�{@�Y�M���U����o���ϟ)����9ucC#�p�hЦ8J��~��\:��W�(P��� �^��aϖDX�r!���=��
9�.Bu��@�����@���}���Z}�����}pC<��FM�y��/I	1��T�4�dk��F��$��;���N)�r����Og��e�=�lZ[��W�6�`�d����Ed"�*�79gs��<�;�g��y���ť�Sn'l"�@5�%*�
+<Q9�3=���U)TGyn��;��0�%��]�m�$PÇ����
��S�KT�=�wWP�K�c�L��
�K|���D�tt� ��ˬ��s� �t!�xMK��&���x���f;.a6�U���V[]��>7`�r�?�Hl"��*���F�7c����;n�xP���MڂI����ކ�����W��rݎ�Tp����{��_�b������/Ĳ�f �)��2Ѻ��-R��!�c�<��u�������"*ܰ@-O���X�ʽ-���@W�[��L�8��:���#\g�Y�Pn_�G�v� ��}Ϭ��ZkU��2l�y@��JMNVu���`Cb���6Np��P=t��D�d)[�]�UQ`���VY������п����0�t���wmgڝi�5J�[��' ��Z\nx��Ҡ��p��4U���U�J��A����j诰�����0��'��L��A�TD~P�.��I�:��<\/���c���z�|k[X��ċ;Mk�?׳g�ރf��a&<%λ��U���N)�l�,�P�C(��n-v^�ܩV'����ÿ����X�$���p��]�
1j%�Va�w�ە�Ivi�f���4�;�S׍A�v�����0����@�$��np�_'x٢w{�������Y�����R�����4�,�v'}V@~c?|�H����qʿ�"��Y:����M��C[\g��(��	�=�����f�zW6�f���౲��_o��&W�k+/z�*O��ŵ~�DE(�<�B$��:�,��[ry1��t�o��G�#=���iU]V�Z��΀�gE֖Ŭ"_\��l��D@C/
�ƛ?�.>�ʐŘs#�s�r���r
ma�ZҜќO� �Eي~��-�v��;}l�9wF�D�,���I%>�	�8yG]��_}-q2�Y�Ë4��"qy�n|�W�:��'̚���8\�.s�Ș6��?㲻ҥ�b|:�jS ��{��[������:Aˏ?B#�MǾ:Z��,�p=[S��A��������(Y�3��&7R!�dm
��zu�3��P��B�6�W�_M��{���&&��w"GeA_���biv"3���h{BO�2i�t�t'�Ka/`����=<q��3��$6g�k2� �Ӻ�C9�p�E'E�^^�yN�������y��	`�<�x�gΒ�	#]o�;w�u�>�i���G�.HZd.�p���.�U��թ���^�����*B��,05���A���"E>a;�h��ɔ�oF��g��9����ǒ���@��-���? ��Y�ͤMF��=X|�nW�V��M��9�$�p��.4�	������5�p��s@C�2(;~���"���;I=>J���ѧ���'�,3\�.�,�G��t.}3
��E��E���ҕ�j�"W~!bz�� �R��!�� 2���:�r]Y�FMb�� !���*֐MM��g����p����A�u��F
�`�eAU�j9�ry���-,L�>ʹ�>�n G�B�4�8��Դ,�p��>6U	�B�P]��3��0�ݺ^TL��voL�7d�@���1#J��՞I�
E\ݹ�N�j����f�9�Ge���n��@1��3%��9��+��<����(AjNT4ăZ'}��3���O�O������<���x8�77I�LT��nͩ��ᘥ:!{���S���������Z���Lc�.4�j�|��R�L�~�B%�O���P!��i��6x$�\�C�G*Aʴ�<̖-�3S��h,%���q�*��*7�mD��n��)3j�(bc�N�$�hѭ�g6��o�,]b��LG@ N=�乚�3�"S<yD��
Q�զqs�\bG�)��G�&�����\Ģ��1�d͠$(N�!)P�|�v�g���^,9�B6�GS��r�����V�
�A{�Z�ų�~&7hi��vhc�/��i�}A���r�]��ʆ*XE$n��C���@���P��2s=$$��:ui�t��BE�E��zZ�;��X*�Y�!N0��~6�%E�SN(_�б`A�mAXy��7|u����XF��H�%^=-f]�{AwL ϰ�db��n�,h0�>1K^!}�8�N;t`Z�q���j_�ٰ@gZ��s��{x�
oE�G�
���W��̈́ͽ��9��M;+n�D�O���VW���X�&`��,"[��l��gqC�������*�ש��I����T�� \��#Sej�F�۰��(Y�%����-3�ƽ�x?|E�	q�c�ҤF��
#0����.%�=Q����Ҵd��4���ď]��x{��E��N�;���r8�^�j�gx�خD��ڷ<D�&��T��h^�|Y�/�&��p�F���Ya`����A����PFтWQ�yy��J�03��&��1sr򞍖�}�Z"�J���11�:nA똃6�y%�C�t�L����^�F�f8j��t[C�LI��}�g�j� E����z�2[��:zM��?g�UR�-�pK�uɴ�)b�1����kR�c���*ʧ��)���UTP,^�'������bA8D�m�
C���S�=,31�8�]H�Y��[���6�<;/�@�PK���/��?k�!�-x�}�N""�PYy*� M�.'b�!T,{,5?��l�xۃ�]І��*3�) u��j�9���n��a-��c��C�|�ۛ��{m!#�AQ�.h��ďb��G�K&c'�U�.��h!��
�}��Uf1.��.G��e꺨#+��R�>��j>9�O���*�4S��z{�'H�8r����( � ���ČG���ڼ��ܓ�.�5ᛌZ%k�~f m�� ���9Ccr <���G<���ABv����X�[Ud0�&�y���^l�^2JR�tR���@��9�e����u�H�WU��@�����������`�=d)ϧW�`� �K4>L�!ET��:�lP)~,��1�� |]�d�dHSp߀��r
Ƙ�[Q��D1�n�F`|�ZO��+1��(ٕ��Ǜ�����L%����'9z@C˅���`��22%��l�%�Cw_"=�Y
�1�!���M!E=�\��i�L�t��#�[�ur����k�����%���/�K�NF���#�+��/ݳ�TT��!z����������W* �	�7x�o��yJˮ()^2pD����p�Խ���m��~߯��[�C���F�݃�G�
�y�N0\:�����G�z�W�4�[�ZCn2��O����m�̺� ³Gh�����٤ܰ�cd[��R ����3�(���c���a���w�rj#�ԋV��vH2M� 5 ��)}������5F~�/,n�u1�߅��#�3 �n��ǥ����ot3�b�{�)^n}}-��wQ���#��9�qp�����w�i}ʯ�Mɸ�,hƱ�M��������X�"�����kȜ[ 3�{U'��iJ���"J��.��� S�} ��" "�R��F��W,V �&vo�쿣j�w�mƩUa'�|2��C��v�ͬ`��Bn$,Z��Lz={�3[���z��8{����wg���N_x���>N�Y�^����mm��)x���:��3
��{;]6�4K�W���AE�� ��bvuY2�vȎ
�y�=�p\Wо3�_Z;~�m�:-\���7�=NVi9k_,|�L��{Hm�c�
�>iK��S�m�_��>�F��*�u�Y��1P�y/D"��Q���f}ks�[AH�gN�T�T%��J;���)O�I�3I����V����$��I�K���Br�����&P��e�;h+�)X����/�H���g�>���0)��r�Hg�?}i��R�#�I�5���<�wἕ=�aN�*�DXQQ9���D߲�����^�Kk�*����z7!�]�1��&�v�3�j�Y�@��.�󐌯�-ee�(���ֺ�$�D4ğK�+�_�X=cO�PU��تi\k����u���~(�
��e���0����nZ�ٱ������	�^Z�ayz�.��4'l��rZ&��{��_M���[Y6D|��e)v�⌵��lzuϖ����5�ש���m^����I�"ge��r�^ړ�Ÿ_�,7�L/��82�X��z|[��k��`$���M��i�.��E�W�M�yŐ�kx�n���y�~���?��7��6**��[����q�%�M�e�U�;e�zy.��O�,h�m����������?�8l���&�yM�\�W�qas�Tr��