��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��@ό�����t�O�Y��
�*T���]#J����&o����(�=}�3a�;���9 r���ɼX,��m6d-󂅬�ea<^��_��eZ��Ⱥ���^j݄ �܏��3#��<�#R�a������Du�[����,"0�ڥ�3Q�=���������R���_�
ШW%T6k�d�Nwnʅ�qWpf4� ������e�R��hE%&�U~���Ӧ)x~��\;ڂV�o�8�'�k����s�(��MWc�\Ͷ-薛/we�-�_ [���	�<`F[ZԠ�+�|Ϩr�?>�Jq*�%u#��t�F����m���G�h��a	�ڏ�.'��%�+c~:F�����%�0���w���|cg9�J�	n�Yv<����fthv$'�z?ϖ}%�S�N��5~�c�ه�(�ɳl���/T�k�Sgف��&O����8�&�	 �h*�o���wD�*<PH��iR�ֺ/�����F���(v�B�A���'��D�k,uj=DZ�0�F1�R�e��*����|x�z���ܖ�c�O��wL����z��9��PA�#.�U��bڏ�,u�b�X�]�u���%���5,w.!��Vj����x(Fj��`;]�=�hjYɈ1�`�<����7/~�B�����9��	���p�n7�#�%�G-��������4��r�/8�o�����J~�&EBT�9�%��X��O�C�$�_�Ƨ����Y�v���� 4��{�Iz�����&�㞼 �0ҭ0?3��[gͿ��x�z�[���|�&�o�a���cQ�^6즦d����7s�Ɲ`���cb;$� �K�+�q*x}���ݿ�<�k��g)���C*LR��O�4XM�e�8�YNp�5i��CF�E�3A�88N6�:��/1�M�eY�R�1�Ԁ�5�^o2����M�<���<������cd(�|�"���M?fВ�:ߔ6�d)�'��7��~��T\/�+�t�/�K��R2r!w���όw_&�:c�0��1�h��iLo�'���uOj�E�\�
��Mёd�l��ʥe$7�B��*ѹ�;������V�2���� ���չ��\~R�Dq��B'�)��}AD*�:O���mᮊ�cPKs��A��Ӈ����rh@O�ȈV�#�	3�x��]HЗ��E��u�>q>W$�|U ���G,) )�D6Z&~��29�����DՖ��������+2ʩ2�9H�ZO�v��(��z�k�ӯqܮ~M�MV[g���k4
�t[!�� (���v;�d"��ʥe�N��;tC��w�
	S��+���]X'�GӎR�5��fC{�o�'���9�"1x������B�p+涬�ɉ�!ۆ{�����k���|o%JA�z*!�7w�Ҳ��F�߂1[I�k��"5��sԱi�B�o�{6���!t���I��Ζm{���f�7��9v�HP�PP�v�EbA{7Y:��йj��d�g��l�g�n99��D7]�aFo�a��T��c�K�5�&�$�z2)yr��KC�_����e��|�����r�\ģi����Q�U���ްE���֚[�rH��S�:a���(I��I�O���4�z�m�N��m���(݈g-�A�;�b����h�)~�E� V���v8���MB�グ�{��*�7�
<$In��G����
��7*]z����"U	�ɵ}}�o�[�Ih8{�N��!L�U/C�g�Q~:P]�)�^�����D�>��S��LMtGۥ�q�u�S�LS�mЉ�=ї�rm	ЫS���-Z{�LbR���������O`�Z�$$�[h*�SMU@��i��
��_
'����a�L9��.����sL�9}ϗ�,��l�o:P�?�����!fۘ�9�?2bk�ǢҦ[��2��}!ܓH:�(�Id�R�z8�"���M\n"R�]�����ÓC{���8���*4����C�Me2��&��l#j���cXk�h5(�{�9�\6�9�tD����&\�Ȃ�in��٪�k:\�33C�9�������v,j����g;��=�ia^	:b��dAD[Y�e<t��3������Q��P��"���3����f�U~R=I$yv�F�-W�(x�`N9���v/��)�~���F� X��M �j���S�:���ц��^�PI[�Q�\�x���lA)����C,k4a)�!��f0��Q��:I���{5���[�l�nJT���e�C��go�I���nD��ǓL+�$�	�w�oZv�pdO
%�0�(oLaC�����3c�'o���y:�G���ś�LK�����/l�үc�[!P	����x����=6��9����S'��|�e<
�)�}ǌ{n�sҍ�r�%��N��.)V	��y�xrJ-�Χ���w�	��I^�AU�U�b�_2 ?+|y�R1 e��xtؓ6�F�"J�^�M&�˓ƒ��og�n=l���IJZ�>���ȳ���<�����8��J�N0���{"�l�w���s�(įr�F�aY����;c[�&���L�8v�7]j�&у��Bd�-�j!�UY��Lc�a[T߄1�O�εo^&���zdT��8&Rc�Z��0n���.���(D�!�����	���k��44��8 �Ս��������
D��:��ڶK*�-7�(V���ȔI.s��Q#l����_��ߟe9Us�o`� ��5O����}�P��+	Y�����x���o���V�neL�	g�~ha�A�w�^j»��IcQ�c���]ܫN��1T����6����bM�����Y�?{�#�R�~�:THQ���^y�ĕ��ˣ�����~yx��oG��&I}��Z^�d"��"�o�T�)_Upd�Lq��\`=O'*mW�6�� �����*YL�sRn��h(Fאl{�p^�h)�R���;�+�YC�/�)����f%�l7�612$�%X^�O�N�-���1$4����"M�b�<cK��Ɛ�RV'���u�"����Jn&^l�V灨�����i�X|$+���''���j&U�l���!���-��0��h�睂pBqIDg��N�#«Ԭ�y��{K5ֽ�%�]��`bB��T��A�2��(l)��q��K���7?�и��[��8�J F���1eH��k]�ӖΖ����e]��R0��M�{�Q�����FED֜W��ys��y,;���^�4E�ӟ���I�A>��I~m#1(?m3Ɠ8�%���o��C�q��W	���иm.��Y
�w������bH�����5���N�4g���2МnÃ�cR�T�7��
2>���6%S�w�Qv�/��=�R4S�ԸT��6�r#�=�m�I��y���+�ni��fȚ�r��`��Z��T���9��q0�����I\��ޛ�KO�/9��@�Y��I�bΝQ*-�VǓ����
C�^�jD�^ ��S#M����@�f[X�_D0������x�M3�d��O('O�_��Hl����9�j�&�Wԙ6���CA-�*������%���I�.����>������?u��]+����,O�~���08�f���~�+���K��II�LȮ�It���S���#�C�{Y�lrcja�p[^F�T?�mFm�2mn�=����(Vm��+G��Yq)7�i��_�^ �CCaE:Dn�7�D�&�L܇�\Ɠ
���I������TC�ۮ�\F��k��b�-�4�	,	�VG"=�/�T��<��`�_��Th���J�Q[��fq�=��Yӑ�FH�~]\G`ֲM�+S���n.-TYl\?�6�B��b&�[z���QZ�&[>GN@8�d:z"�Y��G��DFG�(��P�"��y�*�..�X �-�c�	��,�B<��p2�G�J��K��`4�C(A�<� ���h��g����f�Y�ļ$�/:�1���$P ^���SY���ɴ�˴=�?2cM;���c4Z��X����0L���^����l/�2�\ޙ�&֫��ߢ�/�Q����ˋ�����)����Ҫ:@j���L�e�o,����WE���@-l�ӷk=�%A���\��h����P���%*�OIn���P�y��?�CTG��� �@:p֬A{j���(��L���D,�����Ĉl����m����yI�91m)��:c�k��M�� ��r���	�����ș�/����.����P�� Jt?��� h���&SPBCG� �a�ڗ*���.��C�B�ĕ����K��N����b��iɗ���C!�Z.�. aG[�*]�����;�}1!!id�Tb;Ӗ]��M߾n�,�Y�E��K�2�����.X�Iכ�l~�����D��>�"{����r�������!���P�k�ӗ�*�[�������n����Bm�1P�V^�n�,�+6ܧ��ʍ�2�Z܀2��� �YQ�^`@A�.�W����!N�/���F�nBx��. d�Bf��.I�G����\.�:�L&��%�'��i�zNjs���^~�䢞[�`��ʡ�n3ݴ���9��Y��HjǸ����乛����:�
&���v�4��G�Sg=Ȭ+0a�{+���
�^g�"�{)���%��G����Ԫ_<�J1���N�,l��Q��u�����c1�񖌅`��V�Lwe-ˢ����n��I51Z�f�&п���9ٴ��w��@.63X�1���l��8��k~�p��T�`5"֜�i��T�W�(0�s-����>ؗ#� �r�۹��|8�\�be�R��v��>QI��#��h��&mW����p]u��W��B��]}��h ��W{
V�mI�d�'�����8���@������S3%R-�E�rx;�ңj�F��Ƨ��Ę0I�c�mb9zF��I��g�7��ߕ�R�w�)�5{��y|��@e���M)Xj'�=��#�H�e;���]۝�)�VX_��g˱�Rh��Y�P[f�~6Uc�&5=�՜�
Qh� %��]�>����]\����>�ܷ�/�!��A�a�O��6���fg>3W���� ���h�b�	�zW���݂�=�N�N����2�	1���j��$kk,����@�ѱ��*ؠ�\���Y���1��#�.wo���a'ʊlk��M�xьM��:с�-��lCM�Ra�^�P3����F��/�j�Z@Ǝ����3%D�o��ry���V�n��P���'Nv5��+O��(l�����Rb�pg8�`:� �\e���?Xg $������[-<,�*|F�'�慈uW#�}Υ�Z�r��j���QP�1��^���?�Zյ��:nV�����<ʾ�w��#j[�[k�(-{���&+,�1�b"@�5���0��!���ڇ�F.��kP@�CMl!�߾����]gi�vt��t �«&D��R>�Q:播���CV�3lOY(t/���b�I��w}��4���<�~Fړ�V}�y��k�=�k�qL�����W7���"�\ɩ/��^j,�D�W^�l����`�I���A��̗�H:��Â��,�F��=�����&�+�t#�om}]�Xƒ���e���zr���n�I�-+RG���D�T��B[����K\�������V���\Zͩ	W��N�X���N�;��g=����+\�s��R�={�(M�]�[��i�ֱ���4YōI�7�SGG��6�/��w�_W���(N�h�	e�u>V[h��ZU{%)�?Ф�i���O�;��A��Q�3n�XK�8wz�}[Ģk�N�.�	_H���;˷�T�i_\vE�=Hn��xj�o˿~CJ��g�YY�{���V��kR �1��O(,z4���-'���}wN�+���10�j1�A� ��:�_�^+l��Z7�f�v*q�J���7���
�ᥒ�!?\a� ���f٘���ڮټ����_�~.�by�p��ef%r�5y�FbwJRtu%npQt�g�u�-�\��>�q/k���N��EKSW�Q��A�h�9J�Q�m=Ív�!��V����1$�����C���d
�S�m�b?ߤ����: Ǌ�^��|)Z�t£�)3����wW?���0)|=��e�Cި��;6�ŃO~HV�m���ja�9���ؽ�.3�� �����oG��Gv!h�1����0��M���X�7dY����*%�խƛ\t���Wϰ��q�W��=]f�R^��}׭�!�l�l�6e|a���Edb1�^I�ȁ�8�W��J�;7�� O	C��:��@�~O�}��(w2<��u)#���G�S��\x��~z#���1��}����.�ǅM��	^�KJ��QCԲ+-��#M��/{�'>��v�*��B۟�c�Էf9ޗ}F��2k��0<���tB�p.6�	��y&��yCq��k
Y��C��k.�^TXr*��x$r�o�lm�2��d�\���w���E�����;��=X��P�b|v���ER�3N�E���B@-169���F~,�[u���X}�x���H�ln9�
O�ΊV���$M�]���_���i���y��<]�2�E���`�����ö>~kkV��`-���%1���ۼ�t�5�:��݉� Z�t5�z
������f�=��`��������R���\�?��@��������G3�c����.������88k�d��xƮg�2��1N�7�����$8R����Ū��	��5�`�GH�.l�����*�D��	�w�S���z
)��Hp*-�@��웴'�ȧ�U��u�̦�~{�gB#l�����A��8�vL����;pԀ]aQ��KI�a��枂�#�9�U�y	����-a�W��`��d���qX���Ȏ/˃b7纖3U��1�@���ۺ�.G2���9��K׹���/�Xd��ƵІo��e��Ą0/�c��wf �7���~��mI�vW�r?�*��!#���I�;��$��,L~�m�s��_S��f��cl7����]'���={�ŧ�8^�R$��%
fJG��~)C䋿0���3��'��X��h=�{���@���wd]0)���m��K��:��v�[����.U�E*����yCm�����ޥ��^*/���2Ʃ�Z�Ǌf�@��e�'��v|O���:D�����q�xP]<Cj��x��5z؟�;�b�j �a��4c��]�+��*,
j &zTM�ĵ҃�)��� �퐂PӬ�nդ�l��y���5��+<�)�&�IKCW����f5͍�DiV2P�~���FФ�G��d���2�D�]����*�J3�DEǏ�f0��u����0���24e6�ٞ�+��;��{�q�[�L�<�$��$ ʒ������z��=�|�O�o|���!�GP�$(�:+t�L
*ɻ�eq��X��b!�e��us
�V<7�O���&��-�B0�S\	�-}Y�G��	��O����N��ô��I���r�(���{Kc��*����ݹ��mqzw�`4?���Q�(+'?����^���'��@r�>��Ζ4r�Q{d!��$$��iG�����UR�P{	5����:E;��͡*�ߐr�:\C@���MA��T%�,ʕ�q�}2�=;��!�����
 o�e���.�����-�5�6c� ����^}��&}ׂh5;�|6�tOPB���E&}E�����
�����S��}=��m�A�P4��~��ﻑm�";�̔��ŧ��l������m���_�O5�����U�xX�).�����g�x��I����^yB
��X��aD�n����<�*��m���cD%�4�80�OL�U폁=�+^����\��8d��{�]��I+kqD6�3,�H_S�k�la#}�����S�Pp�ޫp�*�K��
�r�=>�������)���A�4T��t/&����?�,(~�?P��c��<�����Oo�8��)��b����WOؼPV�ҭ�e���֩�i+׀&�:*���(Re65�eG�O�)�D�]�B����������=��+�i�8dHx�P_�*�������B0��X7+�5�6b�j)5w���>H/d|��LU,��7.ڵ���;pܼ��ڨ�P�]24�Є��GG�D�����K�;�N�Ң��X�g^|YI*ߗ�@N!f��32�!"�N�����	�I��Gr�@�}tP�oX�/_��B�}�;�"��?�%a��|�A���BR�]�O)�G�g�0�j����{�3>{{�%�r"�/�=w͗���0��D�B 0����8������ۥ�Z/kߟ����@��έ$@�Kj��5&D��(��FU����f�$Բ>������k�V�I�B��H-u���������KQ�B��p��%�a�ؗ��:��e=Bt'���?����;QS�a�����ǎ�7����2,�M�ܗD��<��b��c�z�p����K%�B��7�g='iYMnBh���杌�Ʒ��s��%�xe��<�'��6D�,������u�LQ�zt:����S8
Z��(WI��$S9���cb�vo����r8�Z�/��ު�jgv�*X�VHYs?���.�)��w��V�F#z'(|6&F�9�ٜH(���s�Xm�V�[��� �ȉ��Ш���#�MR���R���3�F��nWu/��.!*��Ʊ`7��s��6R'�û�H��ߛ��TYaOz�1f��
n�ZJ!�4WYܬ�LP�Ͽ��X)Nb/=��Q�Z֩��U�l"9g)�\Rb�5��������뀁�>���q�Q��~V��*��	XU(��W�92C��A�N������W�|�[�H����F�O����ѵ���O�{�+������O&Ŧ	a���U�S��fZ��I0�4W�hIמ����ژ�`�@@I�X��r�Ue/)Q9ȝ�UXS��K(�ih��e1�"۰�#2>)���aH���R��p��G��=g}�o$�cQ��!yon��iN��r@��|v�y���ו�����徏4��)�@7?Z����@��E���/�A�ϻ���D�%?h%���֫��".��Nyѕ�	�ܦ��l	���U S��5�z6+"���$!:��MS�#��K@��rΐ�:���V��j����g�l_A��� �����h8����j�p��?�:���F�`,��0�T�����k�>���W0Plv�]�t�5?Vŭ��5�e�r��7&�ڏ���������nmGW����N9:d=���p��@�%���)���d�\!^�a{�8	�C�'��F�Q��8=[�~E�l�_m�`*�rY]DLRhJh4gW�����)b�c�X��,����xv?�P����B4nƸ܉����}�[��B���I4��{�dAVf�!m�L��ơ=�c5��39�.�`���O|mY��i��08�[+�������EY�G�<@�od���!>�}���5�N�~��/dH���+���y�4��W�؋�����g5���%"�����F��~ܲga�����%_���𜿘2��n���B��'��#�GI��+���P�64h�/�n!����d�H� 7F�ۅ��e_Vg�3��!�� ��=�ƞ$�(�`t圓}}�OӚ����25%y�YG���"��p���ZD��3��Nb=lj�磤�Egxq��,m���\L�O!l�HsW3�P1�"�5��k
��0"J�h�!�΂"�5�sҴB�˫ݧ"�$�DsoCl����B}a�Hbw���sTb����t�����J�?�9�V����:� i�/��j�^M�˳��膢,|�̀��O���w�kZB`�P���k�NG�x�?�#l�����r�nur[���1(��k���rIK��W������×�mxr�^Vڈs�,O�����-�%�-�ġX $��hz��Ͱ7��3Ey��%6{����0�r����� ����|��T��|�����09���^�xmk�r��%�6�_�ep��RF�h6��PI�Zٗ��+${n�'����q�Yҡ����9垆:z-���g�]��EkSQ{�$m7[���!��2�mG^Z���R׾��16�NJd0��D���L��1�ߐ&v\Ls@q#��B�=�"I^�A ���`��>�̀v�̟��&��S	x!O�!�c�O��t聺���QVǬ��s�@����	�����`��jJI�P^�"�z�?�H�9�F��>��Vĳ�����)p�����I�����7M`���*��3�&#v���	�f��W���3p�����&_w�W�*�}����	����w�=���
1=�.�|��AIZ�+��'�� ����W���&��� A��)d@��*#�xׯE�*�{�Msr��6�%o[gӃ�)8���,+af|���s��[��3RЊ2�-�ҍߡ�X&�y�=�R���s�&T$�� K�:i���ఢ��t\"����� �O���f'0�G���A[9���E.b��~Q��[�?�JVQ�wc�Bz�s�O���Cm1v-싍K��oG'?�Pc�%`nĮ�9i->/�����b���7A*m�`�R�8^���̇�I�pKs��W%u^C��Mi�"�N���t�v�9��A�cJ$���ˊd�H�ǔ!�� ��b�s�>BF�l���P(�5���o��4= n�Z�"1�������R�e�{8N��Y�;�W��CVI����Y�si]��s^�W%�p�J	͔Y3�Xp�lA��j ??�+G7^��.�d\n�鿧����ŝ��l���x�
+�k�#6�5m��c��FY	�R�y����M��&v�������2�r���j<�,�3�|�_���a���?1��z��$C��R\P��1�9P$����@���:����y;�<<���3�x�tۃ�wܭQ��x7A�ce� �ǵw�Ӵ�P-�����:��l���J��I��>d"S���9��o ����쇤qC�mY�}������gk���𣮅a�:���]�Dc�h_zI��3q ��G3mn���~�<���T
+��<�h���R�9�O�k���ۓa��ޡ�6f��]��5 �YN����~����wΜ
(2&'��qj2�z��͉kV��D:Cp��o��f'��.�]ݜ��N��/�H��þo�ƙ\$��+˷K���S'�X�dN�C C,	�4�h#��Ӯ{��*��I;E|':�������{�꺉�|����d������^09Q��S.O�I�k���t�	�Ǔ�o�F�'���UQq��w��~��~y�[���nb�R�]�m���x��[����Ϥ$�e���4��ٕ�K�����8�e�/��Q��X��e�	h��O0
S�
��!m<�{�E���]�|>��K�S��K��nË�j��J2?�C�p�i�Ӡz�ي��c�sţf(�W=�Z�<��/Sm�`M�ۨb�Z��ٷ��o���2w\{����^\���%�.�c�Q-ݻka���Ѥ��$_��B��5+j::�p��,�����V��!qv*�6`;̗�OzU�O<�s��i�x���%W��������D�������K�%����(7[��(��"���vƔ=]@R��'Dp��=���uŔ6��C[� ��(���aW1�S�8%�Z��K�OE�"�]/���9�c�}�ɪ���F!r���g���ܳDo>���.���/o�2��m��*v��/}k�_�D����o�����=EQɩ����lr�8�k�5E&��e���5)�^i�H�W�]o%(z�0e�u8���b^������q��0��_@��m����Na'���950�d�-I�����I�N�9�@6��:L�Sv2_$��V�w_<:��+����2¿u�d��;4_���/������$#�w�b	�m�OWop��%oC�Sߐ��Į"�ϫ�h���2�W��zi��Ӌ�қz�W�@K���O�!	���e�Ꙧi��S�6d���j;�f�T����"�Z%�t��^��'#����U�bp��mTr?��}31>�0Eg�g�u�wA���V����;ke�jh��Z��;���.��l����"8�tzR��@�Bn^̓9���uBN"�yE�D~�!߰̈_L�>�a�Z^��c
e�+���M�^F�ҕ^��R��2��|�Uo�BW�&��{�հ��.�H�ҍ�z2}��4��Nf�g����OG��:k\�F�ޛ9RS+�OҒ����}. �l�R	��W7���Uy�e���s��>DG���Z�3�qv��wk����C��zv�@�� ����xg
Ye$�,64��(J�#�V���J�H �Y%\��9丁�h.��pQ��+Lg Y4��8د2]�}װ)"3���$�!�a�}����K]-�x��TL'�&����5%7+��W�%����iX�!���R1�FK;'3��eޭ��E�q/?����ZHi�0sN����)�m �iQJ�?L������R����������]�Y�YBa��U%k�$��J}�n�) ��or�ݹ�èH͈LI�C���жYr���&�t!���Ϥ�����_�iSU
.�%�W;ƣ�U��[�U���c+�3�#1X�X=$���l������p��E���,1m��N��σ���!.	�.�صӾ�D̽�\��6��In� ��I�O���`p����,���t�Q\����Z��+-��R۩�F���eR���E�T��;����7���Ӄ�=�� �]�1'P�F|��?pY��Wڭ�At�o�St~�_XN��a��d�����)�63�h�jP$��M�&w���g�N�P�n�d!(ڸC���h3;O�!;��E8��p#o��ʠ~4c�H��C�l4�h����w?���mZ|��+��5�|
 ���)`�
tva�|b�m
C����q��,�z��C� {��-�>��M�t>�Ύ��J�9.�zT�	��N�>���?⿿�	�5��K]g�S2l<o΍�Ī)2�'��Wܻ������k��xw�-�9�_6�G6�]�/��_�� �� ��+��S��0´ݚd/Kb�j�?��^WO��8�|�F����̰Iu���޾�A�-���k�^��}3r�%��!��!C�mڥ:sy�ʣҊnVB�@9�ˣdC�S��4h|�����C��I�[��s6NL���J�$�2�^rL���0>z�`D��~�ގ�;�C{o�rD�|�-�����xx$e���#��_��Q� �J��4s̒�2��0\�G�5c����2s?����_tl1���5�!�n�f?ꔀtd� ػJ׋�$���?����B�a���4=�v�\c��׵�ĆR�9m���� ��j]�	�Q��IT7~�Qn��ڠxFi72�{h�)%�o	a�z����O��fʙw�(��-��q�f�
�[}u�߬$G�bC�y�ϼ��e5��6���0PMk��I�s�	�q�_W�~s�̔�83�v[ߣ���HS�im��'$��YaP�YJ�}�\~�f7�{`�� o^L�B����q��n��%��d����m�o��!��d,��
��. �<�c����]������U�O�f���vӻ�ܣ��)����^Xb��X%���	�a�jCz�^̿BA���i�!�k:�o�qi��͔߶�6����r�0�Gg��������v�(�鄐P������0�*u,�l�TW���Jr=��V?&�Jo�weU��D�~�D�p���7�ܜ=� c#�C���46�F�tl���_�Kp��?�z�?M}��I��(�ae���\�$�a�+�x��Y���q�?"���{I�7�y��6E�+����'��G�?$iB,.Tm�!B�ܻ<ez�١tf8b��&㑫-�졢�"��1���e�%# p]���K���{@���2���͹cq!k�5S�]����-��3�˿=��{�իp+�YR�=��ĿC�,�8q�����F/����.���2ك5ze1�ys��$݌G1"d���˔�8��4ݳ�����!o���#��р������qt↿��>e?��*��]>)��}&�}ڗ��C�n�l��o�������ӥ>��Q���q�?]�.���1�y��+�q�0��H���2���<��3q��t,B�����t����~���n��^�f;W �u��PB|l�bW5S��T��&659���~�j;>
��ïA3Nt�g{����<��7Y��.xt)���,?�h9)c�]����xP&�3�AS��+�."��v�2̞��k�i 6�%LB�oi�Q�%^¼�P6=8UnC��6	��Rk��������a0�Ո�t���J� �U�Dx� Ůz����@�^�E��2�[�Yx��~a�\	�~t�O�
�p�����4G x�����~���\&��`���~ �/Nt���ߝ�htT- >PŤ��|vBW;�;ִ�!�]�(GFG|�1����lUB��&�b�0��k�4��8�j�@K!���4Z�r��S`�u�Vi/�=-p3Y�@��tR��5퉚*���z5��,�,lL&��[�����D��,�m������>"	��k�~[K7,�ƴb:�����`�V��|[�S}2y�^4���x���]dS��T���6kﱓ�9Zmn���������� Q ����W���;:��E��¸%3V�=E�=u�vh�RsE�G\�qZ��*`�����<U�������>*	�Q�H��uc+�wD�<�"�/kZ�k�f�؆^QemĿQ�3�jص�ؖN]ޗW˻u�~���{�Q-�������d����{���͠��$�hu[�K[]�wC�&�]�◆���0�z����ف��(ƙg?�N�>g,��c��n�5�>�>
6Fa���:�}f�Y���ߨP�X{�:+�܆eƃBJy��L�]�@�N�Q���Ȣ�4V���ף�J���segTYetU��{)�ڨ�Ag��fVD`���;Vz#'Mk�;�Ζ���e�9�� ���2轜�7����I�ԒiSCy%��S�,���a��U�}xa��;�ʷ�2���
���?���I�����r��g���)�O������\@4�g
���>�H���e^aM���M��2E�)Z���2��&ִV�i�|JL�{��-�Zɸc��1�r8��N{$w���D�橵<��E]ӛ3�~gC�I?�[jE���{I���PFgD`�� �e@�S,��*��h�����,���8�D��N?��e�=;~�,כd?��٘2��l�ˑ
"�a҉&�
�M�e�p7��K���Ɠ~��8>������*�I8�T��1�th��\A{�r��?_ڃ>��p�^�|8Bo������x�/�H��KJ��,�W��L�3_�,Й���ऺ4��E6R5�h���g�u	�#1�.������F��>y�2T"S�W^�'����vV�;�[�Kl�54��� U��5L|�����B"k#`x�Y��iY����f�������:~̉4%��2Ɇ��b:�_,��M#�W�3JוMMsM.�����f.&���4�!��;m�@�����˨	�8�4d��4�!�l���?#�FX�@���ꑶ�bIu���mB8qo�����x��Ҏ k8t�>ן��³v,9����R7���N��G�H�F(�=�@����j���������.�|��w�}������u��`k��Cu�`����˘��=L�"_�o�����̼�y�-u�9�|,&������ġ�S�]�a�t�ë�
KY4ظ��f�#v�ܢ�c�%����&3�[�B��L�H�����g��{ �����]�)&����8a�R�G%Eܖ�OB�J'^�O�	�0��v鵣H�b7�VQx�?s6�Ǒ��2y"���I�g�QV!4}?v߹����S�}
CO;����y���I��N6�ju�W��6b��&=nSd�g���K�&�ǯ��nP��SP�kCܖҪM_':+5l�6�q0-ɵȴx�U���9��ppD��FL�H<{��Pli��n�O�w?ne>�/4��ΛLN��ܸ�|�zP7pk��f	T���5���y5v��=I`m��|��V��z\�`��%%�����ig�M�<��&N�����!-�L2��N�x�|�h�ORL~��F ��=A�1�f-g���K'����iW��<s��h2Ř:h�Bl�\��)������"����s;�>� _�
�r��l/5_�▙�nJ��j�n���,g�SR�D#qX%�r�D6�C�n� ���d����/O�P@#Sݺ��H��Q��z��w�$��l[����l�X�˩�@�'"�&`t׀����w�ûLF�"�ދi�zh��<0��� �60;|���6�9l�ѭ�5������T��1l6Oȸ�.q�&L:������@v�K�A.L�J�N��^�F@l�T��G�5��h�wu}Tʹ��q����YC��I� �|�,��=O7�ت�mPF�%x}pP��ݚ�sp�]���&D,�xL��F,�o�E�
��|kG��c �4���훪fWEF}$҄���Y���L����Nԝ&��>@G�G�3���]	u3vm�Q5v|i�����$�ё�����y��h��l)����܉�>��Y���ͱo��_�x;�r���ؾg��JV<�ڕ�.���=Ŝ��
QX��8�/�1\>�M��O2��B����Z�k�x��F��r~.�9	�	�E9B�~�˝� ��
_�A��i�����py���#��0�8�����W�e>ŗx�{}vh;�c9ѐ i�+\�?���M��Y���@��7~��a����� ��XL�(`�&�/b�z�'��wӣ�_�G���cH��0��:�
��8�z���8�q��[M�2!�����XT,��o>n��א�Wtx���e8�φ�z)���j9��-�"c~* u�,63�߱��[�h�qߵ�g�kM0�ُ��/		�~f� ��VG�<���lw�j��E�ۤ-�U�P��j�!�����|'X�$��V��ҡ'	V�/쐼M ��v��v{�Bo�%�D�GI����Џ����byWǪ}���tSM����F`��Y�� �za7�H���n�d����$Px�~��_�G�|�O!v ��������#6©C�Y73�k�Ƃ>l�ke{�Q]s��.���vBU��8��Ί�}��/�~q����P�)��[/�����~vƯi�L��ں&::m&������)�)￩�f߳�q�����95��\K�F8�$�%�7����N4@�v��u<GXq��(d�<�cgd��[j���@�Y<������u��/��u��|��Y��'��`PE�k<�-EV)C�t(GY�8��	Dn��݃�"<�����:
ނ��V^D���C=�C/�YݭdD���w�Y��;�iַ�j0�7�Q�!����G[��5]D�4�}�{��t�CQ��l��S�/��/D��Ycم�0FZP��c�[���ޫֲ�lB�Nf�ft�wԲ��o�բq/�#����8�n@���ZN�/����KIV��+�J�ƻ�4Տ:2�m��j����-i�3�q!Hm��:�.,b�	��c��d�lŏ%� ��Y�P �r�낝~2�:�Y ��	�����	����-����A�`���Ԥ h�qԋ���k�GZEU�%�}z��7��l<`݇����4dg�SH�7}�h3i|rV�0�K���A���&墏�C �e�aλ����9m٨��tK廴���kq(�΂�d" ��6ݺ"UMۦl���I����j���{Fc^�����ǟ�1���R��lB��7u W��~���=�T�,﬎���PBg��V�&�z�̨��	3:� (B�Y��`-t�Rr��	�Bg�Mk���l	�"'`��sM�k�W�Y�F��ei�⧑���3�L�^���΄&� T�#������G�B�}��jAZ]!T�!EB�.o�
\c�QtKbq�J.�S��߬TX��=%O���z�a?�m��]�ʋ��@_�Ml>B�
�3h� 5g�y���-��ǩv$�r�h��}����gkݼO��_�?�����`�/�������CX/�7;?C� ��?�	��E���x�Ĕ�/^YX@�:z����ǯ,�r������b�Y��o���^��>M=����&K;�
�"�d���$q��?��D�o&z����!ذL�������)hLTlZ�~��؊�T�� ���֠��M�T�m#�~=YՍ���6Ћػ�|˳n�Z֑�P�{ǉ� ҟ�òğ���ˋ�Y���� ��F���*�Vv����d2n:k���aj��2�tKq)��# ��O����R4�ǒՎxhX)8=�
<��`+��!�e+],H�6�'���:��n>XQ��j�zȲ\�4)�C/S�;��!�n�w|�@�)��e�3ɗߞ�M��\-Q,�`�ݿ�w&��R�OX����J@H�� P_�֍sG��e����[+p�����3�����Á?Y�&����n�G�q�����\��i�k�Tl �cTi�j�������O�N�+ۉjf
��B�͑�"�J�L���"щN�r%&��&�Τ��讽�tq�ه>f���ڶL��1x�9S(k�&7�"��ECS�w/��J�G�ц���l{�;t���T�PO���r|L���+H��B0Z��1���:��o�@�a�9e���'��E*��W�",��Dm�1�l���9���g��3�c��	�m)B1|^52��H��[s�oh;-�ctI���� ����7x��B$ܱ����7PX���:���B��k���_����D(�,9�����r�p�a��l�ܠ���рc��.�4B�ao���$�}�6��>�X�24��F'���%��UI�b�<�L8�;�mRW��A�v˱3�x���)����H3�@��D욨($~�_+��f��cn�v6e��w�S�`B�����3��`J�ZmF֭J��yK�����u�3��<D����hQi:���_����x��/t�|�"�������_)|�w2��U��9�,TH��F�ZL)�qRw:f9�K���A�����KE�[%-��ddqM���=�u���4�G���֎����.��ZC0�ß�Waz��X�Y2js^�<����C�M��GU��0u�������܊�8ֳ��3���i���h��۽�%e�g��^c��#�Nty�Uw��+�D��>�>�;���S2���-}e�0�6���5��BI����һ�1�s)g��d�&N۱�^�f�/?�?H��t�>Ll>�t�b#��J�0�l䭳�����񡉙HXf���{��L5'�$%=K�`�F3��t�֛�QpE\h�w���v�̻ �z+�$_o�)��FM`:�V�cC���H� ;Ɲ*yG�s��eЅip�lN�~�ib��:�|ڑ(<��$�&�N��Z�G��b���yi�u�zF��)0�eE��55�U:$  -�9��K���Nr��$>TS�����$7��f����Y-�<��=�mRa��]AyPIR��ş�Z���q�^���S+ӌ}3�#��.ee����T��A�]�KܷD�d=�Sa{��4�m��"�}m0&�g��1u���Yͭ�"��}hE��~0��;[S���9U���m%5�f�W�!3R� C��l�����&&3ȅ.�+kH�*O񮴜���2�%�c������6M{���������Z��[��1�E�;�K�e"��
���:fT�)ӵ������^kt�@������K|v[veBf>�G�[�vr9��N̭A��	$2T�݉�V��R�f� �m��8T"j���_���7�,�q�*�r�:ɻ1�Ya�j����m�d�n�䂔~�&^t��l�5 f��/��rv�&9�QL.��t��t�0 �Z|�8��E��uV���i�����L=�0�N4�o���~���q?_�|Ƌ���Tt��Mt�95�'u�@�&qd�i/��~���p�����x�"[CL71Z%�N�ڴzQ��C7�u���'� L�u�p:��G99��^x��D�g�9�y;	�x��F�ֶ���1ƛ�*��G�jVv��h��N���6������c}M=��b�#=��5�WI*\A��4�+��4��]�L̴�����zW�R�����#��1Xd;aɕD�wZ� xi�����P�a}����������GL��_`�*f{Q�t�C��˳/��tg�h
�ѐ��s�Yb���䢴��pk&`��G
$��S�KK�n���[�S�'��\��O��։��d$?���\��47qaM����z�*���-MO��n)syX�����)�\X�2"4�̈m΅ ���p;4���	��V�W�O^���Q����$��e�LJ�UWZ"���P�Xևt4w@8�y�ɲ�g�x����>9:��W����EJ�bݪqm��R�	���wHo����ᐋh�,M���`Ja<Mq��������4d�t[��쵋���SEM~��zs͇s=�[`��_�@f�?���B���#�����?�L婈b	,,JyM+������!�|O;p'�3�U�ѵcE�ur��9���.�Km����ؚ��I1��o�|,�Q�����zw�Ώ@���T*\~%���L��c>�o;��_�fE3�i1�����9Q~`72��64����Z�.���ӿr�2c�j#�n�����]ܬ߸��jLˡ�ʱ��}�Әw�f���]q˱�Sc��7!��KѭE��.�@�nc��F���G��4Lա��E@�EA��D!]m�����l��z§u.�p] C&�u\)�4�I㡺����Y�S�}�͜wS+�2��(A�_q�W��0:d>o���_�8��ܒ��8�K���ݠ���8;oZ��+�T��*1���bͿ����ӕ9i@�1^����Γ�����h5;1B
Y��|]���H:�
m]]1e�l������p_Q�'��%9��.s%U�d�m
S1W�z��1�j`C
6�9����І���V���b�a_�a��O��4o�O���)^��Pp�Х��yܖr52�+T��_�S=O��U�y�j��y����tjO�X
�`����O�93Z})w���FBxB���c�G����X��a���N>�J`�'� ���R B������(ݝ��%Im"f�
R���h]�Ʌ�G�V%��t�Z/T(A=n���:+��fg�t�x�m؞�\i^�
�<�b]�ae	l�&ˣ��c�.�ʻ�h.�L��CX���pX�^��y�������Ụ�_-d�`F����k,2�)S'�����8�f��ڐb(vV/ !��*�@Bz-W���#�#c"����>ǹ)�>���Tj�6*�~"������GU����j�c>�_���jw�2�8��g0h�-]F$�H���:S�8�y0�T�E�*;��}��2e0��߫(��f
K5[�<�6׭^s�/�}�qb D�$�C�����g�W4(�����=���C��Rw�NF-�)����O��v�#��߉��׊��Gzu������!�w�_�C'�4r�1��� ��s�k�� ^u��'w4��V��ar�j�l[r�(.�㠶���x �XSj��X� ��2l`��e��O�z�Q�s���T�INw�nU%�Ф�=�wŧ�h��+�e��C���{�ɹV��wŻ
�9C=�� L;��e
��_��g�#�l�
�e&��Y�'Rs�_x4�V�������ZI�y�=����O�3-��eˤ���;T�ȣ+�V� �!q��M�8�^�v.��vpΊY��Z�A�a%5
N����Bu�rΌ��s2��JqH�B�8��]�-�Ba�71wf�~!�U��t�(&$�l*=���|޶��^g�IoLD�*�
�Aϱbd��XZ�&z����T?���5فv�v�{آ>�,���������dt�VU'� V�$��'D/�6�j��T� MmC��n�N�1�Ehv9��!)�V͙���S?&�Q�'���FT$�)Ń�)'�k$�$�D.��q�	y�p9�.�0U�EV�l2%�|��F�FO�8�^^j�jr�>��E*��f�O~'G��s�Ɣ}�Z~�L�w��Z���?TW���5�T�N��'�D�i�i��2�F�����
���X�Ꚍ8�Y�i��JQ�V��SA;n}��<F8��������O������СXt�x�w��䝆�����I��g��ȤT�;v6�A))��ް=�C�QwI'���[�*������q`�Ԛ�~��&,{@6kY�_B�S+�S�S�b����e�ѧ���'y��0@ل�j�*?H��\
'�)-���Ai�t�ؓR(�A�����1r��<��ੜ]g�޿���؍��ʭl�5�0	'e��`P��1DN�B�s��ip�-��۟��b�ة+w����o�P��?��it3_]��c�-Y���~0�����G�#�>���\kW�F�݁������@�>�$�\�/�A�I?�����''��}� 3
��L)(=�Jiv�w �9����7�Z��f-���G��>�냑.���*��X����Sk�&���� (*<ǖ*��]�tP�d���@��!���{��c]�l��	�g�T��Q�V�vPV<��%I��רMU���g�_��e���{5�ْ�Y����iW�r �����؉FD�ܦ7��1��@G�4��ų�ć'���o���9� �<t���1�N�Rp�,�fg#	Qb0�;8�~���,<�vg�R��'�7�����]������YT�<V�f�A���5��L�o*WI�E�ȣK�(�t�Qtb�-H�����P�AP��]�{+05���Oi,h2�}�������8b9U4�ǻ%rW�;�E ��u��ʻ)�ь�'H�-��>�+���v��ezwǝ��\J��)$"`��s'X����3I˿9r	e*-ҫ�b���|���҂�Ly�Y��K;Gʲ�J�3�twx�#V{�Ql%q(���ז��zW�7Vm�z��j��80C�\�I߰��?J�sj
���}Ndzk�?�e�;�(Q'e�R�"���0��:���2gW"g���29�7J��5+�u&�/Npǟ9����^(	P���~%˼��q���(�yQ`�K
k��*f�H�Λ���jb2;4��w�!���ȼp�����ς#����x /~j~��C��9V�$0}`߱ g��<���$�Y���6��ZzUé�3��Y�V_��k��^!��#Wg7�w�F.ô��則�^���t�dԙ�M�EY%a�=ot ��|
�ę�(�;��YG�<����O��n!�
��3�6h�'s���m�+�4�Y�\~��1*�j���2!s��2m�	�zƻ��yCn�sHGhmZD�5��#��Է����?d�$�^W!vD��� ��?9��h�|JOi�U�6E� ՍU��Ny�|*7\��QW5��~��Y<m�qLS*v�Ju[�4�����KN���#A�}��w��:A�m�}����/��o3�%j�S!�&s�-�:ip|$V�w5Yf�Q��X�D�@�D>.�S�Yx�v����Wz6m?�j����x�5�|�n$�u]mω:r�7B��w��[���F��ٖ0���d+������ �۸�,��mHz)�(q�F��L�QT� C,is�K>[a��dp��&1;�T�>\�p"�x����v��^�cҺ2���P�ƌQ�m8�T
��fZ�.B�>?4�R�����s��	o^�h�G�a�����\���O���kH�e�ҡ��a���eX�t�S�x���%높2ac�'�K����QmJ���ՃI�x�L���é���؈1�3� ��GAe���Z>�E��R���؎�K�l֬����B�C~���,����`��Գy��G�8g�l�i�����%���vA�u���q�"�ѫ�_Ф�{b�!��w�7�����<	�t6'�up���>Y��]�A�w�k
e
���+�x�U����gc�@Sy�m�P���/wk�-�����F�,�=su�s�D	!U��}zIB߹�A�NW�6{�y��r��[^##3�S��M�	EЪ�
�� �iM�.!��fJ��G����SM��G�0C7����_
*	\�`��ODҡS�w�����HNBM�¨�޸�A[��C���/x
�у�����m.� �.`du'�ۀl�|�8��xΘ�7��-xRK�_����� 	5#!"�@E)�����Rv���;>k�X��p�����X�}�B7[�[r�r��]�mwt��؎Қ�Bm�3����p�q��!7�8o<K+;P�6Pc���Jc_�Ҟ�u2���s9�5F���4��V�;HG[9����-5���7_�3i��6���K0څ�7'�>��i�+��6�v�Ҥ�ce{P�'��������Ɔ��ؠka/�����S'� |��;y����\˫3҄����,q����G��u��e^�w9+[,p�)q$gJ�txxizϰ��Q���^Ed������q��U�<�
-$%�ʥ�i�u�pɆ�<����Zju����������H��i���l·��V�?�����y!��������`��]'�-.%��д ��3��!jF�3�C�KG�<�����4����DMI��hOg� TlW��H�y����5p5����bݡoo�$RsH�_x����h��$��>0�����ެA
�?4�D�	ճ�v��&��|�R�����h^�&�)($��)�W�������f$�ۜ�w��eZ�?�.f������
߸��ڐ������H#ɚ���hB�{WkTq�Y�u������b�� ��㆛d}]f����g���ޝg�����`�~��:N홈'��	�I��@�@#� ���G��,g���tD�
K�Fl�?~"�0�7e�ͷ�\�W�x�[���~��@D0ٝ� �}�_�D�����-�F��x�e�FY�d0�С��#ݶ�8�!p��ô�
��w~]���h��i&������c��}@�:19@��K��;�T��:�	����Y�|�Y���zKa��˓����բ>��v.&�*����#�s�����E�'l�����&�6{���Wf#�\X�WBv-!���Χڇ��rr��ϰ�᭭��o?�+�_�l�S��F/�8[8�}�xI&�NU��/re
poX�p��M��N�Fa	�P�c�_�ǐF���W��x��~6�'ψ��K4�?b���~�(�3���$�S:5`gJ�?�My��ej�6mk���IJCT{$������T���1,x-�^�OZ2��z����'���G���k�u�.2�]�UE�v�=(��d�e�s��	_U6��$ϩ{bjd��AM	�Z�v���ݽ��Ut�^�a�Γ)%�Z1bT� H���"ͫ��VF3���Ơ?��9pU?�F6>�b��_i�=��^�{4*yUsH�l~���m��g��B60�MH�B4�ڰ<b��o�H�ޝ=l�	��L�{���.��ȉ�_�h�sD.�Me�&�o��M��GG�����?
���>���ra�\tU�n`wB%�	��msa�W��g��i4&o���f;�-:�Y��g�m<�"&��I�l�zEY* ��(v�@� �f������N�}�����19Oްp�i	c~f`��TpM8r�멗���a՗��D�� zĐo�R�icL��+B��ė����J��� ��:�Σ�6v5偈��n ѝV��p8��gk*�#Z�t9U�(_*�L=q:O��P���*g஘LÏ��K��W_��Y�]NܫZq#r����˖���v�����x��G=~dO."�4b� j/���$&�&�(�ۘ��}%�Ј����q�h�����2���!`�X�9K��w���7��!���5$C��cB�y �S-����L�X�9z���u��iR���S�}Z�䂼�~��^V��tm9�;�����[K5j��rV��Y�z�p%�h�g��48�~c��RK|� Û3�,���x}0�"N _�J>y�����z��
�h���c�̖<c��@>"8���Z<S��������W�۫��9>��۽�z���a�`�]���f�D4bR�Q��J���a0zਔv�}`�^I���BR��Y�#b��'���x"�V�yդTp�_OE�V*�H������k'�֮�:�U �(��J�1��`}g�}Z\4�"jɒ ��i�-Юkd3�[O�<���~�qM�_<�/kQ�}����}�k��;8M��ȇ��K�<���Qn�1ޤ������U����l�:ó2�1�j;�6;���V=��uV��˂ԗk㒓��d���t\**CDZ?�kK�����)tU�Og��&yzd��'�>�=��7���?)H��8~#S7ꛎU�\�d�?�N�/��M*�+n�7�P�NZA`iE�[fh�h3`�o� ���w���J��x��d� 85�a���Aŕj�YTɔ��/>w����n�/՞o�<S?2�1Xʰ��e��/�8�)["���ymbŵ�6���,���CF$Ճ�-ba���ȣ���N���o�v�U#Z䜾7�;:x�Pq ���k�@�=�`Qz��	Z�8���r�8�؛�Ug�ˠ�:�9�X�-!�*vv9�n��7+�7�&�*�Tx���*#�	p]$�iQ�����K���G��dH�o�ӫ��2i;�xvCNf�����@76l���e����\���C�v�~�e�8�������a�S��T���?9��,([j��� VE.6U����R5jZ�U�ݠ�FQ��y,���� �?N�vN�ϝ�@{H�i�n\�km��� (RK��`��4�r���ʛ��FQ[�)��Ɯއ^�ӏ*	oOB���zl�IH�{mvD�%�1駇��iD�����x�1�]��d�	f���+�0*
W���O�v*�b�(��j���{6�h�¼#|F�i�'K�"����`
�0p
*l@!�_�_fQ|�VC"��;�T��Y�T��V��6AG�ʬ��dFn���,B�2��)*��h��B
�w�  қ�oW�M����Wb��U�����ga�漥7c�cā�R0��i��2Ax�֮�}\�����Oݢ�����'=�Ahk*�9���Cɠ�֭��|z{d�E�e�#f
4�_r�C�)_׉Ե4�;�|�Td�����?I'xj���ԙ���Ն��$�����j���%^�hwB�ˠ� �Ζ��}���q��:G�&��t��`Q��晠�8��9AP<"����H��	r~8�M��{J��b� �t��
��.B�����P��SmK�-:Rj�մ�9�$�@�
]4u��`�Q��V��)cp�Y{/����6�8D�������@	kʳ��FC�7�C������wD��b϶�fL���6�/@D��,�;$��x=����qLe�qVg�q�����m��T�)��R��B�ފ�%�"�@�"��鉫�����(ځ��g�^�,�X��(a����Z���r�4oL\���N�Ȓ�B��hW_C ǐV8�x��~4&���N�C��L|+�R�,
Z��o;+��@�F�dP��>�$��6�ߢ���qz%��-J�k���Vr���/{R$�=0+X�E�бi�ȱ��x^j�`���6�*9����tD|���a�=JEY��A�sdvA�� �p�k��;��;�}����*D����$ w���A{�����o���g]��-��
��,�������I����'Y*�#��'���{X 5H�n�����W!����|0��������R1��2�j���ڶC⊦��	��k�xYPۘs^Y�y��Ot;0����(�����?O�w$c; /ڱ��~9tm�[���C�ŅL�9��-}Ʊ`�H���C��YG�{�f�U�KǬ|&Q��]�D+$L�I�����m��O����C��4��?�4��4�KZ~��䘳���3B'FZ�t('��P��i���/&����.�nGd�	B4���A��ܤU��zò3f倅(*��R!{�VF% :*��b�j���ڲ�
�]C0�Ǒ����Ii��N�z�7�Ģ��0b��Vʬ�BOTL��1�ImFz:#T��XN$n��D��ry��
E'��X��w��r����Y+˜�"ﬗ]Q�r;�-�C��D�h�7@�lp@L=�,�`9��X�UM�q��8<EHS�ٵ,�P$]����V[t���]_x���	�ƊV:]7R�L~��G�Ao��U�1*ocO�[ SrF�1(rM%NPA��, p���u�_7���g�zoKۅ��!��F�%�r�(���8����e�@�.��g���h�:.�m-�u�t�"��&���asZ�l; 8べg�wj��?���ٗAQEq���:������F~Y�6fW6�t��vY���a3��ۆ5|?\̩��:��',F|󘋢�ж�z�� {��C>ȫ�u�MTUm.����O}d<�Z|@�@�r�Ť���^C�����eiY�c�e��0˺���ןOY!�"��@������ �L����ƀ���+ 4�q�+���"\�P�w�|�z�""�pu��ӛxe��'�g��|H�Z�?����87����p��z��UN53��&�:
i9ʗp�&+���)n7�;�i���h���2W��[�>l�:���2 9j�ꗔhS�B�K�܈Ξ�?,0X;���B����¬��9	�+N��w��Md���Zs�]i|�[���?	����^ٹ�%{@����Q�<J�$�kpl;�Pi��S꜓ı��8sF���8 ;E����}0IMXڦd&|�_kY'���s��q�`1Oa�XO�kEm=<��I��ɵ:s��c6�F �����a+��a�����$�/���<��To�[������C�]���;Mg�]qQ�[:r�*�C�̈́ǧ��:�s"�RV%�`v�L�����������o�1(-���=b�1&����R� ���-,���#q\���_9��w��p�jC�H ��b8����zI3G����ϬYz�Չ�R�Ҽ�[fF��r�k�;Q��)r%��]�pn��Z�g�`�rR��e�7PJ<cÁ�y���S=�o�~-���\2W�/���"�N�*1��+��1G@��E��y�>r���'xhG�C�;�5�e�c]���︇:��}���#Ou+Zp�H�#�?���E�AJ��#�G���lx��`h5�x�d�m���� ��/�9��yŚ4��«;H�b�h�,����$�%���8��	S��nk��M,_��(�jO��w���z�ޞC\!�X@�ѭ��K��m1����3G3
���j,1��gǏ�j�;� q0\�����SQ�*�8�#�]��.�;0E� �%b~)5[-��Ē����F�K~F�O-̀9�eJ�s\� ��ON/1���o䣟�7d8P>��j����%+�` Ghsg�kG���(�%'��r%n5�@q�vo�J�m_��uy����t��"^����'����Ȭ|C��l�,ڰb\�q��Зq:_�Wu��*s9��7_�l�r	�$��'��SL�A�7��նZ$`�	��yZՆ���>��c�g�3z77_�+F���I^���[S����t����391�s-n�w:;�%��!*�k�*\a�ߪ��5�r$�{E������~�:nt�v�d�R�'����[����Ո<I����U�(�F1���"&E� o��SL�@v��l��T?�֕��$��k��,I��
�|b�$9��!��0s��R����׭���W������낸^l����Pz��t��v�
����`�zSݪ�g�&kW��K�$�{Y�)Q/�0ul#Z�L:+��N+��mp��<�<%ڄ�Q�R
&_�i �(�=;��,�7J%���K��=�M�@�g���%W��8����G�̌�H{\�G�><R��J"�G�N\��f�xqJ�G;�ҙ~r<���8[�|�ם���jAsڗ��G�P�_aˮ	�Rt`�Tc{p{�w&r�#.��G;��53���ٔ�ff�E�Hr�B��u6�h.j�F�㪻}������kuzvK���ȥX9j/�]�M-���Wx�����7k�DIuN^6Z����<K�)�5�t�A�#&�St&����D}X��%j,ZEk����g��[�r�Bq����k���`�G������jA-�=
��z"��/�I�t��Z�S=* f��0y$���<w����}n9yb����'ë��>�k�Լ%c
�!��z�������7�@�	{p�1q���fn��݉c�AF&�W��%"Q#9e��*w0^�'�AU�.,�	jϏ�sa{��!�F�;B�J�$��_ù3?"&4����9
K�����}�"r�L�H?gA�lUAJ��8ǟ����8���>zZ�v��΃���SU���v-~h�C�f?�W%	N<?!׵��e5����{�U�>�6��iT���@8])�:�h6�=�XI�_�-�"7"�i��|�
VM[�����R�9�D\����q��(�ahK��>���±B��x4�^ֈ�S��Y�hWd�<��J��*���խD��������S` ?�\����D3�u�W���Q%����k���߸�輗��Z������D�O��prN�G(�7��t�	m�4�BX"��@D2�A��ˠ3G�ã��ܪ���R�h8v�z�4I�ox�H����h)vEN
����5�^�������IH� <��-{�_�~�_���-�GK~�ݩq���'�0%{\�J!�)>�ϝrN
�t���ݤ��e�BA�M�B������t"q�}x�Ч��LJ��b�cR�0s�G,r��򩍇ۜ��;���j�Ix"Fa����Vy��)�����2+ˉ;%�$d�)͋z����BtҀ[u��R��P�c����l][^��C���7/� ������B�����6�^_�o�'����XC�������̉��O/�=��ǓUϹ].�;u��!�?ˣ�4/q:����a.��.#4���/��dAσ�9��l*D�
��C�8�F�����x���JAN�ߣ��L�*_�"�������k5'r�<�퍙-x��Gm�o^2%�F�ģi��Vɚnw���đ��j�σ=ِd7b��u����ɓ>�ԉj��]1d�\�M�ڽ��h����0�}�W+��{�Rڪi�=�m���<_hS�@a�I��D6�<��M�G�I��{��-��{�ċ"XuF�γ� tHxJ�ËҒ�Uq�46�ڠM��UG:�D��2B\�	�v�2���n��^*�vx�~�r7Qa���K!p'��%�u�C���F]�
co����Z�*����fT�9�-i?Oi�8�DYia�Mu>�Yz��: I6��q�vV��8W�'�Z��[���ay���Ӌ�m�Pu;�d$�%tql��I�0��p��ĵ��z_�? �}^�L�T�k��p!y����E �#r�fz�A�b�8�Jz�����4CV�'e�%h�N�i|�+٥��ȝ�?2>��|�]]��Q*{704�{a-"D¿�t��?W �]�Fd�p
�(6����4ݳ!ga��bZ|%.�'n�/<-�Bx��F\�?�����Ӈ?��n�U[b�����<4Ck��'��:��C�L�C����fAw<K��Lb�\(��<��YB�Z�r���{)d�����r���xn3 7�����o;�y8+@�	��_|�-A /�5R���3�_}�4)�n3䜘l������B˲W�b�*r�%�{����)1�4�?}��ѦȯD��z��wj�݄yL�����A5.��\ɩ��Mr7����TE��[�3�$�;=�b��+J2���]���	��:B�㎴|�jcʑ�K-�|0�b>?u��%��ꌣ�|��]����ϩ�Y��Z�����E]�^�u۵
������#A1/�5�2�+G)q{y�ϧ,��v�6j�̹�!<h�.�y���
��`�Ph�?�;��NU�<&�P?���eM�O�'&�V9�<�K.�u=�MN����[��x��-�MͽH�$U��IP��f���:CU����H�G��{����t��o�{$�ĥ3+����2^"���`5�����훮����yyu�UZSF�$C76�v���ƒԻ�~�K�\y\�u\^B"˩��ٯ'X�=�)W���O�h��r)ͅs_�d|�niڅ������X��4�%ܬr�p����ͅ��%�؄�-��0�"_�>d�$�f[��';�`�3z���C��F������9���*,�KM�
��0�p�%�i�$�TȒ��Q�y�~�<y���m��7Y56���������
h�!�� �����,��d�Ѡ������lr��b��P��j4ER4_��v9K[�J����N��ڟe&z��}2Y�)�r��<��X0��]4��o4�5�y�%e
�/���rXBi��p��A$!�@|<a 7u+������+M�֣��c�$� �ơ#jb�Υ7-i3���t%���rt��Q����^%vM@�Eٳ�?|�s��V
���A�V��:+��A\�V����%j�J�@�YC޷5�cv������̕j�T�>�;pM���,C��|ϗ�cY���]�3�#4�v*�җ���Ee�6~���B� �WW�N��,;��r�r�2pa���AM4fMo(}^�N�X�E['[U�ִ%52����Ve�<�_p�bR�ϭT=O�
%$���{�JdO-@eB,	)���ٮs::�c��3Da��7C�r��.��r���lGEEA����dw��j�v�rn��)����}?���v������K���s�M> �ϝ�Nˠ��-3I�sC�@$s*�X�*����R:��M-�M��o}�������]8���a5�D� �
����`_{��9��(@&A�&�z�)��7�[?Yh�#(a�=A�󅡱��?M)ᩕ�^6ٳ��v�W�D8�~d�/�3]�	P)~��q��E�/Y���O8��2�0)5u?%�:�~��W�^�ꖛ���E�D#Ն}v��� f�q���#}����4to�g����V櫥�1�+�j[ؙ�����G@[)y@(�����ox7D�	h�ޞ{�]��i�Vc��J6nIHz{�SJ�8Β6�LF���p�n�B����]�`��ԖI�0��;�_�<<����w�_� �z��h�_�� �v�D8��Z��,���/������h�n�|���<D�q�$��S�@��L��5R��Q�?��h=��-,��M�&�r�:��D��w#�0-
��>�k?Ǩ_K���Hu��]���k%^p�vdk���ODN���p\�(�H��/<n�3,�t�9m�*�[�� ]�r�Z��:�́�c���FO&���f���x �-	�N5�	xe4��&BcE9�DoEx8:5�|�z�j�}�O;����Md��n����.�p�ѵ#Z��U"�����r6
�%xNj�g~�+*�R�lN�
�4�iT1�""�UISˈ�9b79�Q ��H�{/Y��_gK�1q?�-#N�p�ޏ�e6�D���a�%H��"k��oC~�,��-]���ƄI��got�5�� EȆ>p�� }δ��+m�7�2�'䴵�>o��y�B�g����|�=L��h���5� ���+!��s[��N�&C�LR���%\�d�� ^���٧�6�~Hlh/�:_+��u�����Ͻ]tE��<NH�����ۗ��G�y���v��O�=�i��+�j]�a�A+(I7V[�m�Wt�Z�8����NA�8�$��n�a,���-:�6�IFyT;`$�hw߶�hNt�������DC(�aI48���.'�y{��+�W�0�g�Ӓ1�2�����rP32��c	Oq����Lc=����x�t��;Z~:t�!�d�F�7��c��k24D�S�w�(ȟ Rq��V3k='�o��;Y�/�>�2�=��lӱO��V�4T:z�:���;���,h��ԗ	Ub�]N.f��SB�þy��kC�oNG[9L�B1O�}i��k�50� �0?�Y�7��fU���󬃳��IEBɹ��ͅ�ã�oz��3}/�m�M��ʹ�J�B�l��s۫H�r�~����9�P�s�(#�$����S�MX��<���u��,���,B(-�r�y�^N�ڱ��%-}�N��m]�����)�#����>��BM*	�1��Ġ��6:��s:)E�����j��sWڧB�UtD[�#ߣ��R�Z����r2\�S�<v
1�Slu ˈ�fYI<�ѣ$�_,�uC��*�@U�.��Qq�F�5_�7+�m��,L:��r<%B��G�%W����E��x<��%�S�Ā7���{U����׸	C.P^a�Ӹ� �ۿ��gv)C�^�,���j �w�Rd���y;9���x�PD�V .P������6D�|o�X����l��"��n��� �>w ÐFRN͞��фؠE't��#��R�xv�P�ΨT�{��z��S5j�~�f\I:o�|
���u[��)�E���L���
B�#ELtȪ�g~��� �W#�N';8�D�	.�B�������r[�Q�S�u2ʼ��'�4K������)�&^�l��5Z?���L�~���fw�^Ԩ��U	92<���sX=���T�*�\�A�N�^d3ϔU��Թ��*��	!��\�໲ꊾY'Ǜ�ʆo/	;3�O+|�H�n����r���r�,��k��z�?1��f���wT�WT!���W�pU}��ԫJ�*��bD� Hf̵6�
��N����s՛��{�]+���X�v�A�o���UQNI�������w�<4=�摈������v���h�f��'���}k���>�(1�:)����8��p\K��㨇����c^�]����
>�� ����9 �o��6�'���D��<�Kh�;by�s"�T�l�4�.Д��?��o�B�	�<s�G�֙s�Qp�v��X��v`:{;�z#����oF�~��;���1eDOg�O�����-M���r�g��HuQ�Z�H���ڎV�'Zc7UM��y8NT�T�GaeLǯ���e@g��Q�Ip� ����fx���XyS������,w��g��rym}�:���vd�!EBtdV)O0.��O879H�JTOcȇ�j��	�ő����+I$b�Uʙ���򥍠_eU"���6���u��c��SvO�D4��SP�iu��bj�K/B��,_Z((�	 ^��KHر�� �C��>��.�+�OAjGMM;�X�L�eNs��{U�6o� M���AY[\��@#���r]P8�t��?��֟�/�c��î��V��;���@G��9ұ���:' k�uR-3!	Y˙�W��H�;\�S���D���r�+�
�rgo�c��H1�O5/�=d��!M�"������L���K�7!�1$���[���;p}�t��a����c��Yy.��+k�fqG����G86�ݡXa�{��~>~D6������U.�R�L	����g��"�g�g�����Yv=U+u�t�X�����U��n�#�VN��m=�㰶d�fm��6��c���t����w��rD�ðW=�fx��;���.�f�oE(�*�g~a���	�,����y!4�,��,����[	S��&}���VK�%�Hk)�{q��;ꪰ���,�LBo��xE⦞�j9��s��k���
eeH��(��q�����u��0��|@�'�9�;r��R(�]�e��p��e%`ON�̫wE�nhf�>$N+A�;�=��8���U7�
�:�N�T�0ʾ�����`ި�X����0o��}��\�\��Wv�J���~;N�3�ft�K��
����{]�(b>?FɬNjX�A��_����d���E�g
I��މ/qdr��5h0xm�py��-�4��RS��]	JE�ˠtJ�����)��}P4��FG�fe�EgҾQs�I�j�g�C�܋�a�*����b���5��	�>�R4�k��K���\R{#O��_��J�����6}�.k�c]X�t����_Q�5T��=���
D�PQQ6�T�c&i4G�Ҕ�P�ђ'!A�[��{X�B2B9k����
t)�;�ۚ7R�����ד,B��{�j!ښ��й+�	K)x��zY�Kg�[���Rx�'C	�fU.��:j�^�7�=KA���;]�
O���%tQ~�����8F��&n�v	x�����ء�<Q�׆Qཏ�*{{L���1�p�t+���`��"�+���MK�ze��p��l}[M;����6�xG�"BB�-o�����F��e�;dR_'���R�S�"��j�f���!�*�$y����毪d����J���ݒ���t?R9P���*�O��GI����/�q?�5�a�)7��A9�	D	�d?�4�GqvaU"t�p�ےw&���$�}�p��'M�����.�D|��/�vY����ZD��Y��);w��jrk��������?:�+ԂW ��NU�hdc�VSb~��m���"�8��:���T_-�	��b�ٿ��4�����sb}ձ�=Jf��vc+�z�-��\��)b�C��H�A�0q�f6�Xb�b�c�]�5�>�:� �	w�@�e!��7 �k%�$+�MJ��]����O��1����%��AMF������E�3⸩lg��B(L�2�m��Z�~����I�K��-�x�����>�׋^�N[$jH
u$B��� В���~��*����U�b����7��:���32넔{;m'[�m��;����L:'�v�x>�Fg��|rg��໮�w�=j����Ε}�
Rp`ʣi��������;C����r[t�=+Se햭ϔׄ$
���D�R�&�Å��G���cs�6�$ƍy?�mW�ğ=ѸIV�e N�������� d?+�7�(:�ѣ�M�����:�&���X b�L�o��^ڣh��"��FD�(m��� c�*��h�3>��@������]�Bd����.
�T��.���j)}�Q�!�����n{Jt�8�aݳ�j{��/��>�y�Y�6��n!����Bb��A��f_D�4İ��Nꑼ����zT�E�6��^u�����捶�)�-����z&�V~δ6nK��>@%�TS�n̫��*!���H���$ �J�:5K�:�$M�V�ݞ�ˀߕ����f�5qo-�-��TR] �ƽ �|��_�1�,����Y�AB��-y�Ԛ���N���n
�f3g6BL#�p'?��Mwc&���1��7+�d��'�Y�&E�Ҭ��X�p�tx�c;�J4-��٪*3�|��f�X��Q�*.(���+kTe�ܡ���x4��Dy0b����.��FO�
f�����6f�k�*<�-ĠM䑵��ٲ�%^2��!{����bەE���{|���� R�4�z���窉��TU��b�We�GN�sO-�Od24`�4�5H+�'e��P?šwr�[-����GB�V�ZXx^I|���)�I�t��CNw�3�yQ�S3������� ώR�+�qu�!@������Į���N�!JǮ�4Ѕh�	�����$ɫ����K,X~��)q��_1���:�wU�|���<�TKBC��pQ��&_p@��f���"sk�0�Μ,�����.��z�%��V����m�c��y*A���v)s�d��m|���#��gR�fHnh�6]�"ux��'$�1�d��H&� H^��������C����a�v�_�0��	/�6�6�AI��7,?'��;���6>e�b�p����i�5p~��ԉ����G�1��,ŧKF%��KV	W�(��(���D�dpVyr��LV:f��v���~�F�i�����v�)c_�}��_lp2+h���oԈ31�j�dҸ#�>��r��_6��������/^��0 ��^Ϩ2�K]Q۬���&�S������؏K�AkA����T�;�^�n#�D{�Q��-�W����T!`)���X�� =�V��8b�#A��-����	`�+\cLR��G�=o:J�wOV��da���T�ƌZW0p"�p�2�w��1,\GW�&�'`�B�����@e��/��Y��o�>���G'��.{���0Oi�ݼW]�"p�}� H��?P�{ӢFW�)ᓮSa�Ieւ��g�l\񻛑HupJP�>WC�P��y�?�G��GjK~���Ҡ`O�a�8�X���-��I	���U�ϭ�?���jz�g%��ٰ=7�_W�B�q[M����:��05�h����ؿ#�8yK����W�����M1B^�0�?t(w��g�:�o߶�V7��
5��V�no��4�)Dm/\�IO��ʒZ���>�W���:Я~�<��ߪ�t()�<��4�jx|ٖ�����R�\`��r�6���=�ש�=�-��sG��R;�|���2+Z��P&�2n�a8.H���5�o�R^r5�$�#��P�j4���Q�q�>�K2j��yclf�<�}Ԩ�-8z�բ5!�.��� v�Rm�e��"sFLo����k	����G&iH't N�NF��7��_��$�X��(f{ˌ�� �>��eUD�=񸔛��0={j��בb�찿I2=���N��h�C�����C*ɪ��Y�!l�#��7���t5��\�a7�Ϻ����^h�iY�ӿ ��K�[~�r��ЁBl��l�Ѳ�c@��ت-��恄&F�+�P�a|�_7�\>]�jd;ޥx]�N�h�v���Q��X�;��O�X���@� b&s��)�֟kFI��X��dE%�~���^�7f�A���9	H�7���X�1� �f����0zM�!teo������F��
���@���:�9�́p��&�����&`i��ԣ�G#D(j�o��ApY	�8w*�DEIX�kX��<�.��0Vۍ泹��Þ�(-�c��+X�ۋ�9�Ӎ9�kz�Z������7�+�Nې>ox�?�\�����]��(�A�vk}�������E6�#t4���=�c�VDb���0mz��Z����ɏ�7'�B�֟�0bYM`�,A���#́�|���0\�{��}U���l�-ܪ��|M��iiUb_L�s>o�=Z.�zr���P� |�g�jV}���ڌZu=i(#�_BL-o�{h�aD�ݗ����<<EV��T!�竸X�ݖ�*bb�n�+-�߭�ڭ�ܗ���i�c�o�0;\fgյ�!�>�Z(u�\<����5i]V�[I�	0={�c�TL�y����K�+6<n��k�.32�L��ҡIfc0;�k!��'��� _��1>p?>����yuƍ�:?�+#U�z�p�&0��W����_E��q�}��&__I�����IE�0-��̟�a92*���(C|�wU��:�F����LM�G_�UЧ$0`h�#H9��_⤰�K��2���!��4���&��J��'�}��FV�vl���귐~���{��, :��*�Dپ6�>�K�լ���RU���yx}b�Q���#��7���`%��7�40���L&O��4U�(��>ƈ�/Wح�6��l��c(�N�����)J������9B؆f���5_������8����.��h���q�4�7C�c9
����ʏY��ӵ/��ɉ�����G��1��2��╧���p
�iRh������ނEQ{M���/jlV�C�.��1��ǰyH;wѴw.x�c���9�s��Vt�a�t> b�P��h,��n*(�l��C�����r=U�}+-*�yW\qu���q�8�:}�f�G����R�����&L��;�붝�~
5�+y�Ś��9nni��֡�V�y�7Z\P5�v@���AO� �&�F����m���W�}�yQP��[�D�#A��l�O��)�(Рyo>y^��e���fn��y�<��Ʒn/�vڿ�D�������1v�"��7��4-04<灿�֮��2�]�,�"�`+$]i��3[%JҼ�����2��W�����Ik���$��;�a|rben���"��Dī���mc}�)�����f��E ����̏�"	�,���W	(���g�e��I���aJ�FW���%�G<�}i$�\	L� ���<=��S#l���$\�A�3Z��KhGQ��:7+�m=������h��h��r��_T�c>[�|��x�~!O���P�p(7)7R�[uc8���
��F��<uJ��z����%�q��dPa�.�B�@౱oceH/�BG�U9�
$"� ��&�����ؙ�܂#1��A������/�{�&�@y���=���-�&+�B�� V�5����~�d��_w�b�������w���!O�U5s����<;ߕ������^�X|	���%�A��Ŏs�������rA0�\�z2�u{�����T�Kn����:��Ú��hL6����)����MS`ˉSS91�_gx9i�A�h���㏲�:/�I���4����=U{��j�@��M�I���i��c�*q��:��S٬��ԙ��o��*�1{=-�:��1V�����
��1�j,^����_Փ��?�-�'�s,2����#�ΐd�Vo��.��F�2�' ��d󕄜a\���sYI�0^�i�����Y��3��=�C�n0��6f ��eLp�o��#im�^��؀�?�퉖/	.oo�n3#|^��L,����A{k���6�髣>P*/90��xC4���Z8{���(�J�]��G���Ml��d��bUF����/{�sZa����va�eD߬eá�Im�tT ��q�?T�'���� xm��c�ؠP�𫊇n]��c����`5HP~ｰ�<1����$T��{X�~��AV"7��Xft�+�`����Ȁg��GkPx{I�W~���}ll�JHϹJ����"���Y(���΂gq�(LN�B9l�ㅪ�#���t$:  _y"6��>4	^��D����rd�*��G�~g,�����ǳu]����c{��
�A�>O(�'����9�s�j�"u�V���6��It�� �;���Nk��� n�e�Wy��|
���+������Nש�MhL��So�p7A��7׏l��������( �O��˕����K���?4'�A��>OL��5���p�@a��]�n�=f��d
��v>��tA�BR{!y&�Q5���]ɞ���|�5Z9�Y;��a������rh��C1�O����KƌG�d�ȭ�:��U��ݵz�
���=l����t�Ɵ-��������pi���0���5�	�&q(�_?eF0Y�l���h�tf�U��T��Q;T�s0�#�j�+���i��]۽}ɩ��쮄E��Ðk����qݹ�� l��q˙5E�qH����?�N����"�*�8 ����ۼ ���:F��G��v�"C�k-2�U|�������i���;����<%?��w��P��?ǟ�x�����F-���.�H�oA�44�Z��\,�9��\�5%����]qۭih��+��el��H��v����]��8\�V�<1_r��;�RU�Eep1�gV)V�v�oF�Irl�z!BK��H~�>�\	!��,5��o��_[���҆bET�٣�������@�CT�|�v4�Met��C
�>�z����r�^$��ږ����}��Tf<rq�Ŗ�6�ku;W������_���5�>9�O��WSO�
ѣ���ɺ�hX)��:��[�TE�.r��Ps�wv&8�k�D�T�嗱G�	��~�پlzQs��7u�b�ͱ�%�ۙoRv���F�J�h�]���q���-��|��n��oZ��<�j3�Z,�Q��B�()���MʥH�����L$�sic�g�0Jݧ����K1'������3�@��7����~	G�f�NO��oQb��x�xT��ŧ�n��n(��-�,�Z#iL��� �1@V����dE"�maG�E��.vfCΘlRhq�7q��X.iH��Z{u"�V?+�T�&_?�����Cy~�E����c���7X�1��7�z�E�8���q��yV�.��C� �I�Ky�?rA^���TdL���-�5S2��A�3��R`]��m(n��KeEږB�����5Ь>��n��W�,	�(I[����~tʴ"��9�G;8��&d���4Qd!���G.e��N1��V:���W�L��^��'^m6�׊����;^W�4�]�6�"P��}��l�:�����	��Ms�Nm�m��]�'O�e������ ���n��G�#���%?I�`b��������zK
����ڙɶ62���N]P�ۇ�P�R5a�AAh0��`�{�_!�In|��Hܺj�;޿��L���]z�I
��1�yra�0���������cS���b� 5���0�#A��pX\ Ӷ��g6�zT���`���X�$�	��9�m-�����G� �F�����(k-�XhH��+�Ys6�PG��@'�Ң�xǑ�'L�Ԏ����i{K.��<�3Y�� �3ur�$1ʒ!��d�Tׅ-nA�c�
�E�z���E�n�H�xaF���7}�]���t�:h�l"� �쟺�Yȭْ!O�����bW��W�U����$�y�1(�΀x �9D�	��ɗ�1�p<!A"x`7��|6%��B[6�!�}(t���G)݇�p�9$��˨Z*��3߁�1m9�m��Pv*��O
z4���8��6�Lt�SrO��>��b�%+!�U������C�uOY3��(N1��4�n�`����fZ���+�?�wE��~fx�0�����$)�j�5�ż`܀璢m�Ɠ�*��$���K���$�S�i����o�3O:��Y���'���u��>f)ũ���S�E�z�fAi#�����2�!�B:%�TR��K�|�'�߹�K\��]A�yGX�Zs.�60e"��Ǉ����9����:.I�f>��� �NJ:���w�vÈ����m��A���5�w���2��"k]�ƌU�����YSX"���,�_��]��"AF1p�����y?���Q�W�9��!���([�i���m#�4k,t���(����T����,�{���ۢkK��gH�]����q<�s 7M!ua���'����(ޙ�<k��N&@�T�.�\�$xf������`v���F`)2�#U�f�
��Y���"��LJ+�P���蓻�'��+�8�����]�Rz�j�2|�Ï�|q�&��ۋӣzs7��K�Ǆ��]��CZ��M�S{<�wt��:��ΔQ��������� �� ��٥�
s0 ߧP��F����oV�a�tNyE��%�Mݙ��)-a�n4��
!�����M����t�U:����e'Y/_,�,�$�3��{a�$��[OgHqM��J$Y��G�X����+�W�e��<�ڿQ�"��>�E�m�R>鍰R4���`7�I�0�	�v�Q�f�Q�z!" �E�o����zԉ�M�-���)������4mOO<�Ŭ���1��1����#s5CՀ��c`]'®��d`	�.^/?,W癅ah���$G�=b�̜�,Os��N�ڽ�7gtf��VVc�����rIpl%���ϢQ�Q2q+v���4�5YֵP6�$*���9��
�r��O'zν�P��V�o�~��	�u��-sA������b�M����~30B��r�o����{u��5�L�3����g�<����� yC{�0�B���d0��rn*�V�����+��Cȱ�aS�����?r�؄^h�X���H8g�����~���R\�kՂ�r�Hh��x-�]�L���8����G�*�=.'9������W�~�Wd�
~mT(�����~���k>?er�Nm7��� ��R�#/����)x�PK,�!��EYvX߬ti��"��8�VA��;�cXU���R}�(ڧ1MJF����B�f�M�9'ܛ
��5��9��n�a�^���!�:]%¥�L��W���_I7���f�V I�N���l!RiS0��l�BEH:S��[���,�/B?�]:H��v��ŐE�b�F<�Q�����SU�_LG��䧲����SH�i�[���e��VǷD��)
�e���P�U�1�b�<�Vq^-�[u����;� �V�����"���˟c,4�%�ά��8�o��	�+*S�c��}�\nԥ�^�ڇTϓ����Uz��iI�f4�=14b��g��1=��������vt�+75婈��)6���؈NB*/�����l]2��r D��K�g���Z�ғ#5d�w˜p/&+1�Mx��׺�r�oh�����*Z�5�[�6ͻ�d:�|߷Fן�I<��8�_�oex4�|��
�M[�y���'���<7��C��.+~�z=�5��i}�k"�����%�kRK���l2�5����J�L��W����Ԁ~�2$+V�Dzj�V�2��8��#-i!�
�������	�tuТ|�\�����(�5i�ָ�GO�a��2 ;2�D�&��x�0f�ncH�Ԙ(�Zj�%��8�:|�H��/�z��K)���[�s��<aDRt���21��Ä[W���-���:]�#�'�I��V\ /��ET������;��ݶ�tK�!<*i���/$��S�^.�ɿ��jVy�d+y��hÃ��/BI㇋�
�	m�H��$Sִ����PL;�~twcq@d��a�b+)�hS����&�n���ip,�h7~o������^��(�l�m���ւ��tL��C�P���v�_1Z�'�u@���E�J���I9p�j��)Y���(I6[e�)�4��E�޺�~�_�Xʟ�y�S%���ۉ>��`jBiͶ�<���s�֕�Z4�χ	̥_�2	��P�A��G0����.�L�U��)����ǔ�m�k���/�4#C=
����U�5DNQ��w,�ա�M9}g<
�L(ィ�{��^ly��]���̇�;+mL$F�8��@�޲/��U�A�%�g��!�SI{�)v��y^��W�s˾�.�`XK�(��Ê��O����,��k�Ō8!r��ƶ��+�ۿ�/#����b
���/���Y�FC�Љ�U������l]~?D"��yO��_��ZHǨCWA�C��j˚%��m��H0=K[�8�d�_w�B����/�'�489�Q2�6$��q���&��M�N}�[��/%9�%�E�f�a��b��$lPN7�L�G�Ԗ�Ɂ�J��d"�8��f�C;��h�Ǵ�Ә�˩c�ҟP�a���@�z��E���a�1.�j��r���ږV�>/L����s�hݓ!��0�?{H���ė�.$ɺ�#9��G|>��m)@�J�j���x)����3*�z4&o�O>w��w����obـ��8�S�'Z;�6r�V���O7ѧ+!a���Xc[�5�R	/FUh�{�&�?�B��L��ҍP�)��;�7�����Eפ0�^�_�]g�T[���Ejp��(3��\�s���S�x���BY`�7������{OS!։İa�K�j�}γ�e���íd���aB���t�z�n�Ў:"����hr�8S~�>�>�ȟ]�Jq�W{��zA]��A�UU����^����${���Q�Qp_kM>�-"��w��F6�5�K�/o1`�����ydS���
�� ]ɟ>o*@l�f�do�����&�Z6�������=I����D�2���eN�h�"�4�n���S��:�47g�s���>�R����Blg<.J�cJ�+V��\��G%���P!O�� ��=��
��fa���FpA�g�q$��z�m�sH*��{k2�F�L8nE3S�L��F��^YE�e����Q=�,�G�c/�8Z����jW��5'5�?FN�֞�ww3Ԭ�=��q��0*�(r�q����g7#�Մ�wU��X����|y���HrA���k�lK�k�c���\�R!��ϖ�WϨ��&x�U�IW�'����~J���L;��(~o��Q�g��(2/�G�|eQ��pNkp���	ח+����NSA�ڞI5�)%ᐡ)���+���o���;��r��%�����&�BX2��K�����~�0M�]#���@�՗�߇V�(s��E��~k���i��)��!��^�	�)77R^��Öf��S}�~��O�]�5���pWb��p8�<�nVCG̒��k�-q����4�k�����Y��~C��b��$-����$�J��N�����fr/h���D��qlv����t'qxk����F�t��rƾ�|�ҙ������묖�Ѹf�h�D���ZNu#��o�Υ�4���E��iO/�X/V�ar��k�}	{r��������Q6�?�� ��n���� �X�u~)F��T���I
Aшo���rHX�_���d�NmM�Sn 4�����(i��׷j�kNbF#� e����e�:$�dg\Oӈ�~��9/q�h�[���Gu%���� d�`���
���Te�E�dI3L�E�R��o+0dH�3H�
4���?��cŉ� �m�;a/ԡ��8�vD�G�u�s�4��Y��j�^В�Iy@�YK:���P�dJ=t����`��]�r����k�m?)}!d��4T��̯���QeL9+�r(=���I�gx,'�jb�&���V	�d<�8\(�2�T�\iiSl�E���NFē��T��O�We�%�D��������	�E���5��Wζ�y-�'�`�ڠk}�`ȓ�M_��	�Vǃ�ˈN���i�X�ʫ2�m�����L�
���g�	i�͠W��.9&SG�b i�e�,��kuR��	�e�'	}N�tӏ�"�[a�����1k���w��9n�cpU`�b(Xc��,Xt�3�~���������1(�RJ�P��U���oJ��]�Xg.3�drM�}�Y�4��32�K�2*��f�$6�g�}4�� ������)����%�