��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������FuZa����cֿ���
R��U�����S3C�G�*{���c0�R�IG�b�`x��<H(�a��.��pVIJ���$NL]c��>/�lN��+փ���^�>W�7y�/�]���Dh��>�;�Zۇ��7��A��0�����4�!ub�0�ɑ� Y�
YY�����k=T��S���?��IZ�c �;��?`=��u�|�D��ul()>�,�ѥ�p�[)��;�cn�a_�ouNf��Z矟����E�
"�M��'e�c1M%s�t�[���9^Ύ�<럨܆�qA���x��\�8��v�4"�cG2����7�H
e�V�o]�J��4w�o^	J����"|=��گ�"�U�Ч��d�Ǝ��'a:i.26�v��@��@���{~{K
�1�9��OS�]٥S]F���N��+\vTt#P�J�P*T{
��oܾH¾p�~���|&�E(UV���O}\���{�4~P�P~��7D��v��Z���`�2��QD6@���E&)t���$r|�Sud�X[2�8/7"r�5UNG"�8Ǡ�o�q2Ӕ����"���b��uz���i,M,��D�MAk'�ƭF=3M-]d{��u���^7"��E2�����Zz�A�beio�ͽT�g���C����Q�����Rð��5A�@<�I�^f���af�/b�)�*}��LkC>˷�߸Ad'��]���*�i�C�2���^��z�1Ǜ�L���m\�Dl:4v&�5��m&�b��,«Ƭ�弃ڧ��3��s�d/���$WNc�¨�`�\�8/���K�<�؃�/��ʩj�,!%��8�y���I��W�H	���V̄L���Z�)�A<�b����H���?�3N<�f����ͨ��� -�YP������W���NOkZ��Z���F��������]�����3ĉq����W���j&J'����d�_(� ?[��`D"C�m�0C���x2��I���+��i��t$�����V����i$XT)�p�!/�N��B�̯.m�E�>���>+K{�ɦj�Vg�n���u.���6�/�QV��4��Ɲ���Mސ�US��{�|75t�id���z�t��%��*�Y�-���2@v�>�u�1#K>�-���X�ל���5p�"�C��f�#c	���<�G�����vcβ}�]��7��󳽤[BJ@�ҍ{�FbJp8/�Qfw�E������4=�}l ��QM�6-z��D�����^NH��˶F-F<٫S�a"���I��]��:S<P<Oq����K��l��� w%��Mͻ��`L�{�ڻB9�n<3�U��B�;�`�4��%�Z�mR�y���nXJ���s9V{���Č���~H�wR!�a�K�����ץ2��sҡn�����!�e��*ng�h}aw�1Lg-�($	����S����D�e?פWii���m�Zd�{�+aF\����S�{T����^��9ch
vO�9�̀��z��[����նw+I��aY�	�W-��X,cb~M�k�s�g{�WL���p;��?)�=A�/F�I�s��"��mT1;��$h,_��e .���.-��k:Qq��QN��=�����\�8�Gx�u1 ="�(�o��!�]���rEwU��� �������-�E�UbZ�U�;�Cq��S��/�}ܹ�8���r%��P*�{˂Ġd��D2�uD��ȜP�.7�܇����nGT���s�7�c��;���3���c�P\h� q~h������:������y�%X���\do��g��Z�(�V	5���#7�
֞F+.�T;.:�g1��sy1�G��ʦ/���Wq;[��S�㓝������� �K� �{i,x/Ek��qB�o,�M�{]���u�5�{C-�.�O�3b��*/���$3)d�v@��N���gLV�+Ȕ���؂�1�:R��b�]��E=�|��Y�$~Yố��_$x�~����9��8g��!��c@0��E.�ixxz��]�N���	�����d|.+�(�5=���Q�(�I�������P;�6��kA���B���t_'4vˁ�ـv����3� �-/�l���: �_\��&2�!A��m-�
���!֐_�"��7K+E�r�����z��E]q��q:�c��C|�t 	���
����������A�%�A���7D�9&�Ǡ�uӕʔ'�{GAȺm�EJ@�r*�w��I�ؗ��7x�d����"��\��+,����5�Lړ+�*�G���B�v�5f5lm�Xc��o�kC�y�ˮ T�t�,Z|GBH���o��W\Nq7\�[��R�hFְٗ��ci����Xз�TBA�-�-{j�6�Ƞ� d�u���A�ߦ�Tnj�5V�{�86|��ʹ����`�ո���ۛv9�ب��ߐ�3�����G���[Z@?��X7It���h#l�{���-k��$؍o�8	�9����*����S���ѱ��ږm�@�	iJ6E����EJ�<{��D4�o�	.� �$����>����+�.�}���oְ(;��k0Ȅ~�bQ��;xÌ�����5)�a��Y @33�6`�n�,�f��̦wN�Nɺ�/�xkzS�qz���$�����V[e����"%l�w�Dі�8u�:e�p8����5[�Z�H��[X6r�������n��l��C��T�^)���ښC������7V��	ڂQ̼n��4ʡ�t`�O��ORX���M�!��!�C�P0�]cيN���&-4�V�Hؖ���D 3��
ت�g�ٵ(=�Rذ���/�+v��lY��֥�f+�}u�Z݊`�;�L�8���B���<����n���"o:ŷ�s��-
H|�ܯl�W�jSL��)X>�C��,��'����;NDgVY�b򁟾#W�z�L_E�>�+3�"Ӟ4i��������p.M$ݐo�d�L���Bd�;nc��ȶ�+����I��7�f|����|
�ݩf�/3�1����;��[�7�=�5	a{U�6�}nR6�u%�5����8��S�KF�`�(�$��H
��)�I�R \j�  ��6qY���zs�D5���r?���Xz9/�b�c��6*��У78Z���hh�&�nBa3�C�&��$1Ο�v0�������1`���@�J!��)���&N���]�$�h�tG��~� J����U���QO�����J���h6R��[_�.�k��lm~��Ѓ����c��ԑ��Q0��W�]���Jl��������#K�ݶߓ�����Sdr��
* �g���T�O�Ǣd誁��I��"�WI�Z�W��?��Ք�/N��~��W��CUj/b8)?�MM��F��TZ0���8f��4��w���AtQr���T�<CY��4)?���f�s��P����Ũg�S�j��ʾ�\��?q�P�,_���'�xlϿ�(M�H��x3���@��}��v����Q	>h`�2X���zD�6	�������iz���)���<9.��%������-��[RT2�f�bW�y���sK���O�\1O����Һ�ew�"Y���c�:E�3櫳�n�x��O�VO��o���X��g�Bj��e^+����ks	y_W��uۆ��}�~;������͟�@���&�kfb�U���visK�����'RT5�N_��N�w�{B�>`Yz�m"<jO�$��@8X62)�9�t�4ya��^J���.�5%"گ�!�_��b�rs�� �.T7~p��Z�P'��Rg�mmS�|���3�2u�+N󒽤��(@.��);�Y�V�\Z߁D���������(���͟��b
P�o�]]����5������-�p� µ�w����-�GO�e����o��3�L�� 8įź�.������G�J��νRw�B^4��(eE�K��. P�T��c���e�~`��	w�0�_&U�5�F`�v��Om�;8%�V6%�~]����s�������d��L�tcE���p,�y����ɕrۖ@�1u�;r��y����MN�hl_�`]��*쑪�w#Xt�QS�^P&�ڻ�`�B��5�� /aK���E1�+��;_�.ľB���Y2����^*�w�6�G�ʌ6��,����ʮ���8�(ؽc�GyzuK��D[�]�