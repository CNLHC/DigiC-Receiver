��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%��XخV����0�ļ����i�$���iQ�ıJds����'��?���Q����8M�� ���n��g��CC/��u�`~ՙ��v=�g��\��&6�t)�c6��0]�
��
DG�=e��{�3���|񵭛� �4K���Ż��J5���)͂�/y7Ji���@ 1B�
���@���	��M%�y��>-H-���OB��[s9ڑ�#�`�h�!0M���B��(`���ˏ>���<P�d�/)�ަ'F#���~�hl������n��4tNDz���v�����\Gh�LaVR��:�c�ߦب&�7�c��U��IqN��+�(�
4L��S�хgL��S-^���$ׂ����I�+r6u��[�Jպ4i�T��fG
JQ]я�8ݰ}N�OG)?�Qh"�c�h#��W
�{�����Ĺ 0�N�FD��c�  �\F	?��o%wi�I}��Q(��<u^g���@��δ�[����k��ޥ����I�q,H���W�j��Y�e������V��z#$p:gR�h��E�U_���Jl�N�n�*ї�j 7�P�W��'zZ� �4~��4��5O���N?T�9T�<��D���*����x� }��G�ig�=~R~JEU�u��� ��ɾ��}���h@]H��Ł�����Ⱥ�4I�ɉ��l�.�J�qj�>�*	=LǗ6E{��\��]���`p@�G�it�'��ȣg�k�J���o��>�Iӧ�'�%o_x����[p�˗j-|��k�������5��C¬��ë@`�M#@Y��c؞J�fM�����K7���\8�\�f$�~���/�����	�5��8K��	/���--%�V�BT[�27
t�c�"���, �w�d0�>��L,�C���b"�f ���J�b)RO���������9�)?���q!����Ͳ���oro�T�L�黗۴�g}�>��y�'��ҟ`?�9���a�֨��k_ﻞ�۳冇���M�ѐ�Ed��f_gv!L�~`,�vYJ��{�9"R>�(1��(��bQ��݊X,a��{T`��Ը�o�׵�ʲ9V#��a��Ȼ�0��l ,� Y�Eʦ'��������<�|"w��Y�!_m|7�쪾W�������t��3�n>�͓��|m�}���=N3�q���6V¥�$����:<h�E3�ViS+���ƒ�d`:n��-���]Y�B%kW��&��̫4�whs�|L�f+�=�֜�ģ��_�ȗ���f+=H����k���v�T��:��I%��&B���h��8H)4�� |>i�'�#��z?D�u��]���K��h�֕!�bq�H
�,���bw&�9��!���cL�QJ4W �>a'��+��X��� �E0|��!Lf��E��<EJ�n#�����V�fK̰-9BN�*~g�r�����
���6�ʳD��J�#7��8����u��\lrb��Di�x�c��qO�g�&��J]Ź��Q������d���5B���v��\��`ӷ^[s�9!Ŕ[L�U��]nED�v	�$g�P�槺�U��db��G��t+l�x����6��݇�|���Sp����q*T�&!Is���z�+!�	ѩ
�-ZW��N����S*� )�ɴaw��`��'2Vi��:����Y�X���%�.��T,��k�v��KR"�tw�W5���ҹ�6N�����@�];�����h�J����ń�H�&�ISv��m�G3���0e՞�%�js�������uk=!I��R���
j���Lj�����<!d���4z�v�d��)7`a��˔��ڧ�:x�K��w��&�T�*�.�P�i!M?���R�R�r�
/;_z�F�s��V�{;���	7�5*I7pwLÇ+i ��b��{��/�h��� k�l"�x��4U/�����H	G���'�J��M����Lw$�h��p9:"�W��A�m�*��"ï�:��a 7Zl��:�l�.�T���0�N_��0���eP{i����l��^t-b�C�]���}sm\*FІ��ģEI-t�L���w)RҔb�M�K4l���;���R�[L��\����x%��;��ZޚjYL��@0��q���	8��Y����3CǄ��<�j�"RvE�_��<#Չ��ɗ��O�dWqd�I�(��-�D31��Z��fS�a�&0�j#]Yh���fը���In Kw57�F5^��5S�!��ލ)�ğ�X�4�ʔ@���&1K��y&]1:�D����w�ӠB����W�K��2����#��K��.mZ��ߛ8sN=���#�`_�g9s�q%���Uan�i���F��ѧ�Rd
Ei����ueiv�1���Ә�%QN�����mh8>�l�>��T����dJ`�e�m��
���'4��zꦼI���
�
a����$�.�S���t>*]�_��\��A�D��+,�)���G9����Q- M�q�,POl��FV�,5q�K,3�Y���m`n�4��N���jCm⨰s�e6�en� 	5IV%n�� x����G�_-�\r���A+��oڙ#/�����D����i�iO{�,�3	:1+X�����|���-����%.=��u��X��NU�89_&+D�&,ڲ!Cb�f!A
Z8�K�ϖTH���h�9�׶�6�8��1ĭ��qm��2�Uf�w{X�S��5�0l��=˸��a�\�k���k�76�'P:��}�f�ì�a(�-*	
g�M&��L�j����1���>�Hl���¤��*��,?�y��#7��
�7 R^h��Um&�����+��n0ʧ��������r!���e��V��AO�?��@��m�0}#G�_�;S�eڐ�)��^�Fv6��ÂM�9���~#��M&�m��v���G�cO'�=��צS���K��!	.�� �G�8��AK�������Od�Qr-4��%<�Б>f/Vd�K����T�1�6���ɢpzǍhdF���=��\��$�01�L�@C|my�������͟��2iw�	[�,w-�<�c�����4�X��1j��=����F���0����fAJV?�G�E�{?����z�Nzk����L��'��h�1��űS��`�u�̞k�jZ�1�4n���������*;xv�BP%џdI�ø��y�y6	S�"6yX�*Ciי���խ��
�c�H� _I<L�$����G	g�F���m@Z��y��ɜ1����̝	Gҿ�/�MG[��)*��)s7�K���	�S�UF������k5F���a���vz�%[�4�.��r�����HR�0�����������?�?����h�z��@��
�U0q��,Z������[��ⴍ��>�2A&��ǂ6�Xh�3���Q�����O��65)|����Ia���a�����9�E�'��l��57T�r��>����qT�#LDқ4/��r+v�.Q���L=z"p�<�pQ{?�z@�j��b�9��уf�ye���w�J�wߗ�}��&�����]9�ȩ�������=�J�)U쪍�T
��j���HX]0�[l��e��Ux��eL��^&����@O�N#wm�c�ӣ��sd��t�x"A�b/��#��aE����m�?P-����^��U����v���ql�����r��IP∞��	����e���a�>���oIy<R����o�����WA#�i��5i���p]���PH��b&�+�)�0�O���F$!c�I�b������١'��b �]��5/@dN��(Ȟ�a��
�$8VA���w�|���ݱ�C80�kLYg��QSz�,��bM���56�u�����<\��w����ѿp~���2�R��n`���dX��3`�Q�Z��/r�Ə�K�{��XV�AW���~D��\}��Sj���U��j�D�0�hfQ���y��K���k�ev�:����_���9�M��@F��0���w���Y8��zꖦ'�}��c�e��d�v<׹��gB��6�JB���2?ii�ƺy�rԐ�_1�W��
,�c:k��
煥7_H�&�,��E�1l_�.k�M�.���1&9])�8���}^"�ɯ	�Ng��o~�K�Z=�EO���TL��w�5�	�����A����BV�[��~�w�%DX�-4����A���hk;:�p���־�#��	��\o�f��םŢk�
�0�cQ�󎐋{��R��Ė&;rU�7�yTz!��_R�=����s4���1H�_X�_�������� ���U��84?Վg(nH���]��W-Kpa���C8�K(u�&�Y#�e�2w{�W2����]G�sJ�|�t�L~�������־�ܖa��UL��!̫z����;.pf)ik�bE�c����6V���Z<����9y�] �&(8����`��Sv�υ� �[�F��@��Ƨ���ʄ�G�~�{�KS.��#W8Ӝ���+�џ�Mn��xz�c`33)�_�F{^��<����|��UG� �yŸ�s�.��.oHzX4��7�x���sߘ�C݌M$~Y�_5u�	�r�`Y6~�i|�>3}���G�$^�r#tq��|���n9A�g�n'Hy����b	�о;���|��;�����Hes�-nv���h LE�.�Ӽ܋��>5�
ݶ@��Q兖�:��� ?.㩱�\� �n2���)�J\�C���]S60��@���x8�z�,��ťL�
���T��lᵁ�M�)�9H�5�9��ߜZ}�%ZkQ*n&x�����Cƕq��͈�W,�`]a�BIX�r�#��DlD=Lutmu�+�i#&�i<֔�ϔL��R������3��PE�?�T����\�X6y��;���F*��U�Q8k�M�+ 0��@��\XJ_g`�V�f%o�re�X�Q��H�����/���^�ɪ䶎�V.��pD�����u9�9X́�_�|���f��\
$��țӞ����^|��TtUͱ�ǖ�\櫈0+q[�zI'S�� #�������V~"4-m�y��R��dZ늿�L30=�q��3��J6H�E���U�cMM?�4S Z��J1f��r>�D�!����G����.>��A��6+����˃���P;M��M/��_��Dfӈ�ۋ����Ch��&�$�!n]���S�ȆAb�K�5JM��V2���I-Ҧb"�$/-����\>m�茞\�@���x�Zh��j8���)ݽD���&�'���_Q�޽�%�;5�,���!]�1X�D�Ú�B�s^�#���PU�]1.6I4Jn�e�8���"�n�dAՀ�����F2�d}vၐF8R��r�`Ƽ:�����fٴ'����>����e�p{�����Zh�`���c>�-)ެ�8����sM����j����Em�ܶꆇ�^|H9KK��sZbE(�
2]3��jU�
m�_(�1�@��#x���jskQ�&Jl�|yI�O[g�ErD�N���%��Ƌg��ut�n�f�D��b����נ��j�>�pr[��n$�;��"�)��M3�<�P�Ҝ�n]�x�X	b����VS&+2��ef�it�)�E/�m(�$�.���|�@O�K��G�'5�K��t��*z|[�~�k��?L�^�������枽~$�N�6Y�B}��$v ;f�ФU��LHE�Q�Uz����!Cv��"&��&E��U ��AR����<	���=5�n6�8�U��
w�qА�4e{)ē�KE�3���W�.��/L��� ;D�!5��� ����y��h$��D������ڱ�/��V�L7�p_���~�ܪ!���ұ�e*�nc���l�-`q��ו���X.�,�9�R�=^���ƌ,8��(a��(�P"���-�Fy��R�;�:yE���Q����n�lz�uy��� e��}�;	���R`�"�GZ��wS>�ޡ��w�9x��T�=��4�-D fiF�3��u�C�^L>��h�^l���4��{jە����k�>u��������7�6�;d�{����[��G�r�&5P��< pO����ep4�gC�4�!���6�Р/h �oP�>˭̠a��F������f�5����(�]%���@cO�b�[rd�N�,ꞥZk��@�qSA�fv	<������0���`�=i���a��(��H���VJ"��/o��ը��Y;��+%��pP_n�,0��Y.��2*��2b��p��0	n��A�(V�� �������N�yUL�l�bq�Ӽ�j���g�v�҅(ǜ�]0c0<�:�omaS ���+����f�#e�8��A�����BwP�`��o����[�+0=J�)�����Ē6��s��W��O\Jw��R���F��6�����'����<S��U�f�#)�4��[g±��|}��Ǎ���^6R�]_//>��`	�K����J�l�������(�,�~0�N��7�Κ3	+��&�&l���q��7��_:��Q�;�cS'_:�YZ�r��YZ�SmLN7�1�?!����	I�LWd�E>��\�]��4���a�-����ڡ��n��SLy+��j�ċ�ŏ"�R��Фd�t�|	1�pM�ԟϴ09a�l�"y��f?S����#���I�U錪K�2�JcI3�ZKN*���.��"݄��ѵ
 w)��O�d�����CX�\[���=�V,wS���q]S'��<u�ADꝯT��4���������ͼ)R��R��P_������¡&@1�*}�2�q�
{RĊC��R�*�I�ӓ��$"ڳD5}�X�%���c+�	�#�!�9m#Y�	x�+:/�ྤ���X��)z�ơ6�Íp7c�(1��~f=LK�䶤�}�1c� 	�`�a�\�D8!���0�0�����Ǎ��r�'��/FE��HHJ	�@�ЍT��zh��w+��2`q������䋳=̤��XM�Į�V�h�*j��],,���H?T�!(.������,A�do���T,���s��l��Gɚӽd�;qC�h���H�+��
i�$	�TI��7�U�ظ::�����6t�r��F�X�9;gM�8}��k1�:������|v�	u��n���1��C��2�u�{*ޟυ"!3 8bBYׅ�г�Y���_�
j1�+���ex.�M �W�G&�3Uu��?��mC�[�7z��FG�y-E�^�Ⲍ���JK�4�/�Oř��7j�9'�I^n����5${yK��td	?���J���B��폣:���&E�%��6��w���h�\t"��3�����Y�-,�V���׆"��9���Gv3��G��I���1@�rM�d�Xw�Jg���%wp�}�o�u}��}*�?�PV�y�� Ϊ�~GRo"�=
Ç�N�Д�VC���P-���l����ʬQ�=�A}�|e1���4�q��q�6q*=~�_%JWjv���gġ�I($@��qX�m�Phh�,!��������n�# ��$�
���M