��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���5p������H�4�z�䉫,C�=�^JN������oԇ�)����gd��+��-3�:`��Gx�Xv��Sk��¬'�fI��)i~B��P��#?�����g��p(�����$�5�Rv�����}��.뻌�����(	|�I�;��3�CWw�ח3���a�8�i0�x�ʯ�McB�4_M��(���ӟ�oC�m��¾.�r@̭�-9kq���ah &kF��+��P_H�v��3��}`#W>�D�//Z��=ih1p��h��N�ۙ�o�_��Ϙ+&l���'v[Qq��,�����L0��}o'a���j8����]}�ʹ��ZdZ��Hڎ�	�yb��dL��Yٲ���00���o6ܒL�hC�g�����xO�Մ���ꦩ� 'ʌ ���)��x���1�Wl��p3܈�K����=�e6�dƇ��.	��r@����ms��J�x�%�B��'�%� �����ۑB�8�n?3zБ��f��"b���z�TrQ���ꅌq��Y�+�'tNrF��J�9¿2���Y��C���G���J� ���0�aqt���j�}�xK/őS�F,�P��R� ���#5��j�>�"��e]��5P��y�㿏zq`�����V\ �>�q[E��� f��uS���֋_��#*{��e�7�f���w<ȷ��ܻ�[��Q�]�Bȡ8`��5 ���1������"
$:�8+�k
sdAPT�K	�J�qS\�����6DˈT떒`qi��|�z�Y�� ���4��U��)��r+'�O;?V��L��#��jXnK�w������e�(�$Ah-Ϗ�"/���FX��e�NB����m��5"W�n=�ƥ"�2U�N=pLp� ��Lc��;��D/[^��qd������E�3���q%���N ��.�E�&�^��w�IVf��R����M��@1H�!�p���B�]	�m�,��Ȓ�S7�:K�XLǇ��O�T�4���r �iO���@a��]���.��m��j#;B�0�_���^�Ûx��_�tHǨ;�::p�B$�dr(��f����b>�����H���Z1�.��Q)��/��ȳҐ�txj���v����A�>yrL�?�_>�J�_J��+�Vi���D�1�i:�_��Bf�NQ�#������̈���2��^��ͤ�;� +�t�� _G����� L���T��B&�$DN��"薤�y�N�ԟ�[��� ;��F���&�"N�0=<�aT{LVL�',l�d��$�C��?���EkL�`݇:t^A�8�笛��76K�;79k#�����P<X<���/�DQx8?Q�q�I�ݮ�Y�7��l��#tF�mA˒/�99r�Xt~�sm�|�4��&h�P��H-\��sы�oQ�e�'�#�֯����(��rTT����R�����*E��ⱊ�hA�3ٚ����� ���;������$�c�;3��.����AEv���搧��NC�N�Mh�~�˚�s*|˛�K�Ց�jt)u�����"��ō�)aB=G���zK@��_
)*���]Z!^�a �Q�ae�4TM��� ������
��Tj������3�Q���5�զk:RS��� �/��E�Ć��<os�����x�0'@�D	D�0s\V
��"q^�;�n�"�2���+���MIwroq�}��.��Vz�����h�,W+bf������P�tg�i�-	B*��r�T�u[�pXL_;�����pj��u7D;��X>�M��z��O��ݞ1��bs	9G�A�y��|����x�:�P2S��mv�;[AٗZ/F�uƒ4JF��g��"����1�F��h���8��>?N�X~�:u_��ͫv��)�u�RF��G���О#�5�Հ5&761�P�:���.�T�9�=����uVV,�O�k+zRN�I��ׅ���Ap�V?o�hN��
��R����/�*TÍ9��n���R$��'1� ����#0�����Բ�"4���&E�5m�_���W*��0�%7��Ҝ�����s&G��2�k�V�P�4�dM"Q���d�8��01ê���J�l���y�,'�S���m��9sd�DLY���cl��_��{�x"�cUɱ�O1�v䖍�$�9+�%}}Z� à�����s�KAt�!�7�_	����hy�<�0 "��#^G6䨦�m�;rH|���!nƂ�~%��5�!���o���6V��ț=P����w˒�E��r�����T��{�?���9�0��4��5+G(T�Z�z9/E�RS�ғ�'���L����W��01�+M'_}^@����?�y�m(��koY��<u�����&v�Fn]�OqT����&��_de�hZoc;)��?�ܞ�y�e&x�@����C�c�-(։�S�֟���á��r1j��Y�
�a}�P�]�4�Z�Fi0�Չ��a	İ���KheЀ�&�'���x��=�z#l�yT�j��tE	D�5sPHì���)ez��a�u�-E�a����=�H�S�y(5�@xȹ5�M\��T��	� ޻�N�>2��k�G2+���)���>��bʍ7����@�mL�*�3w�
��݇�k����D��@iIW��R����N�\�o�*���j�Cآ��(�,��+ �w�Wxc��x�Dז�4w�d�o0h��F����JH;n�Pl�F��kJ*��"&Kj���@�e³��Q�����%|lӶ��(Xݴ�畳J��~�L�ƽ(���M�D�Wy���L�?�E��v���DA3����V�a�!���Px� Op�^�0RNI��8v�{ aj9�OLbm�����!�>�ޡe|���r��!�Ԋ�|�=Qc%���)� �
�(�5�}���A�zv/@�ͲR#�v('X�V�
/�9v��D��\�t}��U-TX�%M�'��3םuM�O�}��^��R��G�#�gV-�Mz+�- ��3��7�ƚ,�#�VfȘ���M�1aJ��}���6�2�[�#=�P���������)�i7�/|�R	�����5�e�IK���&0h�pC��,���"�c`Oc���v>t��D���\��0	 �X�^Z ��yP��$��#g�L;O9R�(v�ќ��h�r�X��6��4����c����K�넱F�L��f�Mm*�!z�V��
�K�����:Y�$�	~�*:��T)��ׯ���G��/�>;`�W{�e�f�3sƨ�ޏ��ܪgj��?ʴ�}
.�쾘q�K9y�}�7���d���y�����W8���(��^�+b���H��)�N'����D��2h9q�_�C��=�'�<傐�.�ǮF��X��ga���.~ Z����<@O�'��ֺ����55z� G�����U�P�:!p�#�i��%PT�-I�ր^%��f )�)��$L���@�4`x�$%�0KM�Ҙ�Z�h@\�����ze��Q�N.
�i�T�.��T���/��}�1h���8���DYj��Υa��B?d��.�pE4O�R�v���IrL��'�ZQy��[�U2�5O>�C�f����" ~��\���'�% 󛘶���a;���;޶{zqX��*a�N���q�K�f(4�_3xcb��g.~2`l�*oP6�%t6�@E,P9�s�h�d�°0&Ѯ=�1яG�\i�����y��}O����,��W؋1����Q
޵{��X&{F:�q=>�wU����+G�]����K׌7�'g����,X/��|���-�֣��َ��~�x��ͪw��)E�2Y���������3�����t,' �)ю�t�pb�4.�Z����Ò-wN�h��%��w���kð6k;8�K5��u������F�U�)�yU����l�1v.1)���t��	�TH��\�G^b�����o�7k`� �27������~]�Շ�3�O�m��P�9~�����<��S�@rv=�
���[�d�=��p����\�q##P9�z�~=QR1�5xV�B3+�u� tY��x�����Z�N����n�S*z����s������q�οf�ս���,T<����|�uC�_L����gS�Q�E��:�w����5�CV�y)ՙ�\��4�n��������ncɥ�#;�ءP�� �� �����B
2<U�?��C�����R��u�%)�/��a�	O������9V���7� _B� O�<��[W����>�\�,�<���z퓑��GV�j�U�ۺ�� ���\f�@,Gn�'iT���V�����&�Gd�M֚�(��F#��+�s�ʊvhA�<����P�M�s�����\�$۠*L�*j�2F73��,W q[���J�r����Z�A�L�׾���7n�RK,6��S;�G�8����a��9����g杙}��&Dd�)��uQ=t���w�.'Y�{�G�����U�m=�_M��A�킗QdpJD$H�!���mP��BE���(�:+�V�Z~&�X?��(�Pӆ� oj��~��f�,Ei���c�&0|�gѳ�����u�B��<H�E�kXJ����ե��Ws~��w��ԍ��n���T2�i�D�k0H�������hqI;�!����+�)��V��N�_fS�]�Eo9������zŶR9��*��n8�Ǚ�R��5�U*@�)�Y��gW����߱8R.C�z�K�Bl�\����jhy=��`�o���"b�x_b{�������١G�/)m���L�1R!�� ��w��n��a�zÊ0h��#q�/�Cy}�!b]s�S��^Ą|z1�~|`! \7O��е�k�ڊ��t�j�o!G\Ƶ�5�b��DׂM�cs����Zٔ*�̄��i��Z�S����N:[����7�]��4�jM�zAzHN�70�����J�Z���{9}��N����jeoΆ���f�]����<>���7�z�2�?P>�H���S �.i�]�^��l��%��y�����L�Af ������yS_��N7U�]:�q���B�O��A��E~�/����,)��ɤ�Zߡ��W�7��^���U�(9�n�R���dlK��r���o��@�9���/����g� J8���\�u�)��]p��)�W��'��-�\�<� ��y:���<�	�Y��x 7���!o|���=����+�C�O�R�/Ԁ�o����+�"���^�ƿ�^���Fǣ�V��W���iQ���i�t��V� )�+�B���6��uŦQ�$�E� ��|�A'����L|��RT].�\oV�Ƞ(S	��=�����?����eF2����p���\�������Pȝ�h0)�����릛?N��Y�B�(�{��!CԲ~�u��s(�OI�L���Y���f�u��
M}�(Zv��N~�;u�4����W_��	�����̸k��>��aLɹL���J��ll
]c}00�M���c��Wun�2��!����|�����m����s�IOx���A���!�����l�ƛ@���7�h\�S�+������%�f�cУ3�oh�X�|N�?�϶�I�.��d��D�w̓Kv�LCTi�O���h`ņ��T�$'5�$@*$ �W֤L�m��b�U�c�g���S�6�>��(���g�W�u柇n����]Q�<�����]@�ƽ��ź�3U�ψ���j��Z �T�s��ٜf�X�Y�:��'���ii������F��l�R��d���̫X>(%L������%���9G����'�9���G�����d-HZ�� ��/���R�U�ؿ-����f�kÞ�)-�L��FK�������&��Mxf\r�T�p.�?��n��/�q�V� z:acf[�k!;�R��Wр�+�tKA"�
���lSA�}�<�NT��$�����
r_�.D�Qi�z_�,�ݹO��-]�LȞ�f���7���|Jϫ�W�]�I���d}N~ME�4�{Xq��K��#m
O�Ȑcc�ߤ��Ĉ�`T����,oc�"_@�<ʪ��}%�K1�:�P���B�:��m�$���I����^�ŉVu1����M,�*$h�G��H��Bq�C���е������֪�a�n�$��?��� �a�3�e�t�Wh���@`8�t�&O��~��7�b����amh��q���PD�� s�FϣH+]�G-	��Gxa >�BT��>��w����;��J`5�c�7K��Fя�;��d9߭�.~uq��0zMܣPrQ/�M����|���U���R���� lD����7�5��D��}DG�Bg0���X~J	��6,��Fz` T�P&&�N$(�Dd�U;Y�Ζ�8k��I Z�W(��)�W�+7�g���j���~�X��|^�W�8$z�ʍ}Q���2w���sm�����yv�Ħ�y.�8%�:<�`�k+�E�<aw�� ���a��g�{Xq�p�4%�|R>k��p�K�L;��!�"H��?i1$,�x'�l�Z{��9�anD��j|�b奵N�
|Q�`��?��H6j��Q�.�e�	'��ol�Wz�6���et�1���,��b���������}*��?�����'i�����v���2��TP