��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ������
e�Ŗ�SPt:]���/nk�tf��d���p�H��p�*'�!KX�����u�o֨T!���a��7B��#��Li��j������.Vڒ�<U;�����|U£DM����X �f�Q�z�G&������dr�^#�0��Wby
�a�GWP�|�T{��(*~ț_�wmo܎��xS�LU�.��:Y�o����zu��탞m!f#,�1|���Z��ʸ������N�*��	����"�/��LgD�o@��E����>qQ���7����qs��R��|U��pN���Z^���G����IZ����$�}�]hA*	�
+��2NB}ﴀ�q{�H5m��adw���M=-J��ʞ�'��<���@C"�x��p�bK��<�Ũ:OQA1 �(f��Z�`��]� �k�M��kȉ5EA����5�Zv�F�fz�r��DPV�LtsI(��b�	����v"������]�3|f�Vo^�v�����p섶���![����m֕b����zES4��_M�HM�5�����ɡ����1.̸eH
��&02���1F0�,m&$&�Zk�-}+�����X'�`>��A�S��fxp�Dv<�ú����s&uԪ�(����i}/�A����U���K~:���;:럵��V����œ�M�dG�jՔ��r=�B�Y�R�8�ˆ���x�ƛ���>�,�T'Ei�ڐU8|#�1?�	Ed��k�����`\8l�ܓ�:3�R�i�����Nq�����u�/7#]- ��釞��4d��Ԃ��1��ާ쎷\lIC3�޼���U�U>��}���\JzȐ�J̑O=���^*m�~a�
�8�m�b��e!M�
���$���;D7_��.��O�_t�kaQ���Pˇ1�3�r��wx>C�� �nR�hnZH,���N2�bA���_���#|�=��LB.���U��̙q�p8��w��\:O�������)⌃$�$�7�R�tgC��:�D���XR����=zo�����:�
��@"�u���`y�������l���[�@��]�k�kS�����}��0��f�4�p�C�Ҡ�����`Y`�[1u���-��U&���o��K��/�=^
�<�m�����k�?w��W�N���,H���AR/HQ��[zD�٫�'}g�k%�hv�&i��s�]㥂>�c��)]��#!`� >�,�#�͙%*
�14w��+�+՚[V��F4��O���^���1���:��iw��F+|s
mK���{�>R3���J�d�^�e~�G<�P�l>��2�u(n�`t�E:q<?�>�r�+���PĲ���c]�vM��_��%O�����1y�m	�����֑���Ԋn��F<۠�ַ�-Qʌ���$�va�1p�dچ0����AhP�v:"�F�=��3��t3��O��~{��.���~���
���`5�ӏ'm[
tn�l�7	d�5���%,#�LB�q����ݵ�Y�6�s�@����o�*}�����Vhܿ�0<�`��U���٨^��4�8��G<�/������t��*(�"�^[r�R�{P�D�H�R2�D6�0K�|Ҽ��[GF��w>A/�{|�&�2.���	�i������d/O�?t������ �^�3RLUy�Oh^�L�MZ<���,A�m���ƞ�绶(b���u�e�����Zio�VO�$�a�ͅ}U�=P�y����IH��(��$$n�@*�h��uGR>�Ԇ(ۮ�D�*	��D}zL�V���|�(��/6�{���v�D�Z!� d<���IX���{��2����k���=�w3�b�s��?��yby�C3Ѣ�+�	�R�Uk�J��"�ˍ5��ψ�0V���4�B�HT&�G�H�ر�L��Ճe�	��}�^/�1�Lb�ꦈt.��պ��_|Rh���d��"�ގ��q�Y��EAJt�7g�M��D\����={�`G�4`A5��Vbj�kգ̌<�[�����߆$h�Bv_;�/C% ��N��b=>$�i> �� �0��mA����!^k�|�3�饿8n&�-�U��������'F�X�a�4aZ����_�q5j\H�^�:��)��s\�H�ڠ�6ҹ��/�������̺��%@��$oP����&C���VZ���z����8\���}9���#J-X��p�������}���������"�ȅ6\�Ґ������^��+6�Y$9���A��+AZf0i�w!SX֜�Ni�a�{�'�=[�C�f(@悗��_�>`�c�_�j#�9�yja��1��>�mh��7����W1�f�u�_������`l�)gM>��34V��	7�ɂ���o% ���Y�M��H:��ݢl� c��A�#��)�SqϠ���R ѻC�o%��?�Fz;�m?���V�3���L���#�����<�ʸ��ܯ9%�ԛ�;7��|�..eBA��B��Ä���.H�w�oОz��K=ݿ��c��h�wl��{{��5�g�
RЗ1>�'�?H�D��%��<��py:�tq�6�����³j=we1�	�k
������&�,ǹ�F���9��[f&�KU�K�-��ǆ���;��r��Rt.8$��Dip,A�x}�Un��``?l[G��n@�3�.���â�P�R���]�B���K8�r��X/���E��O�;�����a �nb�#���L��U��Ll���\n��-���Y�t�'��|]q��#=b��t�'�&g��jWt� y1���X`��R��4�aI7���� `�k��05�2Cd��!�;EAOW啪:h�Y���m?����c��,�P���ƁA�,V���ɸ�A^ݍ�v̑]�E���"<�106{�o�� �Yv�{WrY>C�4��+��'�F{.P�9�G��j��N�%A�S��EgUI�IL�7���0Q��N��uP�G�@�Ц	�-�����<h���c�0����}���7�8�g_G����b�૓����]ʥļ�0t�ē�GeA�:獓��l��l�Α�,��ɦ���&M@p{���L�Mʃ�w]�v��� B��s�=�7�x��L��x��BGX<��l��5:\y�7�y@�B"=k�v$���S��Ds��k23mI afa.I��%4v��L(��	ea~"M�#]uz�ƥ`|���-P!��fs
���-�����t��a�y�*����`D|�Ny�o�A�*�FM^Y�=�e �aV������G�s�|�i�z��nm��h&o:�v��Jw�C��FP���X�#BF�Bhmt�ڃ<V\��r���}�4�e�������~�+%Ӡ�S`A�9�g:@��U�O�{�"s��8N���}D�| ]��y֏���?#�Ed��m.\!�h��f#2P�6��@U�'C/L��(�E٦G���T��-��~���`w0��YW<S[�Ju��sp��rh�G�GؖJ�~�Զ:���5M�Ox`e(�X7�2�����l��*�#GOh~���Y.�#�qM{��� �Q�@���"Y������s�T��neP�!P������g�@qD��6�-�C��>򲞯|_����5lC��X��b�� '�R�o�V�Y��>�1����קM�w�k���>@Yu?�+0Dp��(����
�޷oX�V�km���?�G]��݆�p��ϳ�,@~#�C�' f���?��d)[���;�&��h>������C]� j�x8��O�៸�z*؋��_����\�A(���1���oթ�y��w�*���������j�vnX�z��F���_���R��,���d�����J�{c���ʓ��O<����F�a�q�QF��u#������TZm>w�M	�^$��g�.Na������=����s�?��{B�(P�5��Wx���-�s͐����0<�3��k�0Mw����(��<D��9�"�lNl��?�(x���y�c���AK&'
9�B�[����lr*~��ʗ�Rp�"�N:���O���� ��,#g����/�7ؤP�ڛ��
��#	)ȃk�G�'/�C�v�!ZA�B�����U�<v��W����6���Ǻa��C�?x��A�;1.#J����;����x2�?����ekL3��I=�)���J�C����k�-Tk�XMKw�&b��x�	V�g~��@� ̟Vr!���L�'���z͉	�I>'��HJ��ޛQ]��o%��=��'ԍ��@q�^������T�\{G8;�ْu�5��Ԍ��?Ԕ�0�Kr��K�LjEa����=�a����LW՛f:����9�^X�35��ȄR��S ��� ��.YZeA&���a�M������%֒�8��ٗ���n]�&��i�cKNd��z\+��x1o�)�@��
y"���FX�M�V0D'���P^�M� $6m�b&�l�"�̉f2�Y�����B�TN��[������L���9�Xy�Ћ��