��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]i��n��R|�u�2�vi܏����J{�p���ٛ�#DyYH��-��������[��4X�8m�8�e��Gg`�1�y[eA�*&��g�T[�y4���!�4��B_�j�A��y+;���4[��S������cL��jTz��op�D�&e��3Mtu_ �qᎇ9�~`_�ӑ=���mg��@�j��)1�zn�;��t׊߽�
g���^��[?�(���}"o��5Ս��T�`&0�5g��y������!�����t�>��L���1m�S�#Wt70tX��z^4Qw9�j�z-Լx9�E�L}a�5=6R��ϭ
��غ�����%ơ��g�l��=k&�d���A�e�^4s`T��*?����&N�;e�mˁ^c��&�;�xYx
(\oUr����XG�f��
K�:���:ܚ<rt��8��W�c��V�pצ����?:�����q�>��تz9��(Z�׋�'�D�!ybN �>ϑ
�����]�Z[��F�#+Z�D�|S��)�J�M����b���W���� 0M�%���g�]��Y��,{�Q2ka*`G�@�^>�+�	�+	�u�+�ߙކ���ϋ�M֛)T�s�6B~���/Y�%�.�B��eҢ�yVa��~I�{K��]�|�Ӎ��n̠��E�	��J����|X�k��1���iD+���
d�<NjL���Y}:(��v��D���ф:hjL��F �
Z[��5�@�]j�Q&��:��Z�9���xI2�6���\��
)4�X�w�g�_���������t�6�R��]H�y���X'� Ru)~���Qǆ#�f�$��!z%�����G2���>���`�@W�"
N1�JH���,e��y�]�Ӯ�����㞈!�֙�_,�+p^j9	l�E|�얼V�J�w&�I��5V��P��|�A2�v��`��s���od[a���|e����;������W tӗ����A�x��mw����\��n�C�k��A��
��� �:)ʎF��MNr=��%se��l*\E�qr{�XCQj�����Cd>�X��w5���O���
�]��h��Z�I�8�
Q۵A�$���d�'�\��iVl@:����7pis���Լ�P�F}H��s�.-�:I�-���j���HZ���
M쩁������Xd��޴�j�7WfY�B�.�����
���Uz~���!���i��}�m�yWȻw��+�>Ծf�,������|ݖ��&呸��&�q�\v��
Ӂs��������x'�K�w�e>é.� �C�u�G������gG���p�m-��^�m�işE����:pL�z�З��4^E���0���T�I��Y�?��Y%.�K`�^Q:�Y5�:
1��"�j���ʕ6Ȣ������Z�I�}�	��k�c�� L��!�S���g&�#/^7�R�I�U��ź�;R�o�$Yg�r�H-13���W��=���%o"�A|0*!�:h<���G��{+<ik��F�"�����:�1�")�=�l�u6���Lc�-\���-A	�g�;��r�/����a�J`/�E��5d%�پ0~_a��t���_fY��b�XjS T��#e=τ���#����ŷ�O�5�� ��_����7��w_Q�����͑�Ѥ�-9N��l��4�����Ѓ�p�/_>�Jc_	�tB$�Q|�"{�LmmP%���ݫ�p%!�$i�RV��YH��2��3�H�,1�Y�0�x�y�\צ_�fN::.z��N�R�i,���Bp|�5�Ͷ��˃��iP�_�>
���P7��ב��Q�i4�?V���PTDHC��6	��'���X���:	�ë�����2HǮ����U˫��%q�et5���P��E����[w��N��1;�^~2=uY��%�7��a����U�'��w�F7J���b?VCR+ؿ�-�h+���ӅbALA[Hl��R�Xo�#�%/�Vo�Æ���	ՙ�GcZ>ÞB��{%��<p��s ���C*��\���~�J��� ��&��� 쏤{
��P	�8ܖr�t�>8fJ{.
������*k�ۄ���