��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �'�(�٦����6M^� y�N&�hM��\�[ʘS���Z���)/r݇�?*x˯F4<2>����NM��o��E�/Y�tBR�S��j՝�ڕ�!</
]ٷ⟯%��%Dq484)�gL�A�)L��@!h�xr�m����y��4�QM�DG�!S$?oH��;f Vl^7LK��rC�W���r�-d\�!��Ռ딂��?��m�-5�I����'sȘ��q�Gs`����c��� :dk#V9K
�D#�n���s!�W�V�#�>��Z2�c˃�{��d�XS_2��z1�x7�ζh��S������I0���<���o�
��Q��)���aZ&�A����x��Qn��ଔ��*N/-1�<""'��J��n�%��g�*���%�&�1�T�'C��m���v�N���\���b`G�Z<����Q���(+����7eo�9ุ��*@/=�l!��^Mp2���:�I����Rx�ߝQ��I[d ��A"�i�>Ø��F��RM��_좵�����&%�([{��s(�	��7
o=�w���e�{�Ċ���H"g��Zu�7y've�)�)~�[�&�EW�e�;�ru���-Y9���To�L&���'(���c�"�|��U�M3�����᧤*P�-�Ea��2�~�����j�{��*Ɲd�A�Q���K8��c)؅���[
3	���ʵ
�j��y�Rc=���L�c�k5�ޥy (6���E����� q�0����g��_7�F7;�[<7����)~�2*�J�Hbwhx�������h�y���1�'j�&�sN\nt�b� ;�z_���r&�tNҲ�����.�
J��}�R|�+�G��R]�?h4�j��_nRfڵ�����d=ut�����Xl_�#�"*��G���BkxQ8o��^՗Tr�D��	����@�q Ɲ%�酏�� �hA{�w�������s�H�.A��7S�����p5 49��F>AJ�� Ì��J6�"���uu%5����
~��9�~��d#�6�[;%��p�x��Ld'��2����|f]���`�|��O<΋���,�'��i�
	H�Ah1������o�M)��54+�ڭ���AD�Y�����7��Jf�cub4*��-ĮC�}2[�L��%ǯE��g%L{�,�  �J�	�#��~�.������~������K����-d�g08evbJ�ܮ��@b�z�υ>C�l�/�ߢ�+n-�~�HO��]�2�/�8E`>�o+�+; ���cs��)��flw�M+��s44��Q�Yf�
RV���Je��ǌk��,uu���W��g$nw^pi9��I��f/{�m�u��3qQMjP腾F����2y�~���O⼐e8���3 �O���^�`���Nųp����*�\�t��8��̅�`�"FA�'�0������K��5&P���/wUȰ�Q[T�(�`�p��n���+i�o;���("��Y�%���V�� n���T�A�Z�,۔�Q��>�w��w	�HR�
_��T�0o�s]��V+�P�A����A�K"�Ҧ�R&�� ''���y��%i�fl�7��}F߀��;N��l���[m���.<o�J���'�;
�nl�1B��8����Uya�\��ֲ4�ko�u���+-ҭ���A)��#n���I�];ظ�$���S��B��v�iB6IT��B��8�p�jG��e*;���
�MN�*�b�����Gl�i+�푎2�.s����T��a!A�$w
߽�B��ܟA�-�~J��R��n:bK���my�N�����SJx�FW���>h����Gh�(�|��Pf��q�������	If갅�ߒڪRn�H�I����S��P�z�`�p.����ߩ�q̭JJ�G��4� �W9Ğ���:���^zqÚ�f]'~�B�F�#b��E���H����Ov5^�o<�مn�Ad+!A��f$޿k�5C7�巼~������x�N��S�c�)����[��
-�����"5��5Ϝ�.�\��W0I9=;��s�j��f꘯f���f��ؓ��z����K0e�C��$a���쥏cbe�`����+v��-�Y>�.���p$i��=h��TB�Ő���v�R����`"�·΂�F� ="���i�O`�x�g�1���}1�/��̱����Ƥ�k�aG�"3T�8a'���>�j*�\��؍><B	O�zR���:����]�P�M9������c�4<��rK�[��&����Prp7:&w�|�v��vZsx)�OB�c�Erly�y�o�?3�Jq�P�&�v5s�y�ȤT�O�ς��5�l�<�tQ����#��+x=��˿�i�_��{/a����D����=VX�e����p�}�P.���Ib�v�K���������(hϛ�g�x�����k>��X��C��,\�������y��� �����]
��_q��l��a���H���Q��L#��[1�bj���۠� ��kC��.�v��ċ�o�#�;�`��w�ex2\IM����#��S�
�_9��V�R�h���Bf�zbw,PR�-ʧᘴ��E���G}Z��~��ˍ�d�9���ED~��C)YP����wǜ��ҭ7�H�� �\�j�4SQ���`� �~�2�����"$��>8��l��z`+QLo�|@�|b�g&�RAt���;b�zsE���$bV�峹��B�ay �����	��DP���*(�4�ؘ� F"���O�?��d�`��3wK�k�8>վ��(�
w#և���31C��� �aW���.1�Z\<��З�GiF�E�֏�[�[��E�I�Z]^��[�)��k���^ ��4��9~�LUgł����Q�����l���e2�zD���j>-��E�����h���`zx7K��m5���P�o�QQ�,�{�C���)��?����2c�E�w(t��7T��K����ڭ�ܕ;�-�uA��;J�o~�0u�.��C����'|�����K�'���:���-� ׭,�6�pS����Q@�T%�������;R��ږ����j�K�Aٜ���)Șk]���4�4�zW��*����G������X��oT�����F"ozs���w<�A%�9�/��)<��l���T~����8�ĉ,�������%5�K��{]L�����#���V�T�������1!�x�+��n�><x���tϖQΠ�"��Wy?t�`=	1,3�@��e*��vVLh��
џ�~��p΋x׳8>�����Q��@G�pf��b��5���1��mm<�K	�=�BJT�<���zgT� ޞ��{Uʢ��ރd�����M�����Y�M�?�� wb�c��N�L{�	A�Uj	���A�Ԏ����E ��}r��ܬ�O���(��pv��͜�j���BL��ӳ���n7�c�!�>V���wАαS��_۹,Wm�hy�$ȵ��s.⌝�v$u�^`���%6�4���=\T�Տ3|�;�@�z-��q?�0�ݒ����V������Ssě�~K�~����q�G%� D?�j�p� �4��;��:�63�l����Q�W�D��E�����Gcǲ�F�X3.�ķ>^I�*+�/s~�iv�)}O�H�l<Rh28���c�Z)K��:)�bѴ�!&愘�WO�3�����Q�"�?/���pS��G ��0��q�k7�N}�)�<��W��Μ�#3_l�b�~�!%�Txo&���DQ戨ԉyI)?זchE<a <U�?�9UY��]U(�MYU�2�9�>�/�-�Mr�OY�	����6N�Ka{bL�/����V�;�,EǱ
�TAr�{�jz'�oz�o��jo逼+�,�����6�>�:���Ƿ�ښ̴����S�J���/��\.'btP�=��1������S��!~�'�9I)� `����HcD��-��2JηS%-�!�!��$ْa��Q]��b{}���n������f��=�}���Q]��{��',t(�@Ǣ��J�w�VH�3��|���DpØaG�^0�
��a�����c�P�����*4��8�	��EɫY��U%=q1Q��V�������E���j���JyNL"��ם��,���z�Ϝ��}�����;��-Ƹ�V�-��Ϡ�ʸ-��۹�,V.ze���H�v>�*��j��ڂ��������Ξo}��p�Ty��d-�v�Ң˞p���l��b�.�{��/�tJFC���諕]�; S0���,#��:����k0�������4xh_*�YxP���u:X�'�1�p.ፇ�Q�Q�k��TI
��?�3u���m,�Wa±}�q\���R�y�����iG&�Â��b�Su���B�,�%&��������G�;�G/��g�:-��?>K�h&��Ǘ��Y�  R~E6�uj%�V*%q\%반����X��j>�.�ގ�眽N����Q��� ������|�ueL�@��o�϶��$�r`G��6��d��#�4C��1BQ�p�y	��y^�E�&	�Z2%N���7Ֆ�I�EG�[#������+�Z@��r������GJ�Ј�.D��q�E[�P!�ׁ\At��i!���Ue悤��?�(u!�nnC�c��gÔ�����W�������h���̿H�8}�����y)`$m��p�Ἲ��>�a�PQp�늩��;�~W�_��E�߅DP�Rbӈ��:67�R��ܠ~Р�U��^��4��B���k���=�j�G\��%R������u\�C`Յ�Pdƪ�����~Q�M*�b�������u���ʍ"$:�"��V���9��}�J����-;#�I�T��Q���
�k}��D��s��s��y7rʽl}�F����d����x3��M������R�Ū��B(𢋖�3�4s.d�i�QYW��Z���>���]t��H�Z/�eJ��'� .�H�I�^#��L�ݿ��V���D�#�T=�׆��$l���;�I�r^C��%\4R��4ȱr+�R�$ʁ��'٫��sc?��y3��N�_HXZ�Zf��h��76Y��� ښȉN����N{9�c4�cbR���aNZ�i)��^��4�Kf�d)ݐ�'eZs��@���8��it��̓�5��k��=D
��e�۬m��侵����`{i,fؐf7�6>}Dj���BUa�\Pʬ�[f������T����j��d֞QM�u�{��$ƨ��(�,"7Xs������u{��9�xڽҖ.4��rt)�Kf�JX�	tN�k�c�\:@����:���`���*�-����u���� �P;�޵TsJ.SP�7�����6�=g!Y*�蜰��'��8{����9? ��T��8���$i�<tI��sx�_2�lj^�X�����*^��d��a d�'v?�f��<ʟ�VH��I�l�g�8���W��C��8ki��aS	*�QR�� S��`��*��� �I�uL��SG��U�p�DY��a�W�QKѠ�� Wk�.�?�=9f���1��݄S(R/��d�@����%`g��Ջ��8Z
j�ַ�����W�ǱW���)�6����9�4�		h��g]�~�e�פ)�KL�@��[��%�G���^*��
��+X����`~����л�`M^���Adw�(����kI���^㉀����V}X(��X�Y�\U�$��㪔<;��u{-+̏�(V�Ρ�1���B;?�.�blV�A����Ѻ'"�Y2���h�Q%P�]ݪ��a�K5��^O�c�K0��eI�L���ڍ+q�_xk8��g�������&v�=�\���9�|6W��C)����I4�[��̗h��3r캋���y%������:LP�yL2RFWxPel^�fG$�(�]#�F&�9X�BD��Le�t�&)F����w�ʽ�ye��9��=a�@L��a�r�d��S�Ǻ��k��������9��f��ʿ[�خ�!�3�e��_��W��
��O[3=B��wa�u���.��~WEW���16F�m�� �.yĻ��]�4��u��1w"h��e�=��Ժ��EiZ/#go�G�ұ�e.�	�lL�r�`c�ĝ��UԸ���i�ἸA���)a�/��- �dJ	�:荖Ҡ�e��-G��G���7��TI�D,�	"3�^q(OeNK��W�O�� ![��;��Ɔ:�};d�
g�?�6�K�j�$�V�%�)��m<��!n���DϨn�kp�t�|E�ʲZv�63ٛ����#`�՝*/���ܝ	�!z�>ard�79b�+�ytf%�c`�S۝�>�0�����H�)g�/D��]�&	���&u^t��Yf��t�cV�]so(I,��9	�S�̌�	��p� ����T�̱u�v�
)���ۆ.�*�4����y��<]�D�Z6��h�n���%k_�����HñQ'Bl$+ϙ��_�zi��gs�瞛5�䰵ym�t܎s����q�@��Ba
;�RcS׬��BT$O���f�9�J���3������RA^H�I�/9ϐ?�3��)
	<Z�m<��%����^��QFv#���㗐���N\�3�JV�[{-�f��RPE&�i��Oh;���h�Bٙb�~��5atV����4�U�`Uh>A��Ɉ�������2@�@��9[?�#�u�,��nU[�� ���C(�f�0��Q�� ���@�n].�걧�|��]mm����'�qnx�\�)Nm�Z�6�ښ-���e-^)9n����,'��IO�����_VϤG~�~"%���S�D���_�g�=v�"��g0�����s'���i�f�3��!��JR�#i2+�9Ky�>�X2���P������L�=�ni`������N�R�e�PP�4��Y�,H==�@#��
�F��W��e�"���K�7�����V=��/*7��$����- ��	X�{��0����M��kBr��X��zH�8*�X �yEz�� d���O
��$ q�"C�ĉ�aJɌu"�,�+eO�x�ӭ�}b��W��D���s�d;,��f]4�=GD�-α����1?dԩa� �7����Wc�;mF��0�[�9\��˷�nΔ�����2��D6ٹnt�{���WȚ�q��D_��e�o�Xb��E�w�j�/;�bͺ����I%�W)|�ʹ�IB�%k�
$'�����?�٠h�Zc:X��/��d�W�<��a���<�	�9�G
��}���x����W�VQ��E�-w�"@��A���}��!8R��x��YJʝ��sm���G?�-6�iu�,����r�^1��p��I�*S����VtW3^�UF��'���WH��Q�B��|����W�}g����9�x���6&����q�u�7� ���,��q�y�W!��++�� �.P}�;؜8��\�4��K'E`��k{����(0!�:Oq���=��D��R&�Q�V�$}�S�k�p<�~���o�q�K6���I���Y�pʰ��������;��HV�.�\��(YA$������cz�K�1�eL���)��c���8�Ł�I��J��_���,(�N������f��,��g�����b�eU-9)bSO� ) ?v��������O/��2AS(���Pk�]����.��w�(����f"r�`60�Pe?N
�p�0���6����\�c��&i��B5��-M�,�e0��4�O\\m9+?}�w�
�ՂX��t���J���$�~O�O���m�:��8�B��y�Zh�
���0l����o@o��D�I��|��p�z�9�)+��|�@�c��-*���~Q�V��C׬���P�b��a*]o�@j'ږ��&c8���Yf?���!�h6�;Dȕ�j� ��=]<���������2�r�p��E�j����;����6T��qwZ�j遣�Bj!�j��f�F��Z�yt���ׁ�� �����^ҝ�i;h�T����OΡ � KXҝ:T��E��	1�893$�܌E��Ps>eMK�:03���]��<�jC�<��g�H6�C�&��W�^M.�ۜ�sG^w���`�}.&�;���+F������8�Lr�QZ�w��6+�XSw���ω���&=OR 6���k[F�ј�������+z�I�ɳ:'�5_�,��h�_�B�Yf�O��I2�+�������!�����n�s�G��]t�,�;�K�n���[���KhAhk)�Q<��C��\J1I�Na��b�ҭ����	�VWy�6sх#���a9��B�#u� ����\op�YN��\���P�ֽ!Nm��#��ɴ]��uZc'�S�-�Q8�X�|��[,������\>I�C@yY�д4*]s>���x&l?� �x("�s/�Aj���c�r#�4;^xo�9ʙ��d�Z� �Z�1ד��ؗﷄ�=�D��(�6��|>6E�zt�v�5��٥=bćfV��0�
 �Zhe3����~�?v�oZzu��꫸��a�u���|,�� ~ƻB�F	��gL��_���ݱ����e6^��AQ�;��?ƀ
�:>�'��jWZWњ.PD� _!;���0C���,���OjܘU��hi&�4�b��p�q�W����Z� ܋>��5�o�c���xZ/�)KO��+�u$[Eu%���x/�Au�o�B����uն(�mN�@`s�<%57e �����ha5��`A����f�W#���h*�*_�3�j�E��#%��0�p/x��W.���K��y�(�]c�,�a��\��mSK����gTrvv�4���7%���	R�K���q���L��� %7�K$���D!$csH��H����V�W{2i�]�˥��J&7�.��%������YЛi��j�<@��=ł5�3EA� /r��ɚ	�fzc��d�4H?`Ge:py��~��)e$�D�ݻK�R��΁���@Q:� �e�r��(���=���I �`�e
�V�$����w����*)�yP�'}F��y����L6ẞ'���܇Os��,�a,+F�y�:�Ҧ����_2������E
ʚ��q�I����}97P�|��x�ӗ��7\l\�AB+�vo!�
 i���[�v7M⸋;�{Ѵ�Z�.y�皊&V�a=���)�p�C�q�O����R���P�?�@��p$��Eu����P�nxK ����=�P��w����ݑ������c��X�nm-s*� �}g��Qߛ����-�׿!z`^T�����&���5]��� pr=�}�����$G���픅�ܔ�!��@f�sU���p�ZK�qr�Ya���Ξ��ㄬ")�\X߲Bh�~aJ��yud����S���I����<ƑYn��År��������-�RQ$���:���ƓgА[�`Q���R<�6rX��9َ��2���-;6(O;&K��ܺVVW�ں����A�X���]G�t<�`�6�I	 t��� AEs�������h��S��uњn�K�U���ct�-!���(� :�L�A �Z@+��³�m��Ĭ��#Z\�_K4C�/	Ø.X��V}��zg,�_�"|ڠ3,a���"�?�6;%t�K�)�73�I��飊p��핱���|Ǧ����/B-��5�6�� �*	X�Q�!��"�B~v�jG�u0W����S�h"��ҿ0mLo^�7�3Ee���x_~����y��Wu TJ�ί�Oo��e��pG��Jc>B?ar`�@�ō���[AԕBV}��Hc:D�
�qLu��J��sS=N~u.�V����/�<S��v�V�Zo��������R�ge5�_��G��諺]�NgR��:�U�L���6]��ǯ[D*4O�	�؅�Ii��"n���6���v���ZY���X0�
�(�Ly2����y�q�N��D�sT�����k�϶?��%,�����ʤ��i�����Cy2
���R�gIѝ���X��㼚\6lܡ$P��!L���pv�)8Nʀp	�ZZbW<�ЎN�15�ZD"��N�`�W��J&�g���J?_�:�ȨB[����X�U �B��ο�+�`v�{�f�ͅg߃�����X�IS�StW�h����H��W()�7s�������پ��E�P��-��&�(�����iG�<���H���U�zfL(?$�z�.��Y�����zvfEe�d�{~X��q�j�eC�
�#����Z�1����bP�����BPA�X��"���%(�}%�u���$� �=��Ŭ-#�E1Y���� +�-[��fswD`):,ad �s���j��H��Y����Π�:/�]��v���t��wf��,�P�'ET�=�L������ٚ�P>�`/��`���w�!dG*�{
�"�Ӷ�C��j�ƿ+1~j:Bs�6�IL���c�z����g�E�����/�f��A��^�բީ_�	�:ng��,��x�����-V��˞.���9�Xu�>D/Sh*�!�!����m�L�D�g��f|Y1P��Oz{⼸#*/����ev�]�=s¨����T����|�I�����5x�����H4d��p�S	=�#�g�&�$��0����\�3d4g*���%��V�Jz條��m.ٲ��>�����kd�1jI��2�K�����˥��!��`�{�� �hd�%"���I�Zpڬ:�
�8�L��3S�e��a����q��X�D%őN� %�\���5v�mc����u@���7k}���a�u� �fI9^�o��=��,�fV�%��&p���T?��pj��
�O��6�o#4�x��J�66v�L�b�&�(Xl�8�Y���j
����G�I��Z��Y���SK1w�z�N�>���`2ю����f�Vj��$$����������!�BQ���z(w
��\��`��,�PCPq�jq��ɍ��n9\�B�h:GZ�|�ћ����2�t@�Q�\&�DC�`�wcrL��g��.�?`u��D�O,�Ī�c�Z��;1p$�u��RvM��r�d� �Ҳ	��u	��+�Ɖ���1ìS��Q�'C(����N�}�MgF��0��m�)5���d��ˮޚ����A���X�ű���Y
,f����Hk���g��-s�E9w�`�7.RP�����kGC�I��V�8&�S��<c�M)�9�kZz
����/xmX�M}�������Wtk�2�8k��0�{�׬�B]ͪ�~:�5m�f77cy��y���8ތ18�q���p�2��~8)���au�=����L��Q꺄52���=�٪0KQwH�����I�ƿA������Ga�=�|s׈�Vz����_�ԣ���8ß�D�;�:��U����rr�9��7ww�e��Y�w��*�\W�{8�[a�H���/#�=J�,�OCC�?��d��*+���R�e�aw��7b�+���|u��斉zo���I:�~E�q���Qi�)�g7�_�ahq$֨ԠlR���������J_���L��)V؏��f�
t|qd��
7W���w	_W�~�4q��kX�H7I~���Ze��y+"��x����U�4c������#�h�c=�
�U.�K�9�:P�~伴u!�Ir!k�6M�A�� NB����