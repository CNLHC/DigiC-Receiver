��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M������O���R�$�lIlqֿT����N�B���Wg��i�ٝ#ei-�#�D�ዣ�I��n�;'���6!�M�4`N���ꚢ�ы>yx�w���r�'��	BsG��/#6���Qpt�!�yݠ���:�2[Hb�(��_@i,���[_�xW�M�����������XZ=��~�d���IV�S>��d,BtL7����c��q� �>�؀���x�%y�;É�%�s)�@b�������At�}��YX�iDk�"���vX�<ts�ޖ0��c��+��F,ٖN��C5��Ƙ�V$,��̯�Y��߼�-<
��7`D��ds�bNP��oC���(��a��b2�,����lҿ?+�
<�ck��)�c0�as��å�����1�8��?Z�1{"�c�?\& ��Q�>�;���: �1'��;/zz�k ����Hz^f�^1�8��8��y"���>�uȔ�d5����i��'�4�zg.��Q���g���.�7�<���9w�������N
�B�μ"F9�`P�����z�*4�"�-�=�y��Z��M�9a���AH_
��g��P-��=�9��
�ex��;:u�8��17�~a�7�����[�:�r0<%�^�Q`[�ΐ%��	H�Y�s���~���ր�_����3���'��
/t[SQY�!9v����>X���,܈D ��f��p�<%սq|��y���������Ŝ��F�c�v���\�3{��S	S������ fo�Oc��^<*�W;�I�h&H���&[7�Ǜ���L��3 ��d�z�R����,����k�%Prug���Ҝ>(>�H"c~��%a���E�<�Z�K��x�TA����y�so�_%��������Y�Z�o:��k�4O�C�on���#m��g6FS#wT)0��[��0��=O\�Naŷ�j�p���s���;2A{U��+�:���A)�%�]�1�2�~�U��W��/���.�Õ��+� ��vEn�6x:S)=�<�'kKq9*A\�m#��}���_k���ͤ�2��S=Y3̪k�b�ЍN��)Uװ��*-y����ĥ�̖�8��<zЌ��S�=��׿娩N������Ț�ذ���ʴ\4Z�-�n��E�o;˟KŖ��We�RQ[-���t��n�xŲ�Y�5� �/���zU�7�1�̘AQ:\�^n]|�?W��T� ˪� x\����z�A x��j�<�HN����$Æ@�
��̏��cyXXD	�� ��l�UE�\�2���;s�-8���w>�o��X�������� �!A�Q��L܌b�Cj)�1�R��h�mG,b΢��&�����\*ӽ�{�v��kN�L����#���)�����z8�A�K|������,���)���k1PJM����pV�:Rt&Ơ��Mu/�ա%���g4�h�qgP�B�;�!.�`�orX.�j���n�E�������կ�v�{ ����ӱl���H�&� �76��K�5���M�nu_t�'7�+c�;�b�,&�&��?�	u�I��T.�9�$�EA��~T��l�h�X�E�l�_�h�,XA�?�:�177�z�.�3ڦY��V;
h���'���A�z#���9���/�7DÅ%1�m43LR���5�bs�8i6t����lCf)����$R��}��|-�.�
�gcN�<���0�����Fڂ5M��Ϫ����	fdA�������9Qgϱ�i��q�Ej)EC�P1�Q��)��bV84POܥ�D^9�N�W>@#$�]B��	C�yd!�&�Q4������b��}v���Eh1�,���"������_8��y'HǶ�+{��~���繃�v/J��=�Tw�,v�P�9�5U\&��wI0�O�:��I+�.]'���P�4��~pJ@��fa�}�m{��KS{�ic��ʲ~hc�R�>݊��!�)��� vg�O�}S�������(rLCk�'6�S������:ez��U�{�>�	�� �;���L�OI��%��n�
�ߴ���aO���U�y(C?z����%�F����)�zu@Z��1�*����}.��t蛄������ղ\�o�Q$ (d���R�T��
䣛�d�Y>`�@��e�� l�}�� �P�[B'u{���~��Rzx		��y�"���|�t�@��z+���/mb�O?H����d�ȓ�Յ���C`-�P��)�'��N�~�-��R����f���QHiʔI���KC�ii}�8lx7��W������5Â�]�H"��'h�1�C������*R��?��Ƥ��	K�0����_�#���X����K� ވ�S[�tq���¼& K�{E%�P�PFZP:��L|?i��"�q�}xm港��=�l�V�7cq�HQZo���.r����;�iI�v�%J�S�ʊLtZ(F�8�l��ا~/ �UO���Hz�	y�s��T�Z^�[�T�sh�����t	�߰�,\[��%��K����17��m���"���~n�$���! �^N��N������^����w@���@�h���&�j���,e�;6B��63�MC}ȋ
�pE�@6Vz�^_��=�ehG+�<��_n9�6 VC�1|�hBN��I_�Z��׀#Z�@'��k9�h��n�bJ�މ?� [Y[�u'��^��U�0O4Yxi ��d2q�t��OvL�u����7��Ĥ6�/2zq��ƜK��
��Q߻tx.�M"�G��z2��Q���v�<���'� ����⟨�d��9[��x���z������B�|���4!̀��o��h�}�\��0�\
�9B�<�[V����4M�B�c���3�E�߰�%�[��9|1tX���ē�!x^��0�������׏�n4��{���j�x7��WG
�m�:��sr��3�k���6l���ׂ�{� (��c��g9	^r�h�܊�|*��� -���vz�Z�O��j��.�x��i���a5���{?�.�ٶL���SU� A�ӳ���'��Av����;p��5��Q�6� %����5o
�p%�T6	���Ksw�3�^�]�we+W�ĲN�Ûy^�:��y~$�g�9z�9�^�c��HR�8�[��l�j�O[��]��[��Q�������s��S&��-�.�����>.�1#5S���9�~I!��J^sU6qP���ʋ��;�y�+\�%Vb�O^{��,U��|�|Z�hN�#�\ף�6�-�PO���V�ˤ�g82��+�C�y�y+��F!����9B����zaf/c�����ž\։1�:g����Uk���\:���P�,�*�9�a�T����-@T�����#/$�r���(��E�0����H��o)��e�u�C`YD�˟k�`. ��<|ˏ��Y=��:��n➅yi��5?L#���,ɴ-�A�3�Y�8mm?�Ih�5b�(�f�q�̿}O=��QwR�G̎�����!G��ث>u3+����v$��<����U��.���|w��ͷ+)ǽ*��Q�>wWI�)��a��	�)Z�����9�$���L����Oy����EZZw�!_�NI=7�`��ɪN�b���9B��gP��idV�>�f�L��/��?9�?^z�n?��n�D��"��/?B�(u�/��mN�K��Xd����m�|�ޱ-����-5� Mg`��ˆ���~�r�!�K���z/FRc%_������=
^���q"�줞�h	�Ñ�q��O�c��kc[)lK&z�mp����������Ջ�����Ӏ����R��G\<:<(�T4;k�)4����! `Bu�C!s`k,u�~^p���i. �@ާ;�� ��s���B�ڱ���� 3�-c���q,a�ȡn+\y3��p��ʗl�*jX��8�L���^;.�[aT�y,�}4�u-C'I�]�������|�W�{��c^��:�_(p������PZu|Q�q� {����ĭtL�D�h�3 تg���:v�r�Ѡa�}8������Ἧ�u$+fd�&3|��7�ܛtd<�1�C�l��%5����80��W��NdT:L;R��Py4��B��,@�a�� -�9�=�qI鵇}��m�6,^A�#w�x84F
� ��W����,Љc�;�m�J&�+r@;�G�f��гY�ybS�tۗ�kj�}������A&�E�4��K@�����dTwJ�j�"�4�\k���]
�&�P�&�˲ͿC�����GW]1}�8¶��If�L4��igkL��q`wբd���*<Sh�vLeV#S�i
v�ӊ�/�̀�y��&�O�{9;�\ɶ*�8�Y��7n}�K,zT��Vڇ�*9/����XQ�Lq¢�Z�)�}@�%���6ch��>�稁:����
7�s�h��Jz��׳)cɋ%��n��Rݵ$��׃(�9���6��c<��3���;����Q=&�נ���䝴#�/�56s�wD�ϓ�?z� dD$�x�l�^1"ci��љ9`���vt�?G�&�E�!e:&f��8+s�=aԐ�lsޝ��pV��>�M�*
��Zu�L�yxh3��/���-��k�K��Ǔ;mO<�c	�(J��#���GV5�
.ŬZ�d"<�9^�c\�d��q:@�z�&.�f�f�<�*���{<eЋ�J�5@|l9:}�hZ�~��9�I�WY~�W����[�殘,I��U�B?�'H����L!l|\9�cލ��T�Q��5��d�`r�����~[b��{>K�v"J|�x &}�Blge���r� ���bĕ��q�&��٤�R-e�.�\�|=�6�.�h���h��{�Ic��p�)���L�L��P�(��x����B=���3�żs�:!>�v0���z��S�aL�Ut��v�etH�����T�*AI�RE�{ԃ�,�!o� &jU����ꛘ�\�Iyą�d��Ҹ;2�3Y�*dE� ���:7w�HL΢!���I�Lù��*2�q���|!s�H����ѓ2<�D�)�>�HϢ�j�š�n��'�FL�����Ijx��囬������e�����4�!:��$�m�qN��u/e�Yx�b���62��^i������f��m��G%�����~���gc��G8'��ܮ��y��N)pMe�?�eQ;��?���_�?鬽UD��=��iۀ�{��S�����E������A��,�S�p�q�"�V���p%�Tl�&�$�6��D�hs�1[�ovy{��,O�	Fϻ[/.�w�4���a��g3����n<�AG��>M���ٰ��ChX"p7�҈�p<��|�5�ָ�X(2֕��H��tS]��$����M�.�3͡h��6xz
��V[N��.G,%���2.(/���䞦��H"O���P1ZV��KJJ��|�O���X�<����j����1���B�iO�^臑s�|~�9D#���{ǃ��:�v�;�na�J> uo���{�C�� ��SAx�H6�9b�` �v�d����g��hX.D@6l��?,��Wا�R�5Z[�ت���X�Y�`�j�-�n}� l��L,`����3�r)�?�{<�Ƅ��J삸�L���;�Y�ٍN��<����.��#���F"թV
]<:��J4rAӕ�ΰ��qS�>k��Z]�NT?��n����.��,ѩ.$ �1d���>�DWT�5
`���6�K�2���*����������pi��6�G}Qi$����@|[���Mf�x��
���=X�:Lo+���`�s1�Y�%�뾯�u�������)�zъ}��~�/���8|:�I��и�m�s�,�}F+�q�#G����U���s�E�/�}��'�L4�a�{5���-)W\Ib��E��a��=?b�R.��>�p��N���<n2�[n�Eߊa�=^��E"�v�R�|L��~kǍ ���L{�w������.W;L���d?~%��e���؋�C��Og/e���E�>��楗�?K����쨴W�	gl��q�=.h��D�QnX9�+��mVT��9z�%���n0E�Jw����t�G��{ ���"�%�J?7yE�Y�Z�=��-�c��,I��tRf��5H�A鵻4|hj�:��m��r^/YM���̮���TAw3�L���#���q9�8V4��<���:�,��@��9c�ņ�
�+����\&�F.lq/g���7Ŕ��릜�z�{��R� t�$T�ny���|�ѳ^+�
!؊�B]|�fSj*�Z�&qnY	4y����R�Ƭ6�=^q�'��A�KȌ��/5�=TH+�}�}%Δ��9�g�^-^�K5!�Ĕ핌��n�Ѩ}lohʽ��r�s��Ӫ�O6'���M�$^�.O��U~�y����<�9������Kx���ꎇso.O�Ӿz�Cs���)h�@�`e�Z�{{�EV/ƃ�o!�Oo���X�G@��$*���/9�<�j7��_N��ٕ@�_"u�_hp>U&S6������!�y�X'����A�zb��{�?B�e8UCf��xX�)|G˾?��5c�������5dx��#1�iN������}�X��q��Ȓ��KQ2-��~x��Hbvla)�:c"�i�vS�|O��t�G�{����x���?���H�٤s��:KMLS+Np��>�D�/j����2{t,