��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���5p������H�4�z*Gh��C)��i5=��_�{���Q��7�,S>��>�Uë��
;���1�-^�u
��-њ`��|��f�"
1�0���X�Gb=px�0��0ד�e������u�P�j��\{3��M*0���Pm���?ᐏ���O�9ʰn�*��� �ڠP	��`�;P�l�&��IW18�y)��h���9����8��U��$�l��D�V�ND���
L&��i�S3����ܴ3
!�,���q�����S[H�bž{�+�`/���?@>>�F�J��[ �w��쟎�N��G�i�^�^��	F�}��^�Q���!:��D���o7ߎ�j�V�ᝂ�u4Әknq�����'D���K�"���e%k�7G�&��[(�0N���E��"U391��6k�d}��b�p�}�6�e�l�18���hy�?9�o���l��F�G��.��ه� I1_G��M�o'�i����m�M��;*����@�_��؆���v���\����KO�4�#p��ih2+8);A�t?}-��
�����~ﯱ=Qo��/�uOouY4�-7�4#�����Ȣ��c��z	U���p^�q��#��79ɦ������ToO\��.*�Ѕ3��ҫg�Kp��V'S1�_����zZ_�o��;�3MG�S_w��yt18�}�9+1jX炖�<�*.Jt�Ɏ}��ޏlQ�$�T�Y�VP�s��>nȄ%�L�Ba����Pɓ�5�*��n��˱��e�I�W�Q�� f��N3E�V��ɫ��R�����%�4�'���Ye�
�!�0vE[63�H#a8�U���9�N�<���s�����I9:5�<"��)S��H!��--!�o��FF�|=[!7�PZ��T�A%^>��e}�))��M���*B���s����4���m\ڍ_e������(hU͡�
�צ5��xG�.>�Q��I��c =۽Sy���3��Z[u����Pn|q���fېpFX�?iy��F0��ư��,=�S�L7тrO���\S,�F����Wh����P�t�)
�ֵu�j�(��P:����\$e�E6�ʹT�>�g���XhY�N9���2�p��̴E�z�7��>V��<,>����T�#��������m�S'��i��y�v���S��$$�J{�2��Hh���lЃ���}	�ۇ�P���`�!{M f�5=^�#�4eé�u	Fτ����j�#���a�K�i翷L�>m.ҜU	�����U�@@�V��"M�~�a�(h��x?�GX1��,��^�٪�d�پeъ<����	�F6�<������s��z�F��+;���[,������㥍�A��)�-tYU{uRN�+�(?�1�q9�p���6k�s2[�v�F�J7O��D���<v4�}O���C�>܃��� ,ѩ1��H�2�~��j1���g�L��k��xØ��^B��D�z�~�T$�ڬd1�b��*�\�5t��<��[L�������J6���j��-i�e;	�㋆"���ELj}�U�Ӵ�j��}��l�!"֎Y�d�_F�x,��K��nP)0�O�$ �Z�m�&��k{�<����Q�'��d' ��:[p ��Jxv�ήw���o�~28�f���v~	X]Կ�S�*�29��>|r44t����A@P_J��}��#�3�_M����w�6IӢ�9w?�t���F����!��h�Y��{
x��aN	�����کJ��_Nm�}��j���X��#I��.BT��I�n�|&�u����kZ��>D�4$��ν���4�S�l�LR�k)NA�r=�i	]!�B�R\[��3i{�-a|���Ǩ�t[	ch;���I��ȄK��O�3D ��j�y���� �܋��%�Ŷ�
��ϛ���7(f�0���`�����抰M1�HR�,w@q�t5��c�p >���J{�ݾ�~�]��R�T�SS�KU >����g ��9��j����y5��T3��}R��2(�+�w��%���Q��l[��c��E�F&�Ĉ6��ب0���R,�N�p�>O�%�����SOgΠT��Д��B��̊XBk����o����O������D&Ic�N�[��' ��O���w���=n BK��.��M%�<��c#�QEj�:1(9Ad�ޓQ�j3ר{�0��ȹm<zp�U$���.zD������v
g>���ꇇ�_�F�ϱ4���M&m%.N�Q��4������r(�)��P)NS?Zڭ��1���������f���ST����C�"����3A���S�C�.�b�g��\�RI��%ǁ|ՙ�%I���TRNmtOqw;AiiuF�ֱ@
]��~[ ��R�]��*�����z/ݙ�d�6��7�<�Yn�v��f-�ѧ�g0�+���$	�f!}A�n��qyQ��dfn��:f~��_R9���L�ס��V��|{�%���C�^d�ӻ&�����|�hA�l����{�$q��ȣ?7$�����ԆS�,���
�80��������!�'���,ə��n��<V)j�B��M! ��Y?R�U�@+�Ɔ�YT�^�ӑH���Ͼ�<���d���
o���9�W���I����!'VC�o��lS���ʴJO��y�ǘ��ô-��V��M8| ��t?�m�W׺����H��Ҋ���'(v��w6/?�חD$��<���S^Q a�V���^3J
�>ƿ�l�4Gcyױތu�����	�q��IU��H�P�ڒ���R&�`�E��В���=jp�uV|!�u��!�&�� �2�����yT�P�ln��ӫ�^:&����ZP�[RX�"�K�!��)Ӥ��E��^�Qc=Œ�Z��lW�1W<_g���q�~,ߝ�bỨ�]��믵��DM��>�����h�L$�:��%�劸����	9�5����WP����vy[�.)����T#�\cr(T%�al��4��Qz����������m=*U�,�/��	�L� �KG���f�����o9���C	e�J��Ʈ�w�|�s�;"�U���"7�5����< �G�|����`���s���aȕ/�6��u�9�̳�6�ʶ�^�FS�K��A=�.O;�����s������V/&)���L��� �RԔ_�KO�x�۬A���,#l�Ϟ��1�x�Mn7DK��P���X�� <Z��ٖ �3)�}n3H�-%�/yA��W{~��V`�q�]m�29�U��S�Qk0z�Ë�_�4ns
��z��R{�V<�ɝTKD��$nRS��i�3��
P�� x�)�z(]y����/c�X���G�5�v���WC�%wl'�7
-n)s�zi�Z)A����cL��3��1��'x9�ѳ�0�fU>Npz�r1�k�z��䮥ʖ�D���Mj�}`�`��K����G��)�*��	]��aoP�ܽ�e�=p�rI�g����2��!�;�\���ko��wK˒~���<T���w��d�	ߺ����		N�ל����Y &ߨfE�^g�q�(#}n�S�B0��_�C[����������<&(�ӱ�����v��_c�w,�=��[��o)��<�V�8ZIg�B�*F�90�7ksS���t��i���J@.qE�I�o_^�	��p�.;��ɍ.��y�9�(M�u��_�5��|��z�^((D����.Ю�Q�� f�0	`��tu�@���sC7�&s���h �K����H�4��&���L&x�O7^��TVI��۶�F:(Έ��>�7��-J�����*��o��l�f��}}î[w{�ns��2�gM/���E���\$�'e=c�+���k�t�����lT£A�a�WQ�PX�E�j5�O��-Oa��+���Bꮔ�:7��$/�~��hfM? 	�Ƅ�� ����_�`�GݤEY�D�@��n��%4_^DǸ*+S0߻����T�!;���P
"�͎�$C0�"s�����%��I˺�Щ� ���9���5�rk�����k�a�X,9�Z(o!��=
�-[���.�ڂx�Q�����CB"VA��e���}T֕�����%8�և�ʐY����l���)������{�M�%S�>���j�'#���:�j7�u{��*�Mĸ�g�@��	C۝� �z٬��]')d	e$�B��-J�1��ʛ��ؒ�ǩ%[�qI�ݩḇ��Hje7E���e���g��x�L0 d:��� ���E�:B�l3��RH��{�-���|��$2�C��AC.l��F.$ ��T�Y�y}��m&1m\�����-�?�L��WQ�(K�D���_d�%�����!a�l��CF��A��� �����]l���BQ���@v����;��8���
�X�j�ܰ;�N���Uiؖ�v"V��'��Y��&�biʟ,ǥ޴��ɿ�ߜ�	"2D�Qw��� ���z�7��D��85����nj�8G	��t]1�T����[��������ī��9Uix����%^���G�#7�Vm�3��`�A�߻�m���+>Pg8B=