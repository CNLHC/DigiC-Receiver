��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��.ܗ��z��Ytԅ����Z�ЊF_�}�m�J�����K=�{�d]�����j>B.� �1��\�:��N呮�Mg�d�>ϡ�_ؒو�gQ� +Y�o1�E�4����w�RJ"�E�:yKi��fJ��@�������8�#�t���`�W�u�t(S����=�-%#W�^����j�N"�P'� ���Bc�>k+��M��5�e����)#t�K�j&�6T�FL��],���|����|R��Ā'��?6���Tx�.�~�$�;��2�8E:�tU�z�0"���%O�t+"��,AP~?-�4`^ι��]Z��Z��]c���죓�5x[��ț\�P����(�Q/�×����H�t^)C�C#+��!េLp�+J�x��Ur�� :�=�5
Ī��޲�����7F���7���~����k(����J!��֑Pbm�$rQ��� K�0!�/@��"��p��p���{헖��_C�-��/��|��8 L��^�ȕø����bfF�t[&����2c�e�*;g+������}j��t�(;�],޼9_�GIE�K�N�`	�WO\62FKC`��Hƶ����K\��|�|�w�]�9��7���[A�G���mo\���.�$�q��s�1٩�G0V]�_��9���f�7�����2�(�#fQ^����*C�C��J��c�Iǃ#2x�٠' ��I���:��ֵR��ME�hlyg�!�r���"� !�(�]�Ν��VW��ZƼl$:��X�)��O��ˋ�\>$I�����
<!��ś����3O��y�5���g��|�G9��fz�P��	9�x��vW�A �--W:>k�g�2�N��.Z.���<���a�/�P]��߽�w:n=��	?t���>8v=L�cbM	`_��M&a��4��X��ֹp��N{�xƖNM�s:\t��ҤM�E�J�^@��@� '�r�Fm
��u���&ڠ⊾q�*yz����tv�;���3f#�T��;
'�?�_<R�9��ރ�כ]]���+�ђ�#�a��K��)[��,l�V�=���������/)DST�A�>Y���m���8��=X#���_F���=Z��1��p\�����D
d�Ǒ=�Q)���� Ȥ�~A��mX�Ϟ��5�)�Tfi��+&�����pLK��n2���_���\Lu�A@�|���E!��~��`?7��R�,0yJ��[�7@�;�&�R7Y�z����#�J���N'	A5���<\)>���HF<���gU�@�ߑ��B1O@x�v`i�u�*��^4��AY�]�����0������Q��q�}��
o �i�S�|&m��1\�<�X:��r�ꌯ�*>����8w4��4�������`��b&�t>�.��![�����`PH��O2�i+`Ӡ���Y{���D<�KZi��덼�S��}�w�p�n��,4~�[qX�,oҰ�����vj�OVWvʙڐ�\��t� ��\T��B�d��L-	Z�M[�����?K��6�h3��[9���GZ�9����M����~�G\��S�F"�*�(\_�k���<n_<P9��
��Ë�?m���c���"E���|��0U��E��p5y(�t� B����-0��=ga,�1?^r�ff�sL����9���On]�ҙ��]��GÏ���`-r�/T���I�U�V7�7b���J�7`��j��D�ю���}�k�X�2��cj|�R�_�����Eq��hň��׫��1��B��Q*H��=��Uk����Ⱥ��XXZՁ�8ўޢBi�V���Ac�F�=(h�7���<������4K��j����|���^$��u���Gg�L�!74l�0q�]=�p�@Y�-ا��DGD��J����Z���@ւ���ϐ%ԁi��w��q�M�uК ��7��z��� *�V@�G)�Ql�~)D�?T[[ua�����7�R��8�F!X�Z�8�	J�x~�ۭN�.�t��x��#�&�Ghj%�R�9dw!�b'�x�2�q���9�K�����ݿf������v�i8��+��R�J"MN����Y�]5��h$��=oLʃ��r�ق�K[5�&�G��O�Ӄt~;����y��ʃ�2_��I{�+¨�F�J
����X�&�lO�]���컵85ʻmУ;xYǔw����K�M(�SY1�QCEהLH�icc�:t���9�'�8?5���.�K�'x7��m���;]<�0�N $�LG����	���0 ���2���C.�r�<Z��c7a�� �&a�M	;O0fX�3,C�q�%����WR@��9�o�G�������u���hT̕�G[��G	��y}Wua�|��l,��p��e�w��#�n^p�ֿ�0��t��5�d�jҹ��[Gcq�<�s�M m�z*�%� �`�4�>����Ak/�~e�x�H<"���u3J_0���!q�\��-� ��gE��Aw�t��Am��踽4��d�P�A�h�y�Q��{ρ&������zZ�.��zW�w�LNGA���Oq@w������+���0g�P�������d���P�h��G�0��W�����d!�PmY8GI$��ؤ�v	A����� �h9�J����dBg3��S,�����`r)�D�����Ԯ�KO!F�: 6Id�����Ha�x�V���*����;��m(�0U�Ř)��<8t��u����8���!
�f�rk?TY�>0#翈�7��$J���9��mi�\� ��S~�tL�{.����P�~�1���Ev����h���ň����!�j�n�/&=Cx,�\��'���V%����%׀y�7o�O�$���5�%/%��$�~i(\���kBj`Me L��Z�*���6M¤��)6&��r~N���%�����{ˑE�9���Q�\�s���a2G��n5�+ �A��Y�"����t�ݯ\C�O���WF2�"I��jk'򰲊�m� /Vi/K��x.�H�蹱C��cA㻷�i�kJ��9�Qgel�k�*�0���	���R�ڃ���c-5;���m~��F�l\�v��3Z���Y/�rqD�����rcZ�kuN�6���:M�fs�����v��E���{{�ec숀�}��e4m��qh��W��3d}�
���m*���뀽9 ҏ��Y�����)a8��[�N����eq`V}��$��R iK(�a��j�U�hd����.i#v*�R�V.o�M��H��藤?6��Z�AcSn�(��w�����%�-dmLp�"�S$V���
{�y���e�$�?h�ȣP�*���$Va8V\D>�R�a���q�btr� �I9� �R2���ph�a����Z��7Z�@�Eken ��r4Ax�Zb���T�K�6����˲��{`�~���x�'�����Q}��\���%1ȭ���z�JE���-��3���!��	y�&� ��K���6$�Õ/����[ZaޫZ��M����(r~�E���ч�j�+F�>t��g�<�]��T��`�Å(�u���bL�|�-����W�z�y�ۓ����7T;�Ż:�����6z�3���S<�y��ǽ*"��@���E�r�iD�U�_ZX�D�(���_E�-�g�^�^F��	W��&� ��9��}%��0x��>D4��C !�O���)g���U�)X��ⳉ��^�����:�@��A3���}� #?S��\'��Y����&{�9^�{�a[���Rrl������G����(P�|�W-'�� 	�%S�}A�S�B��"�f
��B6�%��Ӹ�Z�k�G�]��,G��`R6:������	��(�݃-z.o䭠��J�B�[��Ԕt���FYH��*x�U����c�0�
8�d�C�4~�Mr��s0�ae/�H��c�0�<y�9ճ�K�YƟ�F�x*����?N�0P���9	�{��Y+8�F�k�G���.V?��-��U�ģ'���Mp+P��h�u�V�$g��Fe��h	�E��|x5��J ��>�y�=���E��Z�8�b�B�MG/�oczG����ͱ�	\����kуO:�#��a�[p�/�f���u����K<nh���b3|9��տjUK���=MD�F��$�s����!�Iᵯ��ҟ#���P��A�Z�g�w������>� �+��j� �@��Vk��Z�G���,��E�T�_���ZG��`�o0�G{�L�!�M]�Va��Y��D���d���T��m�X�p��A0�7��]���73PM��D��pԗ�	���JX~^�^`�꺞���O E��-�J;N�%EtT�K�5���"䀍^U׹WN��DL�b�M�@�M4�H�y4�eT=�k�	�g
��TK*H��>�5��4���3w�2Z����T��O��7e3J��̗~]�16k�d���:��E��o�iu��|��;=����0A��n�N�6(�Sv�$ý(�v}
/�;�����C@��q�G#�E�	������dU��N������m1�캳��E�C�N�J�vvEd�T��W�%�����.�^}���YP���2)�w�"Z�6a��_Mv�N=��7���.6��g���cgP�{-�d��s�T�旾���+�*�����η~j=N�8!�X/`��5���M����B�E'7'O�iTjc�ұV�}J%��������g���_��'�d(��!uxjO+_�����Sהj�W䟴�c\��,��;
���}f�{l{���c-ʮ��2��8}��씷:�I�t�AK��M_i*�mϙ�*�V������,���ݳ*Q��Sf���:�!�tj�G|9�����ln�l�y�����-�͕"[���k�Ohj`D�p���p3ELs�
�?6jW���(F�@%�fi�iZ+�nk��S\ع�w�< ���JC-K��C�D.�����w<Y����\i,�,,�G�;���vcJ�;|�Z��V(���V8�1L����׵�{����$�)��uc@�x���7�˳jeZ�D�n�|Sh%;\��f���y�%	&��L9�Td���W�� VJ$��|Bj ���,�����R�mJ�+XK�ԅޜ�Ɲ9&�R���¥ac�cw�
�r0ٵl�����*�p�C�u��2r��a� ��3��Ϩ.8Sˣ�)��������g��r}��J���A܌ Ėؚx�!�qĮiגC�~3�y>l���IJd44R6>TD~Hfz9V��"�̄UV�}Of�j�M捘:ӎe��Ҹ�:�Z�MJ����D��JYnz���PoxY[Gq�O��@��4w|&��̔�z!�0a�RҰ�{�&�*�%�>P���+;m�m^Ɇ��1=c��̾�(�����<<�I�;:�*�!x�&����"ݙ�n���??����`<��U�f�*9>Z'���:�K�p����b�o[}/���w0c�to7Sn��Jc?�8V��vx]�Ӊ��رW��'d-�bq����҈@QQ�	�̞
�E�j���8Q�7�m
'x6)��%�3�/1��	<`*�!�n�G�d-1����%�x8Dt�5���-
\�t�r0eM��!��ܛ?#���G�v�s�:���>���*Ic��rc�Į�����n�>�&V4J�ON����Ns�b�8'Q�ij��fQ�3eҥ�7{��͝�n���xx`D�k�Z @"St#� �C�/��k{�S>�����Yc	��!�
^t���]��a�-�e@4���r�9;A�z�Y�q�Po�8���`r��p���D�|M��u'��\�8G�*��J6�l�/�1k�U�֘���5�K*n@�_b���u� ���F(ةXC���]��J���e�k��.갛Ӫ>��V������u5G�Ƽ7����	���q�0�FV�n�h�������J1�z�KM}�7m	)���[�������c=�q���&�<j���5;T(�E��
�}��t��V�D�ӈ���=����*n�d����{�Ǖ����X�R�PA��!b�r��O��rvYP�j|K/s,@�P�2��x&�n05`'�d�H�q������\<*9<�`��ܼр�i�����|�#A��ɕ���1�>�r�%�ĊN��D��Vzo"#	�~����Rhh0[`�����q,ٷ��=pe0AFMa�N�
����U��k�N�I�<�<)��u@Q�	Q�
�t����.�^�!�\��G[���d���ISmF�s8�M21�9&31�"�݁N���O+h�p�OE�^���q����@(�O��;����y3$�+A��0�B�B�Q����a�tՓ��BY3ľ���!�r�F�n��7�S8�`~o������D���f$��V�}�B��p�!��<3p\���&�\B������,FնcFRO4jہ��q��p��<R�� �Yx)V�p���P�Y�f�X����?��7�x)�ݕIs`��ū����	������`uӵ�������5�O̊�%�d��kͼ�	3����@`:�)��3ͱ����*ԉ�L� �d��~���cW���N��y��	��s���lu��u�hY��	�܌��(�G/h�}&R��cB�{�ϖ%Ǫ��*�� �س�՗�g�� 8�H�XQ?{�&��~���@��M�C���q�]���lu'������s�<�D�o�_�'A�p4ִ�Gk92�_S-\S����<�� �;�z�Px�RM�;`�I+����,6|E��"`��8��&+�N��ϧB�ֱ�SPÒ���CɎ�.����8����l���+������v�c>���<���m\W�e �?�ŮTJ��c��3�W��l�Q�%��r2��H��"b�d��0�$^@��\�#K:�a���cZ�G&��`���@��T�L�KV��JK�<32g���Î�MkN0g �����q�|6�7�������#;�J[����P����C�5|c�p]�<\��,변j%���_l�?�A��0NRm�i@t���W. ��T`d�N�C!�l��BvBr���������ؼJ���>��CpWoT\������_�#8&��q�)iǺ;om���'�����MO`�r�MY*��{��
[���x����WRXS���>b�kM�x�*I3�l|#�O4K��c���ߡ-H���&�|�b����j��	s�,�9�ؕt��u[��Bk!p��/�n�'�L?����	c��/���� ���a������c� {=p����^fx:�,�q
���Ro���t�����p���
�sT�o����^39�ƣ���ej�����f�o�l�H��PBk���(NYdK��g+�z� ]��8ľx� 0|
<u�n�Q����ٽ���+��4���y�����b���|�=iY/JIj>��ý�@����q6���d)`h����WeLS��=����/6�n�x��QB>�\���Ck
��J�<$G���8��kl�"Ύzf��g��G�M8U.b�Bl�?��V�C+�/�R���<�2�솆tcƩf�f��T�U� �@�5��X�]�@w����]�?����i���>�i�[� �ƙT#��M����=~�k0q��%��*E
��}����L,	���AB��O.�ؒp#C����1�xI[X[p��� ^�hu��=43t��u�S�G>7������*:R=��X��g���3k�k��d�2�N��qM��b��S�L��IO:Z6uzY$pW��,� خX�' �S`u#�g�ق��bĦ^X:�G�M����9U�B/1�j�b�V*������*������f��=�K1K����{;�dV�`� 8�̫��`7P� 2MKk���〪����`� �z���VQL�����zu��*�ƚic=��D�����'���XW@�����%4L��1�Ҕ-�l,�֣�E@���ց�Ʀ��2��7֙�=(|��v*N�P~�I����Gw��D�=WN�-ڞI����OdV.��M}%��e���~��b7����@�3�1��g|M`��>���!����J:&����"֭�Ć���?�xbn���G�x���A����རn�*%<�F�^gV�	�e�P͍������թh!řͤ�3�.8=wU�ˈإ+�B��R��J���E��lew4�_�H�^�WP����s�0�e9V�w�Ww��
o��(bhg�ӤDdkO�lz1kKo�>�����`�i*3G�(JN=RV3f�I�M��@�,6�yxE,vr5w�g� t��8ST���w,�ñ�4�A���e<��׎�'"=S�**��<Ѿ�T��:��k���������q�KqU��K#p'd�7��LU�
�Ι`������?�'�NP�=�+�zǉ�B���\K��$^��D�)ܑ�	��k��Z���֠�W�ӥr�%�/_���x;���,��p��]�wx0ᣲ*������ �F�?�1�w�$��t$[�J�"�Ȁ�)���Z�"�1ڜ%�V�]����V��`�6-Ö`��Y���UU����x,�T���;�A\m��
�ZM�2���T��@���d��\��"���ժs���s>h�[���gK"���qB��$p �,��{�Eߵ��]��*
PUϮ���^����v`U�Y<�Ee�-Z������8��Ls�����bB·��L%x[��%Y�P� �tW�)�,j&���[���Vz@��f�q��Z���N�FXh��/�a6a�X�9�F��Q�bW����ans��v���O����W����	~Ϋ���1�&��A����e����J��ظ����X߹�vwB�E���\#��[�cs���4�	���ekZ-�z'/w$�Ά�T�7��T{o�U~�dl��ϣ��ƋG��p��y;��HD|z6X�}�))�n���a|�(-�I?*ݱ������f���5��T����cQu�u[�S&@wo�S�ң�0�Ft8���ӵE���73M�N�H"�UAp��n!`H����&E�.Ơ����΃��M�=��q���GEa�����0�#�� ����ׅm�w�I�ŵ��嗢:�E�PG���㎎pn6�~�����}�@�4�u�����.�RC�w%P�.�7�!l,n´9�N<'~������o��"����v|H��='F�D�ү�a-�M�_���! F|9;�	�*�g<�oV=�C��Hrz�&_���u���j�U=K��\6���?��B���p��#��6��է�hܶ^��c�g��<5��6��|�|DnU�5%ls��qbw�����m�?���ꉇ�&4��ns�#�׏׵�jJ�C���gKކ�� 撝�V�]�a� #�=t@( 
@�g57k�&?�n������Ɠ�m#���I�zΠ�"~5���u�����|�x� �X�Cdwxw�v+/j�6�{�>!~��fhA�t�	�e*��n���$F�#��sdƬ�EA��� �6�Ϟ���.���ǽAԼO�PF�+A�O��(��Mo��?�%�槺T*�o(m0K�^zS)��/}_6����Ʉ�p�̶�B)�_�TE6t��u��j:G�'��+9�C�N��P���u�}Y�J3�L�P���yy�|l]��Vex�I�+?� հr�o�]�R\�ے%'G*w���s)�/ݥ��]���W�D�j����K+C ���$����:n��v��*��z��l�C	������B��+����\\��8N���㸖=���g�>��Je�I�T�)5^�"��A��� �)}����.i���*�Ztw�g��0��Mݖ�	��܌���-����K{��N���T0_wB9#=D4x���M���_�3kc�v�@RlB
�œl���rS ����6����-���U� �.�O�:Q�ɼvK��8��ɥ�ij����� k�'�)|�'#v�3>qd��R�d_�O/�%)�k���I%Y%BQ+P�����<��^�%��5T(BT����:=����R��N.ë�G��on��o���������� ��!��Ѷ
��L_�ܭ��w��4�$} ݷ!����H4�x$
rn)�0Q�'��Ϣ�$`[�'Q���ać!�2���jǤww+��]�:�vze�oGY#��0.x	��3��~�.>Q���Z� -^Γ�ZL�]�z�mQŊ����h�(`��Oh��S�Jȫ�#6)�m$v���T��� �d�7F�W~H�
/�R���=�I���cGG��:Iwt����gd��뾖8�[LC�ի}D��N�êt�dq=��{��N�2�_��Trw��Փ/^C� �#�o�Y-�+�x�D�`�!���$\|����>>T�b�r�;av��`ė�
b�l��iϵ��0���ZZ��3���+CT-���{���6kF��RD7Q�m��E8���;��.�K8�(O¯J�6�2Ⳣ��c�ja_8�����M�t�nT�ѢƏ�~�C�.��	k+�����C��o?����^]`Q6����wVq>�qSd�U�D���P&8q5���3�?�/g���*,DR��+l�l��~�
��-����� %[�Rq����=]��-'VH��ݝ����G���^�T�E��ƗaV���k��C���d#�Y�E��>vqo�RU�S,� ��6k��A��74��#E��+�������u�q����H�0l���-r�l������Q�^C�-g-,�9#��m-^�(��\��w���$��;�ݐx8Gހ����Z���%����ο��!��-�����B���jlI����'�	">DZ��un�a\~��S�l=���w��̆�'�_`a���[��YB�\ޓ�&F�b�9H&9El���[;[�P}��<KUv*B;k���� �py_���s0_|�#���Lx\�{�K�z��-+� 9?��-<��g�|(�}�W�rV}1άdN͢�*(8]BU�BB}Y)��޲�k;�w]�_�I=�� J��$�į�(9����LnW�J�0�&��g� E"b\��V��W�����<4� {	�P�!iu6�ΒlQ�cx(s~D���^K(����5��5 -1��A�$����T��"ə�e�hL6p���fH��4�?l� �pbW鑽�u	��t�`��\z�'7hl�^��b�ق���I���a��L���2 冨A��Z�?1V,U�c����	�]jz����&�|=Ժ�#�@Z.)W���q���=B��ɕ{cj�Q_	����k���E���L�E����r"�jk�0�rNp�Ƹ�ऀ��eϿ��/8��?ok�,
�	y
�&sNŴ�F���jܲ�v'`��4�q�-O�ۅ+�v�8���K?X��e�6n�ү>pp|�{<������5AZ+d�Bw�~P�M��Ŧ�?�MZ�l�O��7��~'w�!��A�8�E�+&�9u�
�y��d������A_��⿮�]�Ťn�2������ۃ��#�'�T���^��X'�v�{�kP��f{����X"������.���?T�쒲��v�2~�`[��ݖ^�~���:F�9�q�o���H�
�$D2-�C�[���f��F���#y�3$ҁ�e���]Wo�{�YP�M�D7�>�!��"2u������y���v¸��c1n���	=L�:;�')�ZKJ�?zYr��	��ʿ����Q�`�1@�'��$g:Kߩ�+�.M��O}�K���,r�&8��νSy��7^!���*حA�&��-�?z��k�!;����O�ͬ����fcӢ��{���(y�E��t*z�h:�þwi���A��j�$�̍�+%����z�����ϸ�����\^(�!L��C��ɏ�;F%�P���߶��S�z��~�I���X� ����-�79A��ѳ�D�_���T��Zh���#3��&�	%R7��X�!�
�途ډK^V)��(R":�����S�x��}9��>l����E�!G/�(LY �y�^eWCC󏃽�
t0,��{sP}��^ۗEm
[�6����i����vS�6��jt=�^�y[�\�@�}7��-5��n�t1x�:��T�\Q�Kɫe�h�	p����+)�I]�`�yY�an?(=��q%[Z�UFf�яb�t�WP���n�rAB'�e6o|�"�Q���b���ߋj�>d6,��wW�6Q����P۴dI�o�0E�5�:[��mNr�\H����bs���8r�6	^�m/)1ݚ{��TÄ��t#j��l��qC�y�;E�p��D5�ӷ��o�@l�z[��Lp�#Q1��H>����4��3�����N���=�2�JvޣHdL<�T��τ�I���F��;r������^�_��hb?�߶5˃_�0�}�q7�z�l���:JM���,4{��^�%5M4��"聢�6Ҝm]�= �Ļ6�(��ξ�FY�x�/"z���w����}H��H��vd^�ľ*L�?�	G�ł���ܨ_�� b�GuB���3��ru$K?���_W
X���	d�ٚכ�=��v�٩�9k��RiL�+������Z�� ܛ�E0x�.�6#��q�yaL���y���T�G<����#��.tl��?�7f#�!1&���N��q���hAOa.��N"M�=���Ac���5B��.3߳��)=��v"�5���$f6���Ʃ�.&q�;K�':��ᢕ��}���H��,���6��oC7]Z��#����5��J�,hAS�����9ۆ۲���<����N	�"W.����i9+�(p2�֝�_�x|ou5^;{X���.1�V��R� #�{�^�Kۄ�am�y]�{:3Q�����������f�l��'����˒�\#��+r�~����<���!F=#���~��\b�G�ʉ7u��>��:��~�8-���v�΋t�P����@g���N���R�d��O��<�
��R��Y�C�#�������/c�Z�N��}�AXD*Mڋ�'r`�n�ڒ
d��d�ܱ�;FZ�c���15�J�GM"��\�ܕk��d?���*�b����B�۩�Y��+��;a��v�7x\����Ԭ���U�&9�!�
f�����U�i�tח����;��	

�T7߿ɘ�d�w��) �As)���}�J���'y�Q{ˆ+�4���������8ē���o)i{2DM@�'����0�=vIo6O�ب�(�3�g25��E�~H�1�L�Pi�����w���M,Vʳ1mU�O3��C�gR����FD�U+��!(�s�u3×�-�`D֕A�+	�:)�ǒgZ��7FK�:f��e}�������Z�SU7���ΰ��~Z��܄Jz1��,���_�y�~�z��G=4���d"�~F��f'L��Йz��!�3�������؊ f[����a^.���UY�����95���Ka���-��,Cc��z52eG������������D�{��h?�(���2�^�
 IV�+6����>?�!7W�U��䏗2�/��bS�4�a�BL�(%�HMԥS�Bwq$-j�`��?'z�V+�>̨�����A��ωΖ�P���R� J�Ô�$&�6'�Kn�tY�
<7�-�vF�b	{��亀�\�xP�f.��>�!��1똳���q�8i��>�:�Q���Ƹ/�P��H�f�}5�tQ��?�z�6� ��E�>��Z\��5�*u��f���H�c�6\#�,���D](�<M����b2]-^$�d9ן�o�Iۅ�����;�w�F��L��m7M�+�d�?�!ҚR��U�ݠ�Of��ts�Q����
iR�%Ρ�BUbX_�b�-�r�Ct�o�����q!�[΢~BR��+�T\1Xϝ<��B�I�L�P)>��4�3�%�}��>e� �[>��U~=ESk���u��|��d�=��XXZ�q�-�*=�r{D�G��@>�%a6��ׁaf8�K�$a�f�jA�D����G;^ڍ{��>�(�Sp�)�0J��j��('�N�d0��I*���?��a��y�����	�:���4X���'2� �Cs�<���$�<�s�&�ݰ�M�kG�y�s�1�i��5�,	\K������C�"���at����Ȅ�1.Κ$92g5+����eNJz/������/:��C�k�f�/�[7#�$�p�%
�[#�K����bDY}h�Yx��Ԧ������y�f�yq��	�3�l��$�U�|�g��r��<�,��H�jG�@d��2�&�l�Ƭ1{ƥm��[mv������V�}-ˊ�^��eT�B�ث��xo"�ny��𻄹@3(Dm��ǀ�Xml�����b�t�!�y��C�����(�=�O�H�Z�Ӵ�R;�c(/�@5��E<v>0Om�Ղ#��\4��b��q�C���*Lv��C�k���\�,��`�3�jNZ*|�Zv�YT&�Q��t��"`�7?�xbd�ȋ�Ư��ɀ ���7+��������E��+�^�։rexD]끯;t��q.�Q��|�۴L�l�[��/.�>}_p���\��sA�]3w�s}#'7M�p��H'{����h�c���j	a�Q4L��L�,S���Xċ�<6�����œd�𵴐��=�-{�p�iQ&η��]0��2y�;�f0�h�^��]x�/:b_��I�vǩ�G�Έ�a?P�Yv�˙ѣ�� ��R�`�½���(�����!�J�����C~ɩES��
a�1e<�Pc.@��#�>�@3��?�q���)D�y���%�PM��hT���*]?������YV�m����P�Ad�AP�u��{R�f�8�|J.Y3`:;cF0\Q.D�������}�ߦ�\�_�X�<�SK�dL	w� �N�ܪ~��'{��VTȴ�����k�X|�
��s�ᎹUN�4���
�OYV������̙l�6�w9
��}��׭#��G�9s�ļJd�>|��&��g�o�q�2�� K�QU�����e",L'�����_;Xޥ�ؕ��� �e+��zx<�o*��UD6}$��u@%3�C 8zX����Ug�u&�����&S�������T�@.��Я�I؅
[��%?0��`�Ҹ~Ol���?P��L�M��r���Z*H�Q� �ΐ�C�y�$�^6���T�i�>H�ʲ�t_1�����:~���Q�(�-z�h)�WZo=����$�1�>�d�6pS0�t+�-;.&�Bx�����0��(e�>��0�A]��G��4�N�q����s$&� .� �u�B��MO8`�s�������&8j�]�9v<XL��I��4�3%^-�%j� �SVK�L<R�J�U��N�Irʬ�s��Z^�8�7u�ض9T�^��P[� ^M�À�E���Jy��P9�/,���mq��8��i *4c��Ǹ5 ��Q���
i��,ռ�f=x��o��nm�T)(�ҡ�#����9���>���R�	��(!P�v�������5��1H���N��d��8#�u�������f�{S:1�	�'l�u^5�ۚ�3�������%��i�=vr*h��%�
م�3�԰^��n>&�$E\/�zF�a�j�8�
�9�|�"���@E���8�lp�����;�]��i=39��-r(Ҩ<���<�5$dTI�Dp�nz�k�rAx�˯S�B�;g|S�)_�{��q���wx*c2�\�mѩ�=
ӝ/n�T�=%'�5�BS3��Ę]F�k�9�L$F�&b��������ǣ�.N��ZQ�D�U���Q��r��fa6u�5�����[�r��%7�f�:��@��h3�PZH0�PtB2Yl��j��;��pƶ��j�z$IL�R�j�)��%�����>�>r��{�4׎bhN��	�,)��õ�d���gC*W4wQa'ót���j�A#ļ����<�<�z�U�>]uW1_-S�]DdN
i��I���^�+��	���<t�	������:���j� %VI	7;�j�`�������R�q� ��"kޤf�⼌���jA7�-�H��WVG
9�1õv2��ɛC�ܔ��1���	��BTVJHs�����T���bt�OE2��iE��+��h�F���)>3������>_v����:]��(k� ^�9��@l�	�(�Ȥ���p�;�k�<�L�5�uC�������[��٘\ac,vf�_�sf�ό8��v@|�7�kS���޸��=!E�>d�qpx�of�hF�Q�ɖd���ZA���q0/��l��r��pjs�+�����L���
n'x��>TS2�H-��<[�;�s�����4L��0)�w��,FG��S�L��Q�f3��fX����'nn��5xƙ�N(i%�=C1���F˧>�\>��t6��֣�n�>	���`j2Ӳ7x#�^�,n9��>�E� �|��q���J?�+Y�x��C��Nl;��������;�1T���}�;��[�|�I3p,�X(��Ŀ	U���0*o�p�ȗ� 
'%���1�8��B��T��>AM��g,K�x��Q'�Cϲ�Z�p](��� GE�.��jD^�2�9X�����ٜ�.�F0�}3�G1j��B�w�]a��Ǻ�c$U�{/�����䖁�M�-[�M�O�B�"�A�M>f0jSc����ъ��j;%�	��d�P�s�&��;櫥�x�%�+ �DM��Qk09h��X��$*g��]X�J�Zc���>�ƒ�JyjRQ�8�ث�#��O�n��xz���q0.��d�s����K�]f�rL�	锸S�����-�{��dgl��Ĳ��w��(:m5�Q�df)�y:��lSôL+�X�����[��u�{�C^˄l]<e��p�}��ֶ���j�A���oGSԶ�d���?�+�ŋ��c�+�ڛGOS-d�1�ܚk�f%�x@f�l�Q���m����d�1�j��~�Wѻx-2��?�rg=��k������{.�m�'V;�����a1/��a�o������J���"�R���#C�n���P����h��4?_�f�d����G���)�=�-��G���=��2S�Z��1�ie�r �7rf�T&�U��b���t}5�|�<�޴&(\�	]$�>%��▥�l0���#̝�3�yL�����-���/�?�N�ẵ����Ut\l�J�X�z��1�	K��X��_:]���=Y�.����5L8`9LT	n1���+~��U��aW4���Gn��gH�dm��Ӊa�)���ȯг8�jh����9�"K5h��^��Ap��(�'�'��Y���c�|��f���u�s�^��/U��j��߁8��>�2�rӁ�ݞ���G��bN���Y��ee��~�C�ُ��wi5� [�]ȱ|�����M����Q�$���y�O������K#�5�0���~jm㙑��/��g	��p���ڂ���Bc�gpZ���P�t��n�+�\�v�|�j:�1���]BO.��PB�ۈ��@�0��U@^����o���H����W�7���bgtx�C�qK�@��a=o�#�M�)�8�۵V�W�Ԋ���}[��Nq�z�A^ʧ|�9hX7�������;;#�C*��d|�"�\:=h�<�:|
c�Fk�r��Rc�q�6��+���F7a!��	�A[�m��2hei.��@�ZCGoB���(�%vZbE�89������jh��V�v��6�j�kEk%�	}Su����(�X�K�;�j�cKg!�վ>��<7�k��waJ$�k�:T4� �C�ƪ>��l�g������H�s�� (�%a=��a�l5��h~����tӔ$�I�;o2���h�u�A:K�$&��8����ӯԩ���|�ĺg���"	-��(Ԡ�WU�����7"fT���6����γc��eO"�¤r��=�|	9�-�'�Dp��EaV�e���S���I���V6A�������������^E�\Oi0�)$�1�3~�k��R�{��!Xu�O��+�i����>O"z�bԬ��w߽�^��gۉQ�kwˍ=��r�pm��s�SF�n�wfO:^S�h�kyy����(BTo�	�sB�& km&�{�n)*���Z���	'��ŗD��{h�I�Ib��I{+}��=,�W�I<�N�X�������F�ƾ�/yC-��(B��2|�����ߗ��q�`;N��WpY'��s�W����/9�� 6����{ݣ/�6�↰OL��Nq���x^ͪ ��N�礤<ݎQİޥ�a�8�� �p;�0� e�A
*{�msG?<%�hX�¾;g��.x"L 9��UA�*>c��ISm6=)vPb���9�>����G���{K�F�l�j�=��c�5�Fy���Qb�MƘ���\jd���эi�7����խ-}詊�;N�5��|�E'�r��u�2�	�yxbK�����>$�?_����""�(=f����6�ט����t�Ud�D-(�Rѵ�C|����A}7뾃��v�ɍَdﲚ�������7B��e-�՘m�5A�j��u��ί^�VI�-�)k�D��_f���,���0W��?PE�\�:��ض�����ϳ���F���`��'Ͽ_�I���vk��+|�w<���W��
��sh���7��$��]������mڕ?dem�ϝd�δ�Ak�u[X�a��ģh���gj��=fwRwV~���I�Yr��w��3��@��Y�U�O_7�k��Tֹ��4&�5r�:�[z����~��h�W�p����#ͮ���G���Zt���s� �Vd�s,g�r��y�d;3�w���t�Q�]�̹�j:fm=6JE���F�Ӻ`�����d�?6X����8�Ud�[t��#�u��w�ݒ��#H-?����F��i�K�'s�~_���>B�27*���MЍ�҉���
/��^���V�,�����FkO
�b���������/�^���_��C�Ƿ�T��~�ޕ�~���_u.�,�)��(���j��fx�O��f�BQDQ�B+$���^^��5aW�F�k��%�����E-a�Џ���(2h��U������7��}�-Jm^M�~�@���T'����z_HI��g�-�[8*�R��=�!gG	�-��څǘ��h8ǵ�F&�������[�F�4� {��7��.��d!��pY���nӒ]�] a�[�϶5�׭gJ�y���!�kˡn	�}|iH�@��؃5��U2���pؔ�x�,P�t��c�"p��Ik]d�M�~��b�4��R�GY�#�ɮ6Ȁ荪�	�4ټ�ShcYXE�]"l(釡���Z�r�*VM�1K<����WT!�Y�i�!H��ܾ+�XD��ѩ4󼘈�y(��<O�1-O���� ���h=�YV�컧��A��x�:�c"D$'q���?�s��$c���1��T�fmr_�m�M�4F������d�E=+_�}�*_�u�Ub?j��k�ޒ��o.�)Tjm3b|��*��l�}��&㜭�K�i����8G6�>��BK�̥�l��4��l?���Kͻ�W%�0'i����D�#��y��\O���<8�\"�D��N����G*��1���g�l�84�j�0�xX�Bo��N�����_�K�Ȃ��?�qC���┹�|��B_(�I��cT@���;~t��9N*���o%V��.�>7�|ΦЌ�8���ەU�g�M��M�|Q�;�e�#��N�]��N=$�项�-��H���g�BL��G�4��#����$���̈�}���Q���ewy�W�$�F�Vu#k���C�y�zAh-;5(:���k.������{�S}�G�6RxI�N-�cQ0ǐ���A�wC�7���㗊�ճ'.����b�&��e�����B��* a(˟Ȫ��-��S�w���}JG/������Q���q��?�0Ylo<S��`��7I���
��v�w�io�<g�js�JG�Bcc�� �!���x��̴ٜ���L��nx��r���$�(�@P���b��{����^^/U[�\�1d�[򓝖p�$H%�bh�V�� �Q�G��	:S�{��d�j���m�;�[bɳ��d�kA��f�2�r�0�|�aq4��バ�Ȭ)>����ji��6$f�3����n�'�ޢ�^����I� �r ��&�F0�S]B����>�ɜR�R0xӐ�"ޞλ��ӖC�nzD�(�=^�j踌���&�lDj���kT�A~�t��_�
/8E�$62�3���&��������(S]��su��'�9߽(*W%�Q����_'�M��r��n�����_���#�zy��CM_ջ&���$�>�:�?*Ħ����j��)��Lk��OwS��#߻�F�cHY馬{���p&1��'��h&��e_M�L�i�I���(��Q����S�޵���l�mhGB�.�-�y�Dԣҍ#l��Gѿ�<.�ץ�p�UX�~�D�����4��\��ꗠ�ߤK25}R#��mڲ-�O���R�C�@��6'zd�;�uk�.�G��C���~��K��R���荒{�zg��c�DA�Vס@�������������&�X��o< ��UR-�Qhm���뱇�ڠĽ���[�lCo(t�����1]m@���6�oeĵ#����	�"q�j�fa3qD�(�;%��==�@�F���g��]���ΰ��KCä �"�]Nw�L�)�S������M"%[��B$C��)�;
���aOix�VG ���)��D��*����˅ӌ���+��Vh?���7?<Rg���%��ہ�SC����� s��2/��A���i��ΤCV]_qO�w�h#*�+ `��n��=x�N�����K�xj��Λ�磝�v�w���=�R(}�0��x�S)E�;���^�-t��aO�zE姱3,�ja�
�YK�kcf;>���iT
�?�_�k�*�8#�>U/[m�i���OI�၄�'�c�diJ"�P����DF��js�ľҍ���0�hKK��H r\0T����)��@0~Ȱ�֝�'��8:���Y��6����viL(#WM��eygO���3��zz���@I*�ћx��6o*w*�#�-F?ƿ�[����q��T��r�Yv=Ѝ�����M�}k�Lx�A�zu!`�6Fs����L��Q�v�/���s��.���MGn[H5[偤_�]O
W�Z�-�xR-ۮ��=i��� ����ե'�B5DnEQO�F��8WKB-Y�g�f�dt|s��8Ul݁R�Ʉ�'a�f��Oz��	S-�� �~z%�N_�0�5'~iF��|Ê\x.��iP�QA���Z�f,1��z=�)�%�w�W��߷ �v]�g�­A����Eƚ�O�zл��|g�8O�X�+q��S�7�5�ۻ�"'�@������z����ZOJ���h�-���U�:*%ُ�S�B��i�B�>�>{��,9�4��������X���Gt�=��v:+jztJn��yT�^d�;����-���-�"��e?N��4&�`:��?[ �j��<牛�/�V�*p��*��/��ۯc�)��|7������JAzD����T̒K\GHq?B�-r���Vl�2Q�oU�- 9���c�s]�n��%R�K�2~v(��r���׾�U�T�
�3.+�
��?YZ�%�ȼ�^Q/�:�*ݧ]Z�p���s���XrOV%'s�����6�B@%���(fۺ�D�/Q����ڇ�Q.U�64�����p��b�!$�I��s �:cz���P�4ж,5�$�a4�I}�e/�(a���P�X���v���#S��@| /��))\Tf
	u�y�H�)V�(X@dJ��f�ߍ�M�k�=ɮ���;q�d�e���C��c�L%���0��(d�D�<�Y4J�õ�8���o��#��;~R�ώ'x�B9x>rF��t�����}(FoL�&��`�zD62S�ҩ�S��JK�}J��+�Q�n>���W�a�$)�h+*���\�1����$�xNr����$�aM��=d�Ms�w��7��$D�4�W%�we�s�[��ʒlzw(;�I���\����CQ�U��I;XuI$~��L�!&��~��3��P �j,o�l��
�����V�Wf�M�ǁ��V>w�&� ����_=�T�|B�Y&W�H���]� S0�tm���K5�b�_�"$#i\�R(�B�8f|ܮ��G���N6Z��Iy6_�Y#&�K��wh�[�{L�+N/˙ŔhH˞�u!#/|(��h��8�*�e��خ5HϴӪ�c+z�B�3p�8��C�8Z�> wK���\����e��k�j[w`u��)���r�W�%����_\i9z��#���Ioh4�_Z���T.��5�k�#\\���B���:/=�M\�q���r�V?��7�>�/S|d.�~�<W�~S֞���*�1Ԩ�#%aX�ZV,�����h�[���r���)�.����f&]䄩�R��&��� ��4j�rz��{�L�4��,ҍoȣ`,LPD�Q�V�3�8�!0ɰu���]�g��9��U�{�=+��w���r�8]�CYo";��Q��O��	��POĀ�)'�KXR��=}�F�)������%��@���9���8.�&��|��}��|8I��y�:SWk!1ct�-����*����|v�M@���p���El��NF�c�����c`T~+$d�~�졪p���fA!%@8�S�a�H�Χ6.��O�0}�`�ߐP�[Zm#r��i%n��h�Xj���	����p���Ğ�=��7���H�y���p�{U�B�F�)��ZQo�����k��禁�WHBc��x����렂�vWm��׳� \k�������}�r�0ѱa
l�lf���bX.�Be":t(��8��C�a�l�lh5M�"�\r�oԟ���̂ѩ�gv>s�j�S����5����ϸ���m��7F+}o����|Ԍsp�Mj��쵰a7٬%v�Չ�ɑ��a�>�<+��
[BR�P��X�ed
8,`@_���5}ٷ�3��� IC�R��Vƺ�]���� ���7}��,#��o(��fQ���f�͎a��Z%��N�X�A4���!��;�����1��@�1!S]`}��l���+�Y�k�+�\k�d��U���\~ݯ�p;փ"��҅���<��1����'~O������f\4�(�5��j
��b�;E�������ං�����8�hf+�!qd���P�ζ�fz�5�-C�l�����~���h��� �-](;�,=��j'� 54���a���QR7�|��b���ǽP�V�%�F |߮�	�Ɲ�\S��e�(5o3�޻�U�ށ�+����WBgk�+}���c�D��גH�v�Bo�T���>����?<�b�PBUc�$�`��q��.�mվ�ݲe�i��kA�4��^��j,�]��HST��B�����]6Kb1 ��9�@{�iFM���ߓΧ�Q(�
�&�(MM�[���O�@���uc�����nA�=�g2#f��K�-���)�i�ٷ@��V�#����K�|^��:q���Rx����~S��X�$}�9���
dq>TC�	�I���z1��KY�8�����qR<�.|�)C��~tB�7&]h��4� ��费+�p���ak����c/��\��$u
|!1���`LM���I3ki�l�Gq�=[N�|5u!�,f��s+I&������_�z��`Cd���F��g��~0���u��fF[+t���t$]�l����R\��Ɏs9���\����;TmKimBt�۪SD��G�M�Q��������I���`�Ӏ�]�y��x�И1]��ޝ�X%��#�ӥO2X��j�=������K�E���AƊ̽��$|�����&%t<�pd+���01��	s�6
��?���ܭHb��|��""��L��<��B>W:K)��
;�e�"l=:h���gEs�t�z�k
*׏�D��Q���tY�`�,�����<�%�l8�S������ぼ����$a:,?�e���[ک��Hz�\�]��*±��fh[���m�b��^H�-NG̀7��3���j�����v)u+��-3ᖠ���ߎ4�/0x������ �*���[�,��M.4è-	��&a��tZ� /��w;@�2
B�Z.���3O±���2�L�|��T��C��V�L���k����.{4��z[ʶTp:�D�Ik��S�Sx��ߴ�~���4/ ~p�X�!��3]�p ��Q�|T��ل��bK��(b�����Vd�0��Z�}�*:��_��U+l�S\���t�Y�Q'ǝ��4��2r��+a+W���2H.���z�
:������R���'�b��n6gq�b��mM�Ga���$m�
~��͆�m9�L:S��T��}(�_��:Wg���G�ȲpA�g��jo�P�:9N�z�����:1a�J^"���0�/�9)����-�SCԓ�]�d���(��d�4T�%��.�K��+�$8�?���^�q(@�
(���[_���.�R��λ��&��=��1�r5����j��q�=xT�6�(6 ������U���*f����/�o�h(�x�Ú�����^����mL^�G	x$�K���s�~�����W��"u��e�����bp����J�k�x���=qy������J@v2u�͝:�ь07c%�c�~��V���'Ӝ�-��盧Nj�=��)F�{QO��n�,���MQ���\�T�)u�b�����-����F_��t�-�=o���"����A#�ПN��y��tc/�"=�UQ6p�!�J�����V�}��q�n���^��Lַ�5X�E�;��ΝF�����tWR���ac��W���P=�W@e������_m�׸�"�/�G��i~�'�.���Z��4�����7;��滭���� ���a��8�q���N`�4'칛V�"��-�n�"��W뇤�l�R�R;�h�Z�����><l�S�ͥ�J��mK����P����!��v]��
(�UNb;f��ߚ8��I���a?��})Ąd��ǎ
D���JI�F��y:V�H4��h��t�/�7���c�4�	S0��?&�qx�W�e�9�C.�ϻe�x|�G%�n�Y�Z �*�j1�pZ!�;h
�ƛ����;W����ش��j����GӫR~��`�2��x�Qk���\��Ζ�fYX[-���?���xf�����Z+�,IGWl3�^	�M�}z�E��Ӓ�p�$�sfH����`7���-<и�|��_�!��8q3��U�xK�4]���+ay�{��H5e; `j1�I�е��s���6���V�>�6��(}\�1�ܛ~)�e�S�*�I�;L$2@u��8��O�O� �ֶMy��LѸ8�2�� eF���� �"oc�����͏��ud1�S|vjZ)��Ǻ��������AFC:�3�F���A�E�q��_��\��je�����p�sH�X|�:���w;�Ё�a���e2Q�Rȵa��e꒾���-?|���N4a��]�.���/��X�5_��i�,�`l~�*�N��nd�[�������5�d���O�>�Jfב�|��i����05!��ӸZ�3&x��}�MQ3���xAÅ�JRzh���$0#}��`�&���f���G���A�F,0�����PUp`��n({d�>�{-��E
�����B�-� �1�]�qg:��;����oꡦ1��[Y��J���lD������TFw�㈮֭6�9ƨ��A��z �6�Ѓ�x�l]�<���	�7�Ƶ��Mj��yO��-�F[L[�FX������94W�y����g��/>��Iz�w��M���v�<��)K����m�{-�UZ���d��>�d�O�Fh���K��nl���*a@B�=}��C��x���˟X�W�>���Dj���j�*�{|��J*�ކov�x,,y��:�|jp���(y(Cm��=~��$~�,��ש��pq�� q�v�
�~��6,�>� >$>���ZC�(�|'��v��,��7~<�Oc7�M��ވ"��	[�?�"�o��s4�Ԓ5�0�3m����->0������\���^G4RwT��V�="��ǹ�'����Fq��jI˱EW�m�/ �`�������8�2�n��QF����c�*<�= 8�DD�� ǰ�qκ�6<W9�ݛF����;�QB�Pt��s���"U,kYڇ뱍���)QٕE˧JԅKM
���o��^u�p9c�,S ��u֪KYx��i�<c��=�"��,��SGR0^�8C7�*f�^�S��!vX���7�/�݋3S̓R������A�������*�9�uJP�Dͧ��u5}tS\o�D�m%N�^�V��`EY��9&�b+,�I�qu��*���)�K, "��3<6�l�0���e3*�[�|=$�&n�z����,�bGo({\s�ָ[�";�"a�ݤsR�yj�3��l~�AH�I���^�C��?�Zx��ȯ|"�e껾U��䈛LsRvD� Q"}�9EݵL�Z�	������ϕ&�:�c[R˫aͫo����-4!�2D�c��<�Ĵi�ټa�e�^S_�V��ܯy��L�����˥�5'V�Y�5�b�����52JY8�����lR���ue��͵�� ZC�L���pg6��a��G��Am�p�!��8�K����
z���g���(M����� �Hc�z��h i.�QmI	�Y��b�Y�\�\�]�g9�n��k��:{���>��c�aS������c��+f�U��쀎��]���WFJ1�$ף�e�1�K�X�@)�/�Jp���v�\J�!c�$])�b��`Wq_`�o���W�{��Ȗ�>��s��=�.�������4�(�p�q��DI2D�}�S�9�"�C�\�q��m �ӚD"�	�Qk�z���=��	8��������۽�FZ,bnZ��ytB�ݷ['�m#�� z��1̬��ŕ��'�~�g_���Ї�8J��9�n X��3�s�) aօ�L� ?db�t��A7��e;�:���%im���N.C�J�"PKiUb;4l�#IH�ѯ��`K*�
�a���W��+�$�rFU�p��I$B��`����L>APn�[��FM� 9V*+�_�O���8�d�Uf-�:i�	�ԅ�ƦzDQ�-B��}���3�4�8e!�.���^�E��w��q�[�a�|CF�lۿG�=��ߒ?�&��4��H�b|O&iUz��u��9�׀�������qW�m�4��+�zcK_`�)k���~jf<�c���kw�i��3}Uk�N�i�/,i�Ɵ�p��щuh�ߝA`R]�ffʳ�
!�³woN���
~�/�i]����7�[`�=��Z��!v#@3�~2H�Ռ�ۜ�M�GJYN��rʧU���3�c���<3n��#H!���k��XJ��	�q`j$eP�Z���z��ń�L/������ؒ��q����*;��,���[b����0�`�'|5��F�I�����+��j����H R��
������7��ؽH�l'����v
F�:-�����ح\U�l�L�IMJ�g:��5{}]����ﹱ���M�${$�S:�E�dL���N�g��*��t���!�t���&��Y�~�[;�f�o`l}�� j�(sW����~=fGJ�P��l$�����b�@�Qނ~P�6�P�a�U2�yE�v��������x��ѳxaL:���m��r\�g���v�G3[���?���A"�A�y�D�vhiC [-�(r�ld���/�r'�WŨ�̷r5��ԨWhv>6���À�H��%� ���zű�G�l�5�e�;@װ�5"I�B�U����)}+&����z���ѡ�`���S�%T�%�b͎�g��B!'Q��Ac�s�`�,U�� D��~1���t0���0C�����P��m�ʭ+�o�<Ț7-��(��e�ȕ�[�Xx��B\{D�g������X�?;1��]����n5}E��Hʦ���m݊7���^2��~"�/kN��
��&|�w� k�^���"C��Y�.���|y֒N"vA�8��ne$=�i�6*��"�K�'����t���6�g�jHrǜ����/<Si���?*�ځ�$�n����G��{4��D>G:z��`�;,T~�O"�p=,�CRWK#k�b�Ihg����;���H߯���oU/��}^�x���ׂt�D4�>�}|ea���vɭ!~��(.R)ґ�(�|5��l��b��C �a1½v��3���)������W�e�@��#i�E�r�����Y5���&��K����zƞ�#L�̜m<�k�y^D�Z�[�l�f���?r^�'��D;gVȦ�a�r���wxT�\$�MF$і�x��O��A /�~���^����KQ6��G�b��.�jEMbjIB�����b��"�~�����,�X������>v��P��/Nf#I`1���y�<-&�<�e�ʰ���u¿m�
�#Ur�jU_��(�Ӗ[�S|�:��dw?$wx;�xT>☽݊i��re�ѓ��G�/��[��|;.�	|��ݐ��E� W@+����x���Om*Z\�l�2����\���T�W��B��{��f�<�K�jvo8(`�*x���$���Z���?^��옰f���p��
C�`��?2��|_w�ex��K@U�z�������oΗ�V վSC�G\�'��lO�O�X$@��l�7�F|�l�[��"��R�W��� �4H��bun���|y���`��ɓc�v����N-v�bйꔰ��nJ$h������ε��)h	2Hq��t�/� >�#9�76�Α���Nǿ�� X4Q�(�%�� "�N�j؋�f�z�}#��r�ʎ��wYm7z��P�"}5L�-����IϨ`��� �A���SfyegiX��s�
��V@��2��b:X�5JI�򓼻��7�����ˁ����Zh��F�<=D�@�t@-�R�g=W���W��%Uf�N`��k[f@~dM�=�����zcgE~˸���WE^m�"�!�q���rmĽkp�1#��Kyx��%�h%���Bp��k�!�Zx-�:+K��%f�2G��̙� \�������(�?��R���rq�J��&�a�;�;H��ѫSQ'G�����TRJ��W���aa��Q�h��
���N�h�2�E���U�������{@#�ЃK���L/�����]����p=� |ت����XW�Y+c>���yP�?���{W�܍΢���$�/k�4�WC)~�MS�AJ��T��c�;]V�T�3s�yK��=:�3$��ݹɀE��e�
��3w��t��=���F��������bq�Es!'������c~�	.@�(�d�s��!rb�Z�O!�>{1���2U6��f�_�u2����P����gT[ѣ��>���}}F��8���ə#yPNݘ�uwt����[��^�P*���j������䮷���"k'*I�N�iֶD�g�Zi��x2f}	4�Us�g C8}�sg��/�B0���-���f(w����,��2�2���>���_��;{��A�z��ń])�1����z�8Hj$�-�Sy�{������Wڟ��!�՞��f�i��1��'�}��X�뾩���e�x�HAz8_�/�6q�b�ZY��h$ܬ� ��)�֏��p7��S�N���G!��.9=W�?z{���o,���4l����\ٞ87���;�;#R��v(�C6��T$ؑ1���5E]���
�(����_�zIRҬW�&��t���3�Ry�n�2OGȤ��Gi	�E���M�q�c���x�8q�C��f�FU~W!�M�N�EU�@bq�=�LU`�Z�P������ۮ* �W�t���oA�HB�aRB55�Ӕ�ee�Э	J�����^a�.O͚8�gu�6�wŬ.�{�g*�l�a'��o���dR�0FE�v�i��K���g�WB��4�����ܟ��aPFP����v���fX�1s�*��:d�Qgf�|Za��Ju�j�E�<�B���)�?��Y�i����1qGxIm���U9<�2'"YVC����9`U�Nm��F=��N�nf+j%�r�² d�X|[K�+�Ě	�W�>{����97ds|%�M�:�����J��=?��|�\���kc�Z�Psg`2�]��5C�Ѕa�,�Xl��~�������m�S���C�A���%�dތ���#l�La�3ߥ��ΐ��R��2Pv������O�>�m1jV����O��{Z���Ty�#qHq7ߛɎe2~LW�>�rR���[cW��W�S4�ؕ�4�ɚT�>��U��������^D7�F��&&�4M�G�|k�+Ȟ�廢�5V���u�f���T:�� ��<Fe���ŉh��M��+g�L4����"l�����r�F��j���V���sf'�h�<�8������͟	����^��R��"Cq8��ٕP��2u��|���Q����f��!_�}��k�i[�(��j�\&!�7����5XirfSE1ع����֑@�cn.�� �K8-�o^.�3��=+��ؤ7e�Z�A�W�`o���m�"_�U�AF�*t�?V��I;S���+hܖ^h&(jP'L�z,h�V�R>��]�"a�Yj�����[��maa���Q�񻱇�G��%-��GA��r��ϻ��G�m����/��e�w��l�5	���67���6��Obޑ��B�&���*Ċ�j�+*i�Q�v#��/*�܎,��j9z"���HK�X�;o�$�s�Q�ìm��x�� �|X�Z�9��m���-�h��`i;W-$u�ҳ#�4C�����h.�~��u�ᆙX��re��C4VP�y�-��ihD�]K�����x|b�Rx��Nߡݙ�0�ޯ;����֑�G�ڋ�y�����z�
�rg�mf�ݡ��J�G: �)͗��N	+�gi���.S{h^���Y.�z*{��8�hl���Z�E�I�Ѳ-���S���|�9_�R爹�&�R��`/;E0�`Ly
�S�7�2\F��$�Z�#�!$Z&�Q���ds3w'�uJAZ��J���Ҳ�Bω�Pn!�u9d9Ng�T]7�	�k
M����g�[/���N�0g2Jn��E��e���<q7���0Ir�OJ�5$�����u=�힟P�[4�P�F�S��m�����m�t�q/]��4���N3�.}7�G�Y@����{�f�J��wO¯����0��?D\��.�#�¤�+1�T�,\\:J˸�
uwo%��:�u�s�U�� i��'��l������#����)!����c�;ȝ�M�mt��HP7�By�~*�Cj�����-��M09��m\��e4��(��h�n,57���L~jR�<�s$��>��xC�9�L0v�{�j0�k���Ǘ��s�E�F�uS������w���l�^����7J_������Q툙��L<�=������u[c|ŉ��b��9JR��)�O��xУ	�L?K�yL��;wIN����/q���ց������i/�%S�n�*�����X�����Z�r�$>�H�}ҠǓ[5�ꃂ�L�5^����zy��G���(#<{�
lӄ���5��H=�̻�~Hտ������6�H�Bv�s����)���-@1�}*�����1<��YG�����������)Bd�r3����U��w�m�a8�
k����aS��P�fla������g\�(���!�ְr���:�D��}gT���-��gU�R�W5�5������Î&�&�0��6Q�!v����]̅�ԤQ?�mLBL��6��g;�"~y��l�����z�Հ��� ���LG�27�>H�q6�K����-~�/B�͹�Ϝ�e�<K,���g�< �X���H�2N��P��zH/��o/s���݋R͗�J�j��A�c���_J]�&^IDW�"�2&���t�ɤ��cᮺn;�&��y�����Be��%���u��>T�J�E�K�|4���D��p�U�tD<�?�FV֜ .E{E�^�/��]�T��=h���`��2�{g�)6O3� ZX�1!��+j����(���5��Y�|�ݒ�Ab�c3"Zҽ=l��������\B<�cO>NnV�˵�γmgK�|,�O7doY��dHK�`��a�s�L5�Em�W�VE��'V���~���k�w����ͱ�|G��Y�<�����B�V�Z�Vz��qKS���_�10
6e��|�nٙàA�M{Y�u��Ax�r�s��*n8�o#�P�e�=qy⹕Ђ8<18�,MH�U�¯�l�f���(n'�$�rF~3�?���983�������M�И�`��q�,�~)'�WR�wA@�ahQE��Д��+�ܮ�O�;�&�Q�aA5�u������[��iF俋s�n��hp/�����Z��M�'��X�9�Мgb��L��-�P���!<�V@_v�_�ɥ�~� �F�{-"5߉�z�0��sƪ��e���i:����W����y�ԡ%���Qh�� �A}X$��K��#'�8�]a��?s��<5������זٕ O�GI��|F�y���"@��XwJ�od���Uw�4�q������i���{")wW�o�Y�:��8LL5��'}�+vM���B���� g#?����$�R��k�/��|k*���_�}��O����~��!���$`3g1Œ��0\���Fb\%h�K!�(Br��xw�:���vl��d<��go<��7:�R��#��U������&8HS���jh>�=ƞ�������K_`���sˎ]�]-����m�hMǁF�x�9ێi^WqH���(�� d� ��+���J,$���.�c������:�Tp�վ��30��v���T��ܙ�TC�9W�.Q떓��EK\����I��/�k�8�������L��(1�'o)#OxȬ۩RwvD�ͮx�Z[����ҕ9bQ����{E��5�:��d-A�=zt/s�N̂�����G���E��ȋӼ��-�w��Ʊϼ���B++JP�^=�8�ȃNߣ�'����x�ُ�$��B�d[*W�>AqG@#-����6� �#ܘ?�B��Tp�=�Fϟ�.Md� �pUAi��jK�*�"��S�Ȣ.��d�qج�>���PO7�X�{	?b�=�A�s��	�J��姵�����d��!'��f��ཨEl�_�X�	F.�||�M���k,��	��A�6峉�S[�2��[C��A�+�)��]ǹ.�	��0�~5�+���vWL-�h�l������>�m fZ�Kx W2�֋@�4qn��������Xp���`>�\֤;[a"�q^�oBV�O��X��w3�!��I�������"B�:�nAvBS�8y�P2J�>�c�L��F�bsBR�����G�������g�?Ǌ��/���w	���h.]v�W��h�/F���j��i'!�ũ���nY��{�Ѩ���U�^W�z�� �X=�OևIDX��C~�e!.v�dt&�#L�tkI�r��"��DPĔ	� E�mdB��m��b	����0��;իU��%�ߊ�"�k�V�J矇����|�}%�a�;�q�x�s>�cwc�C� ��n��g�7��&�|�$���j�l��k�u[f������|�$����{�i�r��������[M}hQ���J_����=
:<�*�ى(�0eSC�<��G
g3D�6�Y�f/��e��ѥ/��G˘ԖOWD���=����.�se�Ǆ[2�Տ��!X6�D�$ǿ�P�P�ɪ�x� �epv���V8i.JߑMҥ��
�>�7]�޿�6/�#��N�Ԛ�F'�.�s�����Պxp�[X��{�=�Q�[����m�B�ʎߋ`�c��A��4I%k���I�3	�Y�ϗ1��~���z��Z�{��h������6|�G䁜���%!qƼ�������3�6���rA{,��%{��4&;O�g��|�����0U+X�b���]&/RDa��L�!o��d�a�e�b�9�*�����p��H�����%�_�V�Rf��L�����BW�<��R���+�bE����:��gQ�i��@»�_҂� ���PUA�d]RU�5�6P,'�>�]�)��h���cWE���Gz�B�J����
�i��:?�%N����"��3����8��Sy��u��~���1��~�t�e/�:����	!�)�h�:𾶎�W݆Jٸ���(N���v��x�\�w�_^��vQJ�1J�S��X�yT}_)BC��ӥ�D�^s��������b4��7�_c�fT�/���~A��K�������B���� h0��ȗ�h��~K�\�����H��o���V��(�27f���z�9�3�3�O��)8w _��5[r���(Q�s��+?�^��)�}��Y����'f(��.b#%>�oiH���7M�+$����	� }�A^WE��^�۴�����V�B	�M<I�l�z1g�j$�v\���h�z�9�2BŌN|�S� ��g�}5�K��_1qu��E�rKm>f=��]����0>��&"�+��.�]`��d���eٵ�{��/}�Xۣ�n���5�K-�Wt;�t�pN�f:|VI�.��p��u���]�F���2>o(!�#�䊵���k`1�x`݃5<-�z3f��*�F"5B���m#U<�"�b�=�]�,�K}����8�_��s��@�:($Gi Hց0(dlH���'Ϥ]�8e����Z���F����Fy���}f�U6���9خ㷨�a?�'	��m<;�B�\z�KK�"i�^��xuor�,��ܛ�}Ó�*����K�Cz������-��G�s��b�5���{�1}{
��v���,z�.�ͩ~�ƟEu�kiF"�@=�?�c��s�-_k��{����L���ڡ��
�8M�7��N�H�`sv%(܆|�G�� �{�	��bp6#��tq��'�.��u�3~��@�Cqak�t3}������vK�Q�g���Jm8wڕ��>>�7}�k�_Ldx��FɅb(�h�Q���v˙Z5)܂^+?��+��{ʱ�n_ ڏ)hũ��:��F��ԧDK}Z!J�Gj�r��MI�6.xȔ&&��$�D�ɍ
W`d��l/������:V����Kk��a�S�PT�[��*IR��N��<��E-�N8�	H�������d�V���4D�h�1J��o٧`��M�&�֊��ɘ"�.�ގ�ŧ@�-��,!�]������e�� w�e�.�O��c���pq=��%1�>�\�C���д�ݖR�!�-��,��%y�-�����}Pj�Z�u#i��`f�p��zEy<)�/?����r����g��$�	Wr�^��6E�gP����z�`S�B(
-�P�l���mj?|��`�w=z`C���ǿ����\���O=vØ�1���tM��Hi'BIe����&F���c�3�����	�]��BO;�Ł w.��%q�96�' ���Ԅ�J��Pzc^���s#c�B&DЫ���Q��ao�G�2�Nl��JR���|=���r�:�k�W��������2����n�Xq6�ٶKoU���:���ߡ�I�nKѾ�
S��8��l`���O�6J�R3u��&z4�톃X$��e���z��i��F��k�i�lB �`�B<l?���'��Nᔏ�L�b[�	8{X�$#mM�����Ή)�X37!�[�s֬;F��.� ���MRڨ��U��!�-7}��{�B�2��#})�Nm\���cč��	h(�8����2����"r�̝c�S�ڟf�x���g��3t~��K.a��-d���e��!�EX�	������!w�ҫ�7�zvb�>�W{M�h�t;V��=���Q_`C���}@E{yDz�`K���&NFX���V{�G�֮��g�Ib�Gy��idzg7��^��x^ۺpd׆`GÂ�E}�T�Ts����<�[�`d��l�4��$Nԍ���) VGxy�% #(�����"7�'pѬ	��&n�߂��4�z���Z7U91I c~ܩS�'�� Wy����������ݲ���p�ic@AM[��[Eڸ�W ˢ4�V�
�l3��yG&��)5YX4W�
��|G��B����2a�Q:��]{G|��6i���M�E [�(�k�j�E�r�s��1P�k�@�~��K�+vP�,e�?0�n/�d�+�(�)>7�RV���Ę��j�fkQ޺�־} ��g��!��|Bֽo���m�D`� u�2s��V*�m7^M8�LV��T֠�����ѐ%,��Ѥ:Vp��5�$M�O@��7DV�RI�4lF9��s!M�7��sĦ7������΃����Eã�xj�2��}"�g�*�u&����d�Qʷu6߷ ���(�6��K8�z�!��UX�굊�S� ����q�C���ĩlNo����w`�ID4���ߘ�i�2������v�o���P�v�2����e���e��.n2��&�s?a����9x�Fd�ͯg
��U�(��Œd��ب���e`�M_��e��:
�B�O=��H�����&�{�lǕ@��3�ƭ�E�˄v5�&�"?ĚEU�,�>�Dq�zΘ� 5��Ã����
P��@;����K���'L/�j�����
� .p}�`;Tʛ�ۿ��h�\̹�8娼O�=�Sz� F�I|�C�f2��=ѡ;����ѹ�1;���w�cl|G\Q��� XcR��)s<(�����q�A�p��$��z��gW�'K_�x*��=�Mg4���ޯ�F���-t�vI�`Q-y��Č�-�Wٗ��>�}���ie��LT����ZF�O|���&بM`�; ��J�Z�� a�t'���w����vK���E�'� ?B~W��>[~��e//x̭Wo"�l��d$�������(ecYX����������	Z��W��A�x�Y�,Gk΁�u�-��B���YK?��	�8&�.����/�_]JA��=ڃҐ��39k���LOQ�����/-�=Anv�"� ��B7(��~�an�&�kGQ��N���4�,o��΍H���1��U����v���g]C��3�$W��r��A�3�K5�����L-g��wvwB���j�Ҩ2U�a�so��7�|���]:{݉�5r�ِ��N`�X�̠c!7�=�2�ě�0��H�A&�$|[."X��O���H.9p�D=��r�
4���7荒8}����3�ٽ�KأlOyn����r@�=��B�R��k��Sۈih�cu��Ѹ/�
h�� �&��߆��Ԅ]�NHc�u��u*�^zj���n:����@�fQA�	�ͬt�">��X.d���^�۸�6#�~�9󭄈���}��p�颍�q'�>iq���� �oE{H�.����N+��]|Kq�j5�)���;D�o�'���*�h$�<����QY��*����᫃+�CW	�|�?������YB���X^u⛪��9��6[u��@��ěD����m qˋ�������Z�M��&��o.��ԛd݀�Ж7JX��ǟ8o�9+����i���	U�̆����:�q�A�^/���ڇ�	&>/���^!7"�Ǝ:�ߡ��O�fɀڞKi�ބ�ۘ��ob|���A�U���]����T`��thY�������%~iF�唌KiE��-�ԝE���&��{�	�~��g�]�t�ل����W�����(�%�l�O1�>���EG���l��-0�
e[X|�/��� 9���T��Ӕ����Tie�k�G{$/�E�5�H�����;��y#�t��q<#�������Oqx�z���at�$��Ќ�%�O���*���Pq�4FЈN�8�"��K�9�iDB)�t=�K��)�y����|�ѵ{U��}�N���z"Y���K<?����~r����6�/�*!x/�*MX��O^t���A�=�MTܒdnb��E�*FxK1�3Y`g�C��v]���$�M�'�	*r�Bg�4 %�;��yI�nuM��Gb�G��a���5{~j$�9���^��`@�H}_/#u�=�JF�˜��������c:I�
��&���j#q��O!M��t^vK�1�~I�=��n���������.݉�Ӳ���xn��_��͒{�<�����a'�5SS�c�B�C�����Yv��(���sH2�u��l�#��w��2W��C$ݛ���¶��Q�}����6���("`vb�D�X�l�Ee��Ӽ�\4��u�Tz��<�V���L[I�T.�Q���k�-Ò{�|1%Ms�[F�$Z�Xy��Nɲ�Rl��KL�}Rq�Q�RP��@�R��݅��	_�wv��B/�͠þ�]���<�x��/�p�-�Ϯ���Q����%����o9te\(Ә�6��p_�H�K�\{�9E��f(ש������cE-������u�6���{���8�5e�|x}��#x (��֫>��=��B2�򂇋�y�O�KJ�ߥ4r��{�]�+]p�R섯�Gj�6�2�i��-�
��y/���Ҡ��f��)d9�Q�dB�TB �0 V�26��7r>��G/����]xo����d� ���1�#3n��u$����$���@M�v���{��9�N#�2�,@[����g�G�;��g�墱��f�$M
����86�{)x7��O<���y��X�ܙږUg���f�0b�D�p�Kz(�}ȫ�wM��w�R�.��֌����2d�\�|��8RG�QpP�uN�������pb�%���qOm5O?}��ʇ�1;�s)i���B4�K�u`kJ�69�$�\�v�l0��I��Rí4����k�à��ԛ�����uZ>!��اvi�>I� �����4{��P��Gd�5�K%���f~���qx��ShZ
���[.�z��������Q2o�����%z��z�d_d[�$	�|��.���n�@�^��̭�:��3���p�M�2�+°Оv3�;��c:#���O2j\	p��	S�w���P��'�3��������1x�ݗYp�dX6fР�}��|��.�����뷺�O���;0W������.�\>D%�\�U�0����236��Pg�?o�?|]���V$�aŐeMqv;o�<�~����kt�ƶ�Q�y4��� �1d�+�kAL��tU�/lx�"}���iɼ��5=�V������8,��f@����MԇC�qKԚW��(&������Hv��Y�@�s9�����`ۅF7�K�+-<�O��)4]�_����J���]�Vۦ��s\8���[�VXt���=��	a)�T k�Aյ���
)s��b�JM:����h; ��%�d^%�-���i����Hi�j�U��*2�p(�@�9V[?�Y��6�_t��N_�K����Xq2R���fcy��;��"��2BĬX�k�Q;���/�,=VD6J�� T��\�� <R*d��Ѐt�V4mq�ć���v��:	�
���
Z�^����O��yQ���=��Mc��ي�+����zO����9�fT�x^�P1�"��ܛ�t�0��n�x_rEV)c��@`$Z�����.�:vc;�����&�ĉ��9��뿋NՖBO�h������0�Fh�[��ά��/�Wb��B]f���gg�0WD�����Y^
��-Rim�|X��P�u���z���BS�w��Z5�U_������)�n�~\H�ۦm������10�I �L�e�\X�eip\�EyX���4O,b<[k�_���Q�we]�����J>+>�R�_�����	Y��hl���=��-f\+a�?���V�I�~t:/�L�y9�p�X��ģ��~��ŀ�:����h5I�N�7���<jw���a)SC �G��b	v�F���/�y.osw��� d��n��R�._|v��?j�!� �'�Q�)vE�u몉��\�����Ƭ=�X7�xF�Ov7�B��,S�	���ozB����'�-C����ɏ�3#�,��3v��S�Ã�J��v)���k�Tup��%e4��#�p*���V�V
i�?�Z�6��q�vLr�����ry��MrY�b��O �!6�Z�욅��'[�)T�`��/��A�*��P���Nf&��jʕ͕Jo�ix^�91�U�wVߒ��)Ez�y���:e��`Ug_��rp ��N�"�[���c��~A�'Nֹۻ�} f�f�H�v-@ IS�ZQ����-_���-�{.��M��&���La~���s���hT>��A����.���f����^+/�Ȇ��+�5�e'���::@���ў�[�7�i<�~�(�4s�^�z�y��P�|�z��֍�=�|�̺?�c���C�e��x�fy�iv[us"�?tjb`� [��x�Tk�i�����M�Q���\EP4�ulE��o>��W�~�~0�8�w�eēt0��S���Rv^����U�ա���\qcQ�/r�YZN��V��
��C�|�J`����&��$�A���6���*�Ҍ��5`P����7�}V� �&� 2�TCy�&1����rÆ>��/oo�@}��V�keq�t�Tߩ�S�����Lv��<����y���B����#Nu#wŎö�ĝg�_\���v��E����CyF�L�vz?T����Fc���٫��}^!<oNpm��3�- �p'�b��MZ�l�,n1HCiei�#����H�P����j���?�ǡY>�E{��@���P����ݝ0�X��>�Zc���� ʀ��z�Y��-���`~�6�%�bM���2�dA��}���t"�W��A↗t1�P
���epUs<�(nS�07"�#�ab�!�gW��(�}�Z�z�ņ��Cg�T�� `��XCU�Yf����/���8^
�怪s��.�)��W<���:X:;N�'��>�<���S�����y/V5��mϖ3m�����aA�&�����D7���t��{ͩ��u�"��D#��Zj�x�c~گ�Fb}b �S�Ѥ6�I���݌����(�� G�x8O�a��Ae�b���B��5L��ԜC7�I�!��"�|�c��tyT#�`��6�I��d"���t�@��҈����:P癫-�J�7�B��4��D7NP!3P2j�����Y�!ĮE�_\n��r>� :e���Gv���q�J�M���]�."��������rQ1�v��=g�/Is^�P�d��z�,�50V���lHڿ�\�M��6%������}�ou��5Mr����@� B��f�sx�V�$�v]]��iKeV�@����/`�_�p$���x�����py�(d
ΰ��*�����V�(�|��*c8�Z��n��hYFG�2�)���=�{�xF���J�ثFՌ�LX�T��[w�S:�RJ;ic>������)�LWvn��h�B[�\��v�b�\R~*�S"���cB���	�/�%Fa����hL0
���;���������t���@����B��݋x�9s�6��|�$F	�� '��9&������a�D������X��Zo�A@2�f����;�!��`��%����(,Y�	�Y��:�
ޣM��O�n(ϹL	�&���O͹�͋k�1��p���ګ�z,|IX&hFК�<rL�}o�9�P��u}�5�`ը�e�������/�r
Hl�0	��f�?G������� ���3����S�����$�x�g������K��b��9]�b�DA�Ų�p���-�fm.�n�)RM����_���
'���+u�	
���D`}��4ٓ!�pW\Bâ�A`�[�R�T�`�˵h7S(.�gɉg���P:
b�#��c�]�{��?Zuv�5�6���A+-�+�a�v�8���h��d���з���6ˣ��
L_����
Cb���~�MS*B���!��Bj�K�e�C�@��2�������:'{��f��`���y�eUq���uN���[V���A~�˧�n�1��c���ʝ%��9
B@�:�����ꢑ�U�T��l[~T ɐ���R�)f��^�բ;��o*w<�
�G���h��/ �2�KE~��(,��N�S��8��*gY����)^�D:���~.�N襗�eaB�bI���=�r�W��[���Aq>��-�M�+�eŕ�J�CY���5,��u�G&BT��`U�6%���BT�r���Q*j�u��Y2����o�sT7\�[� J� |��6R�ޘC��9H��FSY�H	�k����{�<�!/����X�G�2�P��
�2i�}F�����*P4������ɐ,S p�*��8�����΄�y[a��Mz1��Zܸ�e!9�,�0����-ؖ�@�n�tS׈]ѿw�Zv�BZu��S��w��� ����g��#9X��YS�1�Ee���s���?��M�T@��~5�lYtD����طQ�TLOD��<*r�(֜�+nuc�׆�Ղ�����^��M� ���=B�0���5���ũ�3%��ܲ���t-���u}Y�䍕� y���#��"����ЏQ��4���&H�q�ls�ۜ�*Ə�Rv|������3�h̙d�I0�Y�C��v�F��J��NsW�ĭ^�a����9v'ݘSt��_	�o��g���^�Ʊ-��]HR�[{�{�ߗ_����#$� `��q�����d`�j:���"��Z��09Z�yG�p.���Ը���0������N���<�`�(�O`�D��6�6�J3�γh�q�Z��x�Q'���b�%�����p�o�h]�S�>ۑ�:)7`A�P�zd��қ���C��%]L���r^�f�/VRn�p@3j�'���:4�z�&'=v)�6��t��]#����J�ܩ4��n���"�o��8���7�u�C��7�_#�yK�k������W� ��zKV�D"k��.z�,����]�����J�62�Da��ϋn����cfF*�E�調[�[��ݭ��|cL�J��������8���-��y-C�Qo���n�}y��%-%��r�)$US;TK�cG)��~_z�����4������w:N���,�:�tghm"�?�cnR8#��L!��ƃ���^��[põٿ��0�m�O��0�������l��M�R-2\�N*�G{�]2��3x�^Z`���-YD��*�\m
O�R�cGe�\KL�x���C�s�H#p��� H�P���a�qp��w��+��L�����X�W���^��Ȫ)~�X��'����Й�[�_�D�d>'\G���Z��1�2�&p�~)��P���h�'����L�&�>\ =E��.ht!^x:T�*�_Չ:A�ZC���ڧ��������ڠ�f��ms:�2�jH5�(~<��ew�+�ۏ*n�K��-"����/��(�����F	��*m���\}��:����q�*�B�bs,+3/Ojv.�F�����̷�[a~�Њ/�G��&���������~��7���)��%K�t�3�y���*�mf/ɫ�_���œIk7d�X#Q=����Wdj�ܜ�ņ�$DY����r�Y-��ɘ���������jd������F�\$��??�R3�=hf�򁛙_�o����V��n�o*E�SMV��z��*|��a�0�Q��"�כ,X����V?��s�>Eݮ�8��%�����Ռ�����C6�"5e��>�5�	FJh�ڷ�	���*�_�+҉�[�I5����[�%i���Bw!��gN�=e3���j�}���Is�r/~�:�:,�Vy��P��pP+as���x6RE��]A{6�ġ�'�E�y���@����S[F5�� �VNO��fH�@��h5�����	+?���,Wt�Q����Ĥ��I-n��9V�*�Wj��=��Uߍ^��rK?�Z-��L�q����_T�����[�X �ͯ������_�;�<0h�r��gA2�"~gN���y������w���H+�X�	0���d"I`MW,�(ydn��.j�ylL�̣h:�U��_��p�&��� ����#���S^������b\Z� j�}2m�N�O1�6ꙹ�3�vJ�N�%dS1�G�������t�FO�Fg�N���;m�gv�#��\9�EO;��
��Q��5������ڑ�	 �����s�HN�s�g���㰥�v��³C�.����x��g��oK��P�z�����������x���������qd�L6� �M^��;�����ō�eV1��@�iG�����T�P���n`�c#C�E�a	��Y�� �o6��?��Wj���$o{�Ljv�8s�{U�̛}�j��_��U�5"����ժ���ޝIM��V �оT��PFBa����鑞��E��������K�"�u!�>��$i�?�k?v�zw��������^��@M�B� ��?/����Eg��B@?=4N�o������%�^k#i"Б3b1�x+��RӖ@��+:��:��!��T�s�ڕ		r8W�E���M���Lg�#��eH�/�M؉�Iyd(=C��.�.l#Z1�l�D���yWp9���`a�ağ֝1v��B�* ~hУ�B��<e)�����ڡ�m��g�~�R��7\5U|U*U|����"�2���eH5�6X���°�ჵ��Ə��t�&'S�˧iHO�U9��ȸ%�9;����Dw
)J��G�f玡0��u���) �4�0�[��ee*N7�̙�(o�\V�h�5��]��3�,�'�x]/4���6�C����{V�`����gMā��U�锤�^!s��HJ��bedL�qOq��2��h��N��Q���@�3�\�� ������.M(@�/��=�1�T��#k�{���|!���?��C`���eFD����&a�5�؉�y|�
�O-�0u�zq�A;�Y�N�)��s[���Ч��0eI:7� �CNg�H���W�nTg��g�=�X��
}�xoݶ�z3���_L��X��
��|C�T�ѬG[0M?]3�}8��X\!�������������,X��A��x8y��z�"#ݼ+���V�n�GK�?C�C��&����*(��q:�����'��	�|�w�0�8�<Ϲkʜ�D�a�"b)�̄��r��w�ᶟK�6*'ؒ�9�Ϸ����t��'�!��E:�����������C��E�����ppKn_jJ'��_��О}����7��k!�!�����0d��DY�j܄�)�_�����I*����D%gk�*E� ��s`��Ķ�]�^Įk�MM��$�[�C�<�}�`�-[劉C(����&xn��PTy�ҵ�~C��ol���4Ն�g�P�n�3f«� ����:���:��ݨ���7�Xϝ���9��|�J.?y�iտgi3{Iո����S��K�HI�����T���<F�S�����I��2%����xS�}w� T��n�P�k�P�4tg��m,QSܵ�S�V 1����n�@$ �ߧ�_��^b`򎍽�g8��>J�d����6�������ޅm�n9,�k�M&���J��VCjj��uJ�ev������bмLu��p�Ś֍kKu�}1"R�!���T����ʷB�,��/��P�tyB}�ƹv{f��kci �jařI�A0�����"���1� [�Rs�Mb���!W���~">s���^X����L@�%�3�y�ň�,p�h�XXg���G��ͻ��"���G��v���k�l��-���6�ݑ�}2��`~�i±%RJC��w*N0��n�t�w�'m�;��Ly�󪀾�qY�[#]뾬3Zrr�k�oͧ��RI�4`����� H���~\�̟�!zN#yb>��~Z�e�E~8>^.o6���ގ�\/�ee���xT��\!�����.�ԄU9ݞ����:�uّ���q�&�j�*b���.qp�[ϝ�6��7d�P
���j�䂸��8@0k$�J�x����3����
�����O,��Cz�!?y�ޝ)b�3�U&��j"r��}y�s���H
�*t�[�y?�лw^�"���M�&�
�B�����f��s6;%�&u3$�0�ݖ�팾����H�1 �����Ʈ��Rr��z/�?�`U���K������:^����|0�Y�<�
�2����z�
Is	ֈ\D�gH��?�ז���֍�B��^)Է�X���W��^�CzQ����X_	�p���xҢ|G3Vj�A�b����" b���F�#�[��885�r�VS�䒀���W�{�l8]�!O�ct�kq"�"L�V��c�p?������s�")�i��<��ko
�ӷNj'���dn�����vT���5�7F�QkK��Q�ԥ -�o�)�"�]�Gb�P�������i&�^p�?�&�ˎ�Y��~���|��1%>�H3 ֓u���y�����qo�~ac�����qɡO@l"���R������#��lR.��'�I��ƹk���$G�L����k�����j�}�����Ε�oˠngX����p6���ӽ�Ĺ��W%R[^8.f�S"�=
�L�E���9򴡺�.J�q8�g��78��� ��.vNUI�ׯ}����I�<J`�W���Fr.w��
 �2�J/�ߓh0U~m-;?5����U��gXQ�N�eA��f��PfO�P�#pJ�K��@_��k���%�Bz�p��4�a� �"⹠�JDq�������8��I3�d�q1�4w�f0g��y��O:��y��`�bVW����V�&��G��'��on���e�Nk� U�����7ƫ��ܟ'��X]�����e0��e�"!v?�v���{?���W�H�O`�{��}���F�Nk�H��'�!��ɔ4X�N��q�^���=�ڊ��ƀJ��k#��Fg��s(���_�NmI-(}B�=(~�X���,���Y��W�K��Ƀ�FC�h��Hx m8� ^����L�f�����r� ��r.��LK83W��l~O@X�ʣ��1�Е�#=��.��)�?_����f���kef.�t�8��B�j��FkSv�jjY��l�K�|���������2�B��1|t�先_��xo�b��\��ɡ�u�]>HC�Q��U�u��,�n�B���j��2,�#/����?W�ok�������`o��,\0�O�r����6r�Wq*o�]R=������Ɍ+��k3�����
�x��}8�:�
���)�X�P�[��J>�V���5H�
i%tn���f�>zl-��)~f��'�Ә��2Q��N"T��Ú�&�<��HN��@;�/�J��ճl��?찈'�}m}ol�,���x��,{1��cW�NaC�;r�f�0�$���	��*㑐0�n$X S��v{�JZ�q����e�h{���Ð��tUyR�f@���EC�r��D
/F"�8ο=�����S���O[u[7�C&�Ȼ��[;^kt�
�,��N�]���c��2m7���{>��R�k����*�h� �(7�g�nN�!I��^;�W��^�d�4(B�:�%�T��X��lM��Xo�dB<^�P��Uݞi��#K���z�>l3�oI�IfE�lP�mNS3�d��e+��/�_C�a�Ӱ:�]�޸3����݀9��]��U�u~��o�͋q�"\I\��z���z��~]���4���=�%�����x=IA�Ak13���ԯ���?�,��^�%�6���KŒ`����<��/����6.��ȿ[S1�B�(�k�uL%�g�H���66&eZ���Q^?/
! ��]9�b.[XkQu����K��&�������1^e+P�H�+��Մ�)2	&:_����������;���NA±�M�A�M�?FB�<�+�.�ׂ��B��6+mM���%������8�9�&���y�rl���w5S�{^���ݤq��7��C����!A�����"�D׿Vrv�O�i
2�#�����J���=�"B� ���D��<o�g������j��t�)�Ҿ�?��Ҕ�+r*/t�ԇm�o;G��g���N��iʋ��¸�6sХ�1l��Z���J��o�ud)��p�c!��31�����r���tԀ*�G�V�m~>�{y���L�>�d�2�H�ڑ��2㛹P���!���� ���և8�G:؈�l��
� [�/�ZQ$�u����p�5�.�z��p�DWл�At�:�:���g�U�f$b���y4����~�T} �(	mYSחN�o^���t��g>�Z��ӕ��L+o�{�gi�`�!̚��N��7�Z��C[��ڡGD�Y�\���y��"�8ң��I��_H��zӾ�My�$-���y�%l�g��b�W{��U9�H��vNf#�)������u�p�0� X.��f.����G!�n�;k����𬖩�0z�;��"U��O#�W�����`Ɖm�i�b I_��q&'y"���E�Q�g��Z'U�F��㌬c��*u󤰽 ��o������M{-o�B�5��wl���x���$n[�4�p �]�� ,��Kj�+q�V�:�S���jb���
h���ܸ�0�`�QC�X��f=Fɂ�C���콴�P&�8��o�aN%��'}�=�nsm������3����X�6�[*���$�}o����W�S�~���vm7B��	��H��t��ꖅ�Ad�燳���G�}֩��Ex*?,�
�Ю�z�ŷn�NpQ�䂵�U��즽y)V�i	�	��^_t�!Q'6���;�Դ���?����I��J���k��������Zc㬠�`s��]u,��oՙw|Z���b���X`�$%bw
�)+����%\�"gShzb�5��AR��N4����[�|�|��4���97�1iVn�s��;ѵ�PpVsؖh{A�Q�^^i���u㞞���Ibf�Y�p�ς�a2tZV6�uv�%��m��I	���5��������{��y�4��kM��:f5d�5�4�
z�V�2�����n���7�k�5����me���f�y�wㇻA�k����#�D�?�)��|�S�I8��z&��I7��+L�(E[%��OW����d�ߛ`8�����k��������(J�e (m$<j�`��?�����Lq�S/��+�`�=[z˛��Bћ�{���_ۅ 3F��e�&V�3ҫvx�"O4��7�:�Ө�ܳ�fL�G�.��b��շb��bp�>@��̓�ak>c�-�^��_����喏	���q���,�-�"�㝙C0
<?�몒U������v�~}��d��bV����`).Pf
��A�d��Q�Q�-+��w)/0p�\9&�7qhi����}���6�-�OCK��$�j��d��ߣ���q�S4�lc�!��=�p��H9
�W�,	��r�����%k&���_��NP�\��Qǧ:c���k�]];�s�1 E���:V/R����!>�@��7S�SJ����,�ɝI��B��9`in)��'�]�7�q��iy�V��_�&EP�2��c��a'҃��Q����]�
�p��*�k�H|J7�e�F5/�5t���i� ͪd\�.=/�Z�����C��V�W�d�4��L5+���K�|K��GoݛtD�N`���<%�`�NOR�b*O>����K�L�SO�J��3Ihp\]+�y,TI^�=3B �/�Nx�9'�}`�'�d�?��X_6hO�����F�@4p� !N:�>g�v�UW�gf��ۺ)�K��AWX[�ẹ�e�Xlgi�M��s��W���O��7E:�:��0[)��HH�:)��l��4n�8��;�Zt��1ܰ�`��&B�� =uOVF���;+����u� ��^��	uzΒ������ii"��ĠYN�S�ҿ�bֲ6�o#	��]0���tG<ٙ��:?�����xц���м�IE���FD�5I������.:f!�C#�\�����iV}�OEB
N��v���2j?'�K�D�oy�	Q$(',
g"�
��XĔ�Y�`|%z-zQ+3GF�޶��5�hB��G���z
�s/d��U�q�`��V���/q �y�;$N�\�
���+�҇��U�R�RF�&q�@�3)�k	��4�v_(L�8]�d�F�!%�4���A������ &R�k%v�nL�>{v��UC�M�dk#A߮�h�B��洟��6�rh�G1Rm�f�5��X�3��NK}��[e�-N�ɛ=�Q,[���C�����!�s�^n�b��6�v���]��^4Q�����c�u;��r���
5�0�b8*C�@x�)������dNm4�����zE���t��o��u���[�#n�.I�G"��v.k��x=ix����1�%	�#֋S�M�w̷1j5ߏ[�4�	I��q~V�&k��^��YYC��A���QO�e;��_n�t�(/�88�G�ج��j`��/Ă�]PC=��m�4������OI��ĩ��1ҏyOa�6���;4��a���a�e���H�*����Ȯі�GzR6`�Y��Cʡ��@���zE!}V�
}�/S#}s7��b���NUק�� @B�;��
\I�mX���뱆-Wp�X���9�0"�Ĺ�,�iv�m�U��Ҍ�Sߓ�ui�3Z�sF�<��s���2i�w�1R܂�r�h��<��-`��x����3�g��Yk�x�wzķ�`��ܟ��N��Q?}e�)B⺕?,����lFZ���r��G.��X��ą$���)�OФ.�<>�5QV�sș�Od4��9��jF�o5�N\�jK�]��[=-w"DnԂǯ]_2gv�K��v�r�7���ұhpY��l��>ԯ�|k47l��W5eq_�z���H���:���"��-���Z�91�Q���.����T�,`�����g��y۠c�������tł�/6�ѻ̃u�!��lF�ᅉd:��T��R�S��L�(��Ϙ~c��j��n[޹�3%%���bf�B�1&�ԇ��+g쌱)�b�P���`��Q�{cL��-	Y�*.�!ϭ��<�z�Qb��6	(B�}ݕ8A*��Wj|��끙��S��B��iKD����6�e��+�Y�<��h����%]����~,^^M�����e%�h(#��ݑ�ʩry؇���Z�X���[��s?t��|������.��	q%^m�!�1�k"_1+5W�v�Z���%b�S��"����Dq�~�<om��a��>��Z[^Fn|�*���g���� ������bޔNs%!��r-�W_����)�1b�Ϧ(���[@��xԵ�(ry-�'�c>�JP9n�S?8��A='S}7ss��d��6��g��|+�^��z�ä÷����"b.��7Gw�X'��Hߐ��	��֯m����9MBT<a��&V�o6�X_�zRc �?���|�:QI�D�7>K'�!/�l�`s:sa~���Ű�����@��x.ij@+���� 4'&"�i��k[�)�%�AR̼��f�O�Mk�9�Bl���/���ST#���2E	<헏�|��8��1�5�bH|�#��{�X�p��K�oཞG����Rx��|sTG:�!������*&��U_9z|�u���B��h KqhٲY?���@�����#��ѭ1䀹�l1���-&"��#�lI�#�젛�����	�3U�']��U[p'��4q��l
����ִՆ�TБ� mƛ���~{i���汦�a�X��w�4�����ʈ�4_	��R;U,��\��Ph��I�X4:����i�pI�~���lr\+�pE|���6M�.{tt�`�<���֣=R��Ik�&�H�Qn���\f	����o՟
@<���
�"'�G�
n�l������(�>!���h��a<��&����
�h�g,D2!hC�0���mB�����^%-"�����ֲP1[�Ƌ���������8���#y	���M�Z��ٜ3��c��vO�`����F�3@����F�?̿���G[�����,ۀc|H]Kh�ٜ;r���[w��^&��z� �3e�o]�����g�#�P�%wD��+o1�,����9}�a9��ʀ���1o�����`�B�!)��nA�|�ͳo%��l���
�����1��|�Cb=����4��	�n���;��ޮ�1JR/e[}aM�LSVpnù#nV�6��}�_� ��S)�T�X�+�䠅�}�� ��Wˣz1F��VV]��o���"5�Ǝ
�Ȼ�.��-�NPy��"簜�*c�u�;�����j�(�6mgj�<��<z˸r'�"$���zM�l�h2
�s�!�"��Ƚ��To��,���6�zF�2H�����̙fvD�u����%��-�\��h�/bX4·z��1�7sI^uF�=n��dz��1��~�)�9)�!�x�M@�=��H�Ѩ�i9n��%��d��F=?�{�e?kx"ց7�9EyO�¹o_��EOMZM�p��31af�Zf����)f�cHT�paZnP$Aஇ(��s�iaہA\���@����ۄו@���r��'��Y3&��H�s�q�q�$FgZ��Pp���{���Ŷ�̋ܺ�)nq��
�Hq
�èY�n��&�bd��1�\5.x(H���6��������E�5�����8�QpL��ş�8����N]7�D���w��*�4pg���@1,f\�p�-IHِ��������������~ýXM`��Dk�����k>���F��.OG�Z6��r�C��S����_MY��5y%���P�{m�ܾ�4��7::E�NT�5�0��[#p�#�?F���p���%<[?0-��� z=��R7J�� ����<��0z-Z��,w^�T:�!� �o�@t�?�����!�s���r�X�Z��&R
�����,[r���`)П�:d�B���ģ����А�e��"��0g���eyN#4,S[��X"�,�n�U	�H,]�� ����)�sB;Y���)�h3o����8�43,�s���r��o;��M
�0�t�Aj}>�
w��Ҵ��\��3p����ؾ�c�3���M+)ɀaū--��L��SŔV�dlI~K����L��蓒�m�fWv��o,  ��>u��E��ao�xp�:��֛�nL϶��8���	��X�m�
*��ۑ߄=�f����

�I"�G��ot�"f?P���yM*�&]yR�bK����sM/�!s����cib"ʞW֜�H���R�&&!���j���m�=�ЄWTq��֧և���r����1(�2c������fdY���x��0s�[��b�:�� �=��~��oe�a4�߁�ZmnO�\�-@��ҁ��͍�.�L��<R��S�$�#1�%���q9`}w��ʾ�/�%�L#:B$�
٘IX��Q�`��{��ة�\g�����c�/Ϸߟ ,��ǭpKU��Q_#�)zю+��BJ1�.�������9	�/���8�"6縸F�أ@y�p��OS$�2�lk9YD
[�ft�
"T��0R��=gͰћ:��E�]�i�&���V�t����e�*Q�~6+Q���'g$�y�nY��:�3�O��X<iƟ�3���g"_���Yl[�����*�U�g}��ma{�}�nx��N���e3�Ww�H¹�Ӻ�~����.Q��|�v�����u����4�����@o�I�q�w/�;l�|�ؖ��0 ���9|�\�9�8���������Vj��#H00���2�#��N�`<�<�B��=0k�=2�RӶ6N��|�"���ȃ\�=༃4�$��vణB�v�2��m���6�x���zs4`���cm�[���T�L���0�g_ATuϽ�/pf��^���S�u����i\�ĳ�`�����9�p%u21Ib�.d5�����9��3��c6��E�vYw�c�I"Lb)�&�1����*�����PtY�*�����+4���c�c���X��3�Y�`���'.U��J!��?ks����$��4$�rYŝ��y�����^��{�`Ey��,�u�@���/m�h��C[��5���b:��`UMߤ�Ls��S����VG~�k �Qr��+�uQ��#��y̔Z��!�v��RN�=��A�$���η���f!y���=o��n����`����)�C�xaQWF�W�m�rvm��ӳM���C�YZl�64�-�Uw�NR�u��P``z=�ݥ^.s.UUD/¨�vТy�Sk8w��W��6ˣQ���t`@y��>�Yk}�p%��o8\��ǈ�wQ��C`�,��D�7V֕G�����	#_�`WH��ƺ�S�Ձ���n���o~��"���9OFi4�h�����n�h$W�>qё��7���Ē �0��uYO~|޲���[wl�;
��˩E���^����!5&>�ŷA�ތ��Bd����k��ٷ��&7����Sg,������	G�w*����0�8��g� >�&�p����0�]�U^F����'	�ŭ���W��Q���n5 Ug��\�f�⼱:I���F��r��]�wh���E�N�+c)���lt�\:�r�t��M{�LD���I�?�8s�!L�'#v9��\���;;���=��`qXZ=sTe^�D�r�il��c2]���'ȓJ6\S�XE3l��c�8��c����0Zv�!e 8��}����R^p%_R��o�~MӈK��?��iS>D����!�d�m������Jr�^7�4s���?:�@��:`pf ��	�K��턀��\�#"k!��{�zb�1.1��;�qY)�t�)ɶrW��;��}LY����56�]$~��7��s�x29�W�1�z5���W�[
b��R�t��ܝ�b4���S�tU�[������%��oA�����?�x咆�$�IdU���+��!���kt�>���.�	����Y93��ͱ�!��_�o�Z� ��s5%C��4 r��U��?��(aq���3���.�Hf�)Uޝ�	�uH$�[�To�Ni�������n��q����gO�l���9[L��k�fF��B�C1n�0��u|��D����w���Z�����t��%&�̡6�� 67���(v�;�\�ŗ|��aol8�����.�mF�U2;�T�}�������\"�%d���'FI\��Ҏ�����G���!���y�O^l�|�W���k�J���G�HS���ϥ�6�td���M;�� ��W���<��펅<,�C�(�Qހ���	�ʖ���/��7���%��wA�{I%�(�5�G���m>K,�mi{��e�:��y���S����bD���n�!ʋ�Č�-Yg�W@Dک)�F���<JuH�D�xY�Y�Кa�՚~�;��?�.�ŁQ-�j{CG��in��}��D5$���R��*�T<���r-β�3j�I����zv��3��~Z_3��⣟^F?�FH��^G�G���;˼�u/	4�ݱ�����0s�eұ9o�x���E8�S/(B9�KW�r8+��)�Ja��MsF�l�ĺ�Ft�+Ef�+Y�]�;W����f0�E�%�W��g����:����p���[6��꩒�����/�-8���T^����:C�o�Nq��~ɐ���0ȑiT�D3�@O���=�1��&W
\G<ͷC��T!�]f*ޯD>�����j��P�cK*6&F*�@A��-�܌�Gd��KSM[&ڿ���#�\(h�̀緧F���B3\�����ɖ�����,Ƶ�'7�Jl�ڳ| !�_Gr����v���j�[�Ӊk�?a�m�}�|�Uk�I�}���q9�"� �
4�H��m*��`U��'ۣ�O��)�L�����dB�+�u7�L,A��/��J2vK�����W���z��awJ�F��L׭a� w��[�G���Zi(���q�4�0$�gѹ)��hX1��d��vK\1��s��Z�^h���FYW���dv�7��=��in+x	G�Ee���2�S�����u�)әo扑Y�w�=�wye��{�Z�����jy�#�5��j�n�U\����|s�A�#u"��? �����@G7�#���#���M���%�`t�8@��y�m��:���N�C��+��~ �񲤛,Swx�0s�4T�"V��z�de���~5���[�T���7^�֟$��^� �[˰\�6����ۼJYVF��.a�s�n��*�|nM���)��e��\�?�����5쇮	��3Jn�`Ƌo<��b#:�/�B���m��|!/�����z�̔ւ���\!j��F-XԮK�|-�G���}���]e��8�g�k^�|���4�o��i<�>4�f���,�XK2�R�-tP7(��At���$��Ñ�P���9�v���BG��8�ʛ�k$(����7����˗.��o�	4�4��/�r���W.[��g�,Ik�B42v�hۆ��ىpG_���@� ����;��_X��|)g�X�g9M�v)'��I�k>��GYB�8�a��b�)�|1�."����i�B���̲�8�ˎt�o�^S�Q,���L�$�Ā5H�?t+x�����h�T$���#�T���7�$�v����D�y遈�����b|������}[���ؖ����C('��Va���*���@���kh�kMdb*>��:�
)����(G�.�?���.SE%(zL�Df��g�<�������R7`�%+�pf�p�um���]+v��6�I���z2���y9ZF��ึ��.��59(�W�a1qr亪3�$��C�{���̠��L�뿲���{㯏�����K){�A�!��&X9*�:St%���c���l���\���?�֠�}��b}�Q�%��m0��P�s_OZ*�1���@�͏��I"��wg8���z�A�6��/�m-��W��HɵR&(��lp/{-0r�=��0�>�:��1]�(S���Cc�Ff�n]��c�V����e}�M�Њ��j�]���15�1fE��`\�쉇��W���ZpN�:���
�������� N�uz�D����,%���<ÆM��u�D����j/�7��ۼj_R�9��
o4&�����#������)�b�v���3(�:� �g
����&�"��v 
r����ѣtYe�R�}�'��|<�	L,��kh�eИv�M˵z"��D�G�E����N�8��",3�Y�:T�ɮZ���0po�e������&t��k|��Ӹ�~�!Z�h�w���vbBI�𯈓��a}6H�݌����Q�l��pwA���x����Zѐ}m�G�N�|��l@]!y?��[%�rԯw����e�G��B,�#fa�,��B2cڧ�0�0h�e)�u�څ�E��xR�a&	�J�A;b���y��=E��"XK-�(�B\�C=n���3F$:w�ge��M�Wש�K��8�/��D+\4���S����Y�/i���:�B�C ����
݌ ~W�=�U�}�d�V���>���S�@c5g��@t@�fV{����јݘӹ���lX���]H(���u{4=� ��J<��Fe�#�FPx;�@�w	qP�Q�V�1�-��i�u�n��Y�f�c&t�Y�*���79���WK7����B��v�U<$?_���߲IJ� ���h"�^����2�i��s*�&��(��/����$w�zG�uK�R-���+��K�?��5b�}�@�8	m�-_��6>��' 6B�vӅ!������.c~��JSf<w�"�~G1��8B��c���e����'eY�_s�x
R�1��@PH8
���pY�W�:N�'i(:ˌ��:�o ��l׮&j*p3�{J�hy�U%>L�Ě����^s_��l٪��V6�Ќ��ȗ�������D�^Ҽ��6�D5 �P�)cc~ p;�QF����:�I	�x~�𸇼G�?�����ѐ
ވ���<q;��F�g�}R�{��>�0�^��/�)�m�~�U.O�t�����%f��<F�$�5#3Pd�G�]�~i�W@}-�c�c#�kL���L_�N�t9юL>��-�o1�7b�a��L?������t�W���W0�w��Uu��.�[dq�oS�'7 M�I��k^e��Χ8[hdzmv�5�}ʚ��%ͮN8�1���*��2x����G���c�=qo|�¼װ���e�&��B�S_�ŧzw�(n��2�bG����Dd�����S��>�lg3ͼe�]G�a´��o<ρ���>�>�!P)nP+���1d�֪6�`�-�I\���aEE��yX�����7Pv�cHiz�t:4�d�m�R�J��(w�Q��B-1��:F�0�t�e�I զ�B��[Z!�a��A�[��f>�+&���!�!���9������w%Z-�w��J��>�d"��ԛ�>�4.���f}C�ĸ��D�r���	$(�>�x�i�W�f��I��G���lM@�tӭ�6�dZ����D����QW�ǌ�3J����OFd�^���h�ʧPpYD@���Ue�� �F쩲ep]�vY|�`T}]R\'�h�VX���+���j�lN����&��������E�M�.��Z_IR�nT;�6{�ڀ�� _n?�ЫfiY�'
c�q�<���9���m�u����fy �=?/�׭�ZttKU�P�R�)5(���l�ȇ��+
�|���QE�I>���R��2��H�\�{^�7��*��� ��#u�]B��PW��jZ��� �S�	Cd[��m�XڪJ)������C�����ncr�y�V���ȴG���v������
?� ��Z����N�W����^��wG��*J����/C -?��d�B���쎕,g'�ˌ��φ����Z�5m�-NV /�g���ZƳ�Œ��2��t2Äԍ��b�]��F�"��jѓ�4���e�&�2xq]^����5����z9��@
��7[,�\%D��*�8H�}%
�W0�-5�͝�f�FGgEq���� a۩� |M�	IΞ쟇|wD�EZ�-'ASB��[�Ƽӓ�f���{�Y�pK�>�R�3C�Z�<݂�R�2{o>o !T%�ı�@���aq��Y������~z/�M$�����CZF�����l�G�lɃ��[��H�s�z��2����11g-	>)�n����ƛҺn<m]tV�S��R���n/,kq�����w*�Ć/O�0'�������$�o��𔫮�G�T�.(�p��X�Ǎ�1T3Q_D�Q0���g�����#�/"1�$#�K���$��v����I��W��;�4�S��^^p��Vl3L�krM�И������pr��S�A��dj@'��D����c)f��؃̊�=�W ���]��Ԓ�ӆ�#_jG6]�`���D�!�1��UL�/Ҁ���Ϩ�s�R�$�-��Z���iy�����z:�~�<z�Ӏh!�@^O��?T\e�<�ܾ��͘g�{W`&;<�#}��H�k��4}����iW;}iQ?g�+�6=O��~	Uɉ�p�zh0�V�H��Է��6+���x�^2������{J�Ғ ��Ԭs6��bĝ����#}�+~���*�95|�0�3�딮���<��Ww<|�AÄ?G*���y�Щx� �����6��I������$��?�w@�%:������SK>jG�G�v8=~�r3l�� ��1�:E}�z)F�[8]��X���)͞�7�i�c}�fNї��H����GT�Qf��J;����f��	}��ǖ+����8���(��W���zE{ �_�l�r���é�yT%��^�*����wb��C����;�}�"2b�mO�`¿�\OpM.D��z�Eo��5E�yD�:�tDZw��@����w�'�GӅ:��Z@�k�RvH!v�'nowV�1������ �X���J6��Zg���R�L�;d�G'\m���,���CU��̳j��<,����uM���"��G}����V�f��d�?����Kd#�8���8?�P5Xg�֙+�߹��-}�� �}���sþ��W����Vo����rR���4�h����R!���GG��l:f�v#�B`��H'��	?���N�Ҭ�Dna�V�3�d�~i3��5���z���D�������38@T�^"�82��MX�Rа�7> �H��E�kd�^���.?�ę,�B[ p`�V6�~����"Qک^�z��W�]z��������U��,�^";��SBIY�����W�%XM(������,xh�k%QZ�.s��Ըj+�߿�8��K����mr񭯁]`�@w��XP|;w��kz�����cO����i�ׇ��)>2@N��۷/įR+F�����T$���f�[z �Ҡ��܄{6i)~	�&�G̬p��(7 ��,z�-\�!3�:��n�	+R�H4Dc���|��ڐ�������p,Q����=Wف3;�Ҥ&:�gU���۹�J�}|X�\���T�A����2��J,K`ktq�/��W�@�W)�KwƵ�Xy�°�+�pxą��o^n� c��n����:H��*�K{��y���(��,S^��H����;��٭:�����I7�ܷBs��/f����iC�/q ����� 3��/%�#j.�� ��C�X� \�9Jw0L2?U�"��f�MO�~��NtƷ72�Lq�h�0%=�ǩ��J*G����V�\ͧP�L����԰��˲�hz���8&��]���-(h����G�x��g�8���!5� ��Y��VL�W�f�)���P/t�;��b(��d����ʘST�o4l����c�%Ӎzļ�t��=�L��n�X>.���haٻiѧ��o����@;�0Ü�;�p��KPVPH����%�ely��ѳ`;ȥ�����M�!�=o'�W���x�+������V(�9ˡ$�,Q�'t����e&�S��-� �X�.j7%�I�~F\�3�,<37����"����h�ullw.<��E������a=��|&�2�7�BJ�<3+�.�eȇ�>�p��E!���]LM�0�{��L���״�t�V�F9a�TCN����oqe�e�,K=ݳ��3X��B{o(�3떶<���j�jn��.���mCh]b�\���0�)�_�������t.�wc<�[��%P�$�<}���d��o����ĭ;�hPW-���O�������gGz��Z=}m����4��M�p��*��E�[���_w��f�׶`�<�cp�UߣF����t@qCy"��Z=8]�,�.2;�������喱3�,��٩)�ݡ��4h���և�,6V�΃�Z��%���n]��5�` %Ň�:rD�l2�g��A<`��l0Ѯpr���(��XhC��馠B����'�*��Bkt([1�cc�uc�s�v�pnڲ�(�̹d؂��""�t�c��>X#�J�R�Nh�&aBP��Tjv~k~u�b�J,�^̯�qH�> del��g�M�0�Я����hG�M�ۮ�T�ҙ8���zb�c{_o�s���E&�"8p'� �Tf��F�V��E�c�@?���y4o��d����?�c�XU����5�#�j`�kr6φ>�F���������O���lH�5�a�t��S����IK-6SSUP]�H�wA��얣�����a�H�a܅��j}�X-���iTP�zՂ*����͈�z��a�!�p�d�W\��,�v�!�u���Jź�L��Jΐ�F+�8 pM�L��׵E9Cpm��'�#'�+9�#Bpі5E�/�	�y��/�<�wa
$�39�Iy�$@�xK�^��;1�r�?2}<	�!�S'��ҽ��WC�D��虈[�ިH��w�i�`�~p@����x0;�kOn:�I�%*(P�雷���1b���r��B�<P,!z}�r���(���+Q�I�
��Ͼ��p@X` �hoi�q��m�;XB� ���q~�z�|��[8��t��s�M��j���-���!��9�ŃhÍ)��(l뚘�W�W7ç���`̏	��b=����R�]�gz�1�­Șn�����F���ȆF���#jK��F����(���lco E�q�tS�DnZ���ܮ9�0ڈ�0r������o���9�=��Uڋ3�"�v0^9��0�:������G`LM��}}�z�dM"O�Q����]a��8{��k�c��lý/1�7�=!Ϗ�ڵ��>5�󱲞l}d�*r@"؉���q�y��W9j֭4��+{@JN�B��qۥ������`�nd?�j/����'o[��W��B����������%����T�mL��!�A�}���$R%�.�����{��2\��_��!���
v[���s2 � Q�f���͋kZ=nx#�[U����X*N�q����I��e�J�n�n�t�io9�'����AA b�"�־�!���_AՃBW}K��R[[Δ�f���B��cP���`K} ��#���8��b�Ѥ�BX;ܱᬂ�J��Yb�ձ�1���1�i�-�ϲ������1m��d�=d`�@?�G��{��0������UX�tqx���z�U��.�5q�H�Z���N=�1d��U]�,4��O��`Ei�)�C5��oV�\���Uކ[$��KS� (ސXJ�D��=��s]�fS�4a(R��
Z[$�͟>���5;����b��#:���G���0w������L?�KP���������x�f��uZ�Ƌ�fZ��K!�M%�ڇ�g7o��8c�Vd��fw]�B=-�$ن3m�� �)?3����p������|z�v�!ʜ��t1h��s�����!�E,�U�j9�2��>P��`���i킈}�[[�ԢS��Kw��tk�\��f�ۖN�-���v&J�K��[�ue�-��i��Q�k02�w���;3bZz��<`�����Z�;�޶�c���j�2�x�4�)��*Y�yp��r�,}#�X#B��^�k�p���8	ܯ�W��%r9����YQ�
��]��#��-�W�:��婕
�a�LҠ�S҅fq;�f��J΃���v�
�r0��(�ϘcTd1�r"��q�[�U+��6G��v@�t���(Z�6���M��K���˨�+r����}�7n�>�v\��
�)P�:���a�H�������t��.L���4oA}{�L�#B8ñ�ʣ�ꥀn�ڴ��Q��or���}ș���DL������B�H"k�|��:{�7�]5u�">�&���މRsL�zf�#eQQM�"��,�	)8�WCR���rΉz8y�ō+�`�qz�?�
.��N[�ȃ��,���,�f�����e=E��� ���֘;m�=��d7F�xh��dh_��V�	�rV5�( ����)���?�R�fH���fس�:`׾����!�w̕,)I7�㇫^�"Ęm5edv6�YM��Ai�R���&L�nr{}���R�^g���;/�''��&J�\��[�PNa2���B���U���8:o1D�t#u������<Y�_8Ga^�L��HElL�|�7k�Z�GX��w�7B�o7V���L��Y��l:����v�1�p�'�)S�U{m���g<�*!�
�G�2C�41z�4�)P	��eO��gFSz�l9#��
ɻ2�湆�f���'�=@�!U(�Xy.#�Ȼ�
�zF�ݲ}\����ځ����!R��cʮ�;G{�,�A�P��l���)��D�/���7��iὸ	�����+Ϗ� �����#z~���?����Vr��%��*��m�N+N��K�)��1ͳP��\���f�= �.�OB��#�@�8���^��t�����3Y=q�����QC=d$K�؛b�\�}��ꈺeW�?0{BKF�b$},��	{���%�;?����3Na���sbި9K�Dr6L�#��,?>��=R�ҭ�4Ib���,��4��n[�:/����[ӝ���K6J����O�i�K]��:������͝b���\�6���;����W��!̻�3Cz
)gM�8R#s�T �w�)�K�.k:g��V|�ᅴG����$z��nJ��ɷ ��8�)Ev�� ���u߸s��%6^zI�� Ul�y�B8<�?T#Մ|���:t{`	&��d���oY�d�Z3Ė)�з-QbD�5��[�TzִL'�/DɢD��,��p��\I}��[��um���"�h�Y,�~���mZ�c��{a���^�3�c�V9@�8ז<F��g��P&<�c���x\�f��^R��T���I�eZ������
�T���s˒+H����F/N�j�3Մ]7���B�A	�i�����w���o%��6N�.V4�A��ؠ�1�����N4�����k>C�x!:/y]��d` `G2O߈:�.֮P9O/���f��3�X�����?���i���B��I<��FC��
R|c����vC���7� n�.�:9�Fؓ FL�)ӥ���FF:55}��������s������YO/��ko��ZL*�ڊa&U(^��#Z�⟹�wN4�O BuVJ�<�]�'�m%�w�6�t���Qh+\@�P�e�m�/PRy	�G�`'�mE*��l�]V�ua]sq($��?��T$�����@�z!��r�����֙��y�{�o6��T�y&��o/�#��R�y�[�..ޡ])?��8�3�;E�w����{;̱-3�j��(}���ݣوi��^�T2�	mL��[^_�dF�8U�E�g�͌A�o"�����|M����tPJ}@l�U���7�7���Z๲�!Dڹ#����8�7����K�s�7}���e%�|����*�������@_ ��(T�߃rĄ�`a4<Z�&	~�<\�j�Finڡ�4Q�֙(;5��'����P�zH!�=���TIac�E�Q��0�ї���c�bAGV�����Aۗ|@�5��;�ۧb{)Rˀ&�:ٟ_�ɛk:>�VvW���� w��:��`*�<�K���������cb����F�����^����Qзi!�v>�<!�i�x�pq3M�}۪Y�R��c�i���\miv�c��I"�P����{�d��8�1Z��}�=��
:�?D#�Y:s��v*��$��+�Ra�j����Ps�%2/���73G�i
��5�����/��D �� �ɂ��[�֟&�|��]�%�_nA�@� R`�)W�9)*�q�lG��I�6-�,��S�I�Z��j��Q{�&�`p�o�c���7}>�^ ��򄣮n��]�Ϝ0e�"N�;��&������>Q��� �z��� w�1f1��[��sE����8���NR����0fc9Z�=hf7��}_ۡ0G\ ��>�1߂���< Ǉ�ڝy�V��*�/��@ә��
à���q��0%b_��R�0�U]���0l�l6Sܝ����9ߦ�t� ��A�By�����6[F�mm���
>�	�]�tS��u�f����Eq���+o���2��ԺDgm.q$���t���8�|@a�����±U�ʛ�DX1�=[�D�����k[I������Fi\b�}մ1>�8oL|���M�%3�dS��*F7� 	"#Q���\Nv`[�W�6�˧�\��}Ϣ{v�[�8W�6	�iJ�i��\���Νh�MAHu�[x9V��J����#LD����5�Z%��d�*���E���@n9����Q���Pjk���{ �}����5\5�Ӗ�t%\2�,����.70�oY�ف�l�v�����;�3����0��9�8o��
/�-@����;k7����#�N8Z�U�m������Aq��\u���S��l��>u;�|��C �K9��r�L��	���D�x$�/��IhB�����`��}�#��o{���
��嬠Y��n��ӕz�쁖�+[��R>V�a�c�7��C�l/���+z��K*���G���mdR������1Cμ}h�1է���V6�=Z���|\��oru��� �8��z��X�o����Ў��Y���7s�9���޽����Tq��9B�W!�Q�5&tU�b�����;OlG� O��Ss d��E��}��f��!]�$�8%�L�N�o%��������ɋ�&q�z��3;�L!�x�;u2�^0�^M�R��4sw84w�8�h�;O��I��n�����f^�l�U��5ϓjɂ�pj�K��ь8)���%5��8��W`r���4 Bټ'�@�jY@{}���Xǌ�vJy�+�rz����v�5�4kLS��+n/L�����X'���� 
~���>Qb(l�j�ré���\dfv��jFe��uPآ��r�t"c3c<Aw]J�P�?�30Yک$Mэ���e�A菇ynb��OM�C�W簾\�&c�y�����l 7
�����jO��,L��/(��"v���.�d�+U��R�[�=����K4Wش�n���6�e�%�+�ڏ�c�3.i+�W���\J����u`.Ȁş4���� 
Hx���[v{���{�s��q8��]{\CG�AoA��BU��J��Y�Ν�BˁZ�o"���F�:"Ӛc��7� ��" -o�R�����"K�z����B�qP* M$�2p#jc��(Szk;gɃ�E!�C�״�6}�k3��v�eqE�*/�
�N��1�[;4��]<��a��|JENR �$�1<��2��a/��3�M&�����).b�{�P���07�*������ %�l�ٛ�搏�!s��:�����[�T����F���	ώ����(��n�8�«+9$��؆�AdBD���n����4UL��g���%Ԫ ����Y����KC�X��������Q)?76���]x�1�ņ�(�Gi�3]���f�G��[e>y9Q��z�P��ǵ�j3';iATu�P,;��>��7���Z6�ϠUe�a4l.���ȱ&Ղ��%Jp�Ԓ��OKX���vJ��bWP�I�0�V�����vV�Ta:�6�?��������&BI�\;�AiY�/;e5QF(-{�~�R��wN���c�`��(���;y��+�,͂�㝮�V�K[�oҿkfy���b�
�����#ρL�01rA9��s�(7-��{�d
�_�l������v��:P$��9�p�=���w��y��]�W-"�\zO� ���[�Q�4Ve���e��Tl��#�x���۳Vy8Kxi��}"��B(@��l��6М0k0���x�O
��u*&��!!��@�D�78ƹ�PwVX7�m�	f��E%�7�f�I9kYsyG��oΘ�P-9�{�*���Dc}WN��hB��1E��* 9���	C*��<(.y�gR���f̇�J�@\edޒ4�\r-��;��sn�G�۳�<�0� z�!X8]~n�j���䄘_�}�*iv�0��7��Ry^^,`P|X���|'Ƿ�e4)a���N���Cl(A�)�����Xy.�%���
eɘEG�t��3����Q:$�N:_�Mp���������x'�����xN�umS9o�D��N�J���=r�gc���2^�$uű9ck;�Qf�G�|�����K�c�j��Ѱ���,�^�)������@���~�*?��$��0)�r��o',�2G�H7�(�$uWN9�Y'�]�6��u��;���p�Im��<�i������n�z'���:�`�ߣ�_е�R����
�r|�T�|��W��6N>���FJU&��v0�;1�)���k/�>E��)	���=&�Uu�m~|I1Gip�GO~1���q�5�6����ND*�;Q��o`�i�4+%����-��[��~�:�#�YDiUL��rK�7�7L�y�4���3���K����/aD�!ʌ��]�ֆ9�nK��<8C4��DHA�����g�^l5�e�!u.ǵ��F?;��g1 N�r��rNU�Ǐ�aG��Xޖ�	�#����%��%�A^�:�{��C�Z��!�H��F�,�ǈq�B��N+����n���A�(�����)���jr����}H�+�=�w9�N�=���h�&b�צr]�J������0��5����ʨa6X&dU~�g��Pn����[$� �Je2�A�س��U�f�:��p��#�Ew���T�8�ͬe#�z�y8o�yR\�)�U����-�*d��ƭCn�D9,yR��#z�'N���Չ�ҹ�oi:�u
���1�bi�o^�����g�(��6�b:>�����Pٍ.����hE��?���!�X:�8~hg� �
��əϰ�vc9���3��m"��$k���3E<w/��7�����`�lڎ�.E��W�d�IȕM�q��К���2c1,O���)�,N%���ǥ��|�J��sL������4~�l�2����7�[v�'fpt)���d��+z�HoN�E���M��k�Y��+�Bޥ!`�L�_U���:��H�0�ȗhZ ��qq_����h��#3�Oۍ_�}�2KSל����ᴨ���N��X��s��ե�������>�MEIn�A���p�а�V�9EL{��g�qkL�.��kq�B��)��l[|�%��KZ��h��l�5+���H�s��:	�t�8��O�#uoPd{�c��.�9�i���.;��b�a��$@�����4|���z���V�nWF���y �(=�s]�Yx�P���ֵ�$�U��]6�x��dJ�q�i�.�g�8J��+�B|!��XަU��6�?u��q6|Y^������ro�� ��t$��op��j�QE��R��������q�V���J�3bH��2��퓃9�T�3%{h�q�5��Sp]|np a�ƲA�t�)�^S$���Wsӷ�if�f� �����8�3GggǠ�Rd�f?6x��*�����kP*b��$Q3<�Uo���L�`�����l[*��rru\���	Ea��۰��,�4o7����B~T5�!MQ�����g��1ϋ�-\���0V?��:\���ȳ+x���ߣ�B�P6����ϧ��D|߽6���cb������e�^�$O����&f\&ܗ�5��Fӟdp��ᕜ�T�kդ?��zQ�Fn?�4������`�,U&w�{�<�@���a;��?k��" �K0��b����LC���o����h�&A���[u���Gv�+�[��>k�JZ��3�3��/@�9OueA���G��X�����F�X��_��9@�:Y7=\��PZ:����#���|ˍO�� �&���>k]"�,�
B?U�)!�oTG���Pѭ��o u�G�����\1���Ed��q�r�v��xm��`��cDmG��ٝ��,�EK'dD���t�hZ6�h�1Nfܼ�{�/��������0Ji�������JK�M�s=C��m;��rb�x}��O�ٔ-�nX*�G��������qk���U�3�v�UE�fX���O}|��Y:Pl$M�v�4B���c�ר�9�\�j|q�)_��L#la=1��> ����[��g�*�w����#�%<95�?��-�ln{ڦ0c���;9r�،ٞ]��Zn�&<Ѳ2PQ�g�I�j@��d=!vLiN-;.R��&��7��Y�0�(�fk��+l[�ĩ�g�5l	?�3�ce��g}U�/E�Y����p���Ҩ:᏾��%���pN�Hܗi��F�s �D>&C��7���s�i�ڈ�!�N�},M8�d�n�=�E��٘W�T a���4K�V�ab�o��j��p	
;cơ�>D4D���xv�Rʚ�X�wMw���Np̒{��������j�X���8�0>��׬�nS��,�~QF&4�0��.RǨ������]�2�:Y��L�m*Cޱ7��#��~�_���a��馡�����1�Ĥ�S=��%��$���Ǹ௴����wn�M���vP=o�bn�P�7���������Zx�l] z��ォ��'��� �GD���;�|�=������oK��}\���5�v�{��}<VV,�E��M���0�A�Q�h������g���@����7��B��-��h��>bL9�G��i8O|��m�0����k��4�� �5�n�A�e�����v���:=+���QY�93�C�P�>�E����`�e�ୢ#�|hΛp�4G+���W�L��l�é�e���p����M�p"mo�3�ՄO��,9�k%�b��]!�p!��@�g9��HOr�̙x�gG̋fu��W[�=ȃtQ�3A�dz���4����J{f�uU��������
��}'��-�?��D��8���ٮȌL<Cܼ(�>�=V��n���v�D��?%�Ϝ�	�#�iۈ*7:��O@ǒ�/��T�˧�`�l�qu���Zt1Bo�Hԍ�E�M=j,GK%���K�hB�N�v�-*+�������I�����nt�.'�=�W�L��8����~+ۇ4�?\����g��-�@C5��E�/�C���ۂ�55�0��iCd��P�(��>��7�L���*:D��'s�?���x-f�A�{��P1�#�4[A�UC��j�Ӥ��K*9�T`��0�Ĺ��=J	�����1:D9dAi-#�F����sSa��ˏ��띞���tr�0T�׈>)xa9��/=�
.�xx���+��ݟl~Oȑ�O�c<�2�9F��D�]N��3��+#K�h���`F)�t�j�˃}~9t�#7��b�b���1�}�=�(Z�
�{a���چ 9O�q���n��`0$Q<}�uΥ/�A����ս��!��Y���3�7ިÎ�X��e����;�ŀJr�L?��B�~�E�E�`�r��8S�췮w@k��}tʋC���OV.�L7*�":@�LD�I�0bt�9����ϮϦri}���θ�1��K�W���<m����|�ɾ�����'�F�,�}�$
����y�������O����/k#T
��Ә����7U��u�b�⋹��ž����8�E��D�/g�@G'��	�&s�+��4��+�'�+����������d�7@�O�)�;��ǡ��YH�wڱ���(<"�)�#h�I�:�4��DV�#�Y�]���@i�4��Xh��S��n_��g���3�^;�ޞQ�em�f�n=�d'��晤�>ۋn��&9T�h<�NΘ��V��y".a��VZL��ba�1�e����,v$�c������@�sʭt��C�2mN�Gi�AP~���n���d�:�מ:�}�J�bQi���FĊ�z�ecM�cu��PG�����<�x}$ZJB��1�o�η����P󮷗F��?z����卥F,tK�thaP�	I����%�h��S$���\[j��ȱ�@FL���.��1>@0�{5H5�?J�w�|����xV�N�Ճr�I�Ad��O� �{ZV��9s�1(@���c���0���G��Y�$�Uh��Y'��5�G���`�I�[&q�\p���9���#]J�����9��Ο'�V����&��n%�� ��`3i�c��ǛX����<ԅ弝�xHw�B�e��}%�����6�+��1��Lmp���@��D��(nA��*��qt维-�f�faK/|��6�Ǩ�r�h��r;�6g?��1vmދ�B^�f�/H�79�Q�4��䲰q�z+R�
��>����z�2��n15i��BG%���vj�7���
D��i۵bV
Ob�:�P�'�Sw��3d���Π�������9D(ûN8� >�s#B��T��@|��|*(c�Q�U�	�R e�:�۳F;���8��Q��Z x+�y���+)�,T�Ɍq�L�4�DPzI��\cK�M������:3�����)�R3Oa�	�K�9����������?x�?S�R��g�u�� �XR�h~PGcKFX���g$�T��tO���o@|��I2��5�P멨�K�vv�:2<���e�@�����:��� �t�u{1�Á���nR�6ug7X��e>��|�YN��>H�T����K1�e�V�;u�g���%{;��N����إj�h��#Q����š���k"�����߽�ס�_��N���f�N�W%��g+M!�p:����gs�>E���q|�.�D2��J����>C$Ma0
j^E�.�Rĸ`���ʊw�@�����s$�ȯ��~��A��D�KXQM�j]��A�t�T���r��0�������0٭	"����K�D[��XC;�hUjz���{z�Y���e
�u�!��z&M��{q�2�U���k(���� Q����{1�)��A��u-h�D@�cCz@}��Jǝ�{�]�S�@ 2����V&��LۘG^{n+��z2򑪢n���⪓������!������9��v�f�_ٱ�i�u�q���:dg0L�qw�ʉ�����c������	@�(�w������4x@�tŲ�7m�:ة��j�oNV!��歂D�Hfic�1?9����,�;	��k�q7�����I,�=�FKe��ߡQ�:�q��/�K]�V�OVx��K�:�FS�[��kwq4���FAj�bz7���w>R��.+�k}F�~p�F�S�n��W���s}ܿ�d����"�ұX
d��:��*�gPRh�Sݸ6lkڍNЊ6�aK/s�4��|-®�Pf�U�j�����ٶ �O�/��h��Xf������G�~�,�%�[ʕo�
��>�l\A��.%����ZK�2n���i���e>{���r��� �$���+���3T���tx��+����0�{}�um��8"�$�{C�_�G_������٧r��(�d����_Ww��/�ssa���3!��!�������#�Ƨ��|���:��?[�z�D"�}��u�+��4V�O�B�v0�D:�p�3��3�dq�c��z����	�4M�wвp#l�n��(��S���n��ԭ)@�h;���
��;,� 6�|h�P��I-%D>U=�![ꇬ�8
��(^ e�j��ez�6ª����=�L�Զ �����(��˂�+̆N˓;�ã�~p������D]|�0f}��{�����|�UD�$�A��*R��r{�T�asb��F
~���
a�����R%��N<9�����]�F����Ft�ۜ��tި]�X��+����!H&$���S��+E��fQ�=1�>w�]ډ�y�ϱ����.�U�'�j�OӪ[(�H�Szlj��D�����'����6�2���(bI�n���n|Ea��Ɯ�/��ٕc��Ʌ/m:~U�t�U�fTE�f0�a�|���� ��nET�Yv��)~�Vp�h�`L:� ����5�y�W7a'�P�]����|u�m8��\�f(%��E�`I���r��!@��u��j���~Ĳ.���h�6G�J"U�O	�Ys������f!�{��M��@���M��ʻ��5�.e�d�L��֣��g{��,�f�	t�Pb��[�"Qm
;�*���%�3�>l�����t����m�5&PU��*B�VG\0S�K�����o��x��"��V�t�X2��E
52[��ڏf�Ʈ�D*������Sϗʾ�:ǚ/A�<\�~��Gb����Xd�d�^�j��E$�u㘨�a�Ư��u�Y��s� ڃt�b��WZ�y��`�R��O�a��zj6,�D:���4
R�#I˧"ä`´����"46��HX�\Wl�^����A�9���3�m��jGT�M.�� �������qq�3a:���5�r�,U��U��A��Jl��з(�OF�;��g�N����X��$�8x��E%�U.�rh�LY��č!Y������ ��L�b����������K6:˗��	�}�T`ٛ�����I'>�i���˼�!��O�]q^��u��^�0����LzNZƵ���օ���n,'Sf]���&�y}�2L�0���'�\ l����י��
HX�+v�BL��������s��JWAa�Fhgl��P�h���Ҧ�.�2p�:��v@��[�=�a��Qu�l�FT���ts�`� ��`�8�=�F�����T ~���}�	��
�	��8dH�#�ҥ�3���oE���0h�_y��<ً�
XJ-7T"�W��{碓#�>�;�|џ;�s$��A��J�edM��X
?lv�F}uk����W@"�J���ՏP�<U�^�a���nm�uq�A���V���:T��J�n&�;Bm�j�R뽠yo��u��-8R��X�	Y��8N�	 yN�sBNp�̅��Ieh����1���5�s��k����c�8�2�������k_��D'i�W#�����ps�+�!��$߇
��Єj�N_�nD��D��P!_)]X ��40����-_>�b&�>ld��e
N��\<�Pާ\ F@F؏��C���.o}{�k[�'Nj�c�a��Y%9�n&��bw���	�'�=��&�_VX�s����q�t<��(*���s�Ym�m�P�]����>����K� �^�fρȏFX����uJNz����~#�[�F������;��O[pr���녨R����9��K���C�9e�G�;]��>E(<ad���}O9�a�� r2La��������LP�c����s��Q��7��Q�;ń^���n��f���
I�L��>�i,�4כ��Aу>�?�ʌ����g'�
m/���c~s�&�bIN?�e�q}y���R{�-m�@D�����m��$��zw�V$m2�$�z�=�T�"�%S�>^�&,Jm�h�#��6h��'Ǉm9Vۆ������	s4p�G��7!�5��6��
lS���/c��b��;=�^��x���A	�[3/����_ G-�v牵�k�(��կ�PLh9|�f��2W N�Z)�la��"�W���b��k�A�K�N�ώz0�ذmLr LD&��$�j���q���X"K�L[&�w��*أ�ן�J�@�
#�Ȅ��	��ֆu��0^n�;�e�-ϔ+����{i]c�%�&�����j���$�����
��	���I�9cyY���?�DYy+��fv8���W�D���vLCC΂��O��  XZ��� �{�������SD=�u��.��a��>K%?+F���?5�<˂G/���|�(��t`�7	q����M/�<���;p����47;�R;L��p�'s�Ŀ �H�B<]ܘ0]��Kfb�����;�\^;�fC�&�ޟ�{V:�2�

�Ө����B�7�a!\E���@dP��Xm��C婳�#��ו:�d� �<�g�ڱ^��VDbQ��g��P������� X[:��<��ǔ�S0-.�L���կQxp��K���k! ��)�^���=��|E8�{2]3l��~�
#��QZ zN0|�k��t���:�9>$�f��	;Q�A�D�\T�-�%2Y����M�¼�랈a��5֌V���i��*e(�����OG�#]a���>աM�M8ܧd���-�V�j��Q�;�J�i�Y�̰251�3(���}QIo����o08z�� �����Ԑ�A	���L	B��P(��v�&TC�bœ��V�!\Y��m��;U$r=&��S�cA���+~�_Dٴ����!�Z��Uy߶$�k�V��||U�540����4BU��ꇉR�_[<�6;o,���w�a"��!�5����!~͓�����L�E;�.�G߉Cj?6��Z̅��Kh$�+-�x|�����}U|��J��{��/��O������5z�0FNIT��g6~�ncj#��MB���w2�ueO�/,�~,|�I���B��6̍�F�׼%9}A��/�?��=\���%�����rus����/$�0.�#<>�_T��ʺ���GVI���;��.�G�q� �u|�/�2��V�k�\r���ϢD����2q�>+ǉ�D�㤡u�s�d�ib�\��'0��+���
Ȫm�����T4�n�H���iUц�8� � ��N��l�}�&�2$�|w�Zi�<��C�j;�MC�j��Dc(5���C�^�tA��:Q)?h���c<��X�W�$Ώ��!��=�z9Aώ�+� !{=�$:�}# �����\�x:�8�r Q���Q�BkBX-�$Y͠�b�'�E�Ɏ�&���*+�����?`�����b���D����D�nc-��Z�eJzP5@n�h�(�l.�l�wͨ��0�|o�B�c�pq�r�9�X<97|��\��73��fC������6/!�wĲ�$�
�0�zc�F�p~̓�܎�YW�#��dh�V2���?WٲW����<�r�����*�>�>��{��n}� $��sa��F�-W����s��+�Q['�	���1z c$5�bΰ�`�}���m-���]�i�1�?E6D,�t�m��KJ9��ڴ��rΌX`+�S��[�{T=7����:�B*-���"+�rmsՙʇJth	A^�K���TGiDo.O{1 x����H4�\v5a�ip�g�,l4D[��p���`�k��r�Fc$�m�+]����/_�s�ľC�cBL*O(g���h8jY�[Y�>Z��������6B�8q }n����<����x�5�X�"�*��'ʚ���e5���I�O`_Nn�#z%̧��]4mĞBW[ �顡O�ZG���H�.���������(t憑脄������,�����#�w6��*��KG��~�H��U�K@y�f*ޅ�hb���h��_)�KK��m./엁ݡ�5<�!�BW	�G��Ϋ��]��M��)�H���Y4��> ׃�-�f�T9v� �d�C�9V�1f��i鈉}#s���ܷ�+5��\O�!!7�������-"g�x�������[<�竺܇a&=�o���Z2��,W]J{�-����'%d&`��!�DT_�D��{B�3����
1�#��~c���)��.�9�#S
����d,�	���7h����c
�8_T	�����Vj�ф%�0P>m��V�zM�%�X�]"I�5 �P�`��Ƨ�Y?�.>��8�M�J���^��ع�τѕp��9�J��>6	Bu8��"GPyUЯ�T�l���U:���9� �E��~��ۣV�=�5�|H2'�#[�|8���=%Wb�F ��E��q��r�@�L$(^�D���1��fэe�׃�a�OK;����)��dt��6�0��3Â��b�
�Z���Q]>��c�˟�g�@Ŏ��q<R�$hw�!,3̒ϧwyv�����]�,rBcY�cK��
�CS�g���$�%ǿ�dU�Sn�R���=� ���j��ӕqd<��Q�h�Ku��y�Mo�r�W��)����?����9�x��4j]%�H��2h��hz�+�$w�Ǖ�t���*�M����ۏ/�N�5D^MB���P������JPP^}�i�M)�Qe���鱄��e�F���M��a�s:�S	/'�MQ���$���G���mc���A�����[/�������-A&t#Z�<�eK�N��r��? S�EU����e��e���0m�$�I��Q��k�y��BFKfB�(j5�w�9�H�����5��!�.Nٖ���;�z����. }�`���#*pkmJ��8$������Di+w�����(����ڂR{g/������_���_tA~d�6��Mk�ޏ֒b]����4��bآ�Wj���?���^+Kx���l� �T���4t[S n�/wW�?C¹�g����R��XT�Я)��!D谧���O���#i�7�����<�&�+F�2��t�u&��+>�(�WPĤy����c	�@J,8���{��ޢ�}�8�3pK@u�{S�x;Q*@����E0���c"6ƂƆ���*�X����J�*e;��Y$�������= e�4~կ����~���*�T���H�i��^m>�xԆB��j_7Fz�{�汿	G������-&�l��o\>O��� ��Q6�BW4L<�Q�B���VG7|]�c\V�2�"�\�,p��~ų���E�WƝr谖� ��Ԯ��(���7�oB'�ꚷ�{K㭒j�U���u!�ω�7�Y�GϏ�<?�:�?2��Nbqi/��:��,Rh'�ㇳO����<�萤�m�#���&��!{�w��X�Z�k��6��Tٽp7V�ZV$�R��>l���>�J�1�b¹'�D�m�m����|Ԝ��,�-��A��1~6�=�A�I��6����d5����ή0�H8ƄG��3����&��Kg�а&Y�$mbs��{A|z0�đ�6��M|�!�e���2S�t}��U�V�2�w�b��wX��(1L�8g� ��].�K�Jk
�>U���n�1~�< �:,v�i��=�c��9a��?~���,�B��}'�^~w5X��}6Z�}����$.b1G�/>p��n�łm���L��\���#�$vb���I�E$��ً$�����<x���D���[�N���5Lӏ�?�n�%�Q/�!�6� b^�@uy
m�tN�h���&;0棈�,3ýe�"��/��f�8O]ȿ���_��^�T��5S' ������c(�:��1`(�`ֺ�A<� ����sD�Sĕ-�ԙ�۷� ���@�mr��k괳J������G�{�f��)�X�Qq�%,ׁ��x��ʃ4�c.���ZVܔ(����Y�V��f1��t�N��ʗO�8ɵ%���u�~M'9����7`��g7!���ڄG�-�5�����(B��R� GF��v�<MwO���>�E��sc)�0����]�3�$Z}��ASB����k���L�_l��%O�(��
�X��ePL ��յ��Lt7�M��@ٞ�_�c7�������<"��W�Y*�;*�IF�;�`�ɞb�{T�z��o���qI�]�n*4c��>@�T�R�믡c�ű;Aɶz�\3Tt�(&��c���p3�%kU�)��'ƛ3Z�ݞ��U�{]���x�@)k,�:ћb�׍]�m�"�g�͗C�6��27W�jJ%i��9ZR�4��ARh�%���d��n�_^s��*�[���4��wt�nK�cȻv�q;�B>L�T�t��2�[�?!��D#�ýsԫR�gr���f*x# ���=��]�=�e���Q�'Of�����e�t��q��=f��U�3Uz�5x/���:(N���[o�`��;L�ϭ�Y�ߞY�\b��!s
 0>h���&|8�n�$�:�.u�(Z��$�q�Ao�+�/(�z��������!�j߶�^(W�fP�_A׾��iͶH���n�����J~h�(���)0[	�h��ti���6�h�ȕk;���$O�����o��l�y���bWm8P��!��]Û��s�;?b��i���r�٨��Kڲt�k���] �$�b~3�#r}�h�U=���������.A�߳�����ܝ*���`��J��V�s��=�1�S��fO�[��c�He�=.V~p��k[ڲ/�.�3eu�p�O����fN��4�{��(�z�S*�x��V��咮KI�K�(/c�A�O��K���}�5pS��ڧq�7=�g&�/ �p�&m�r~r��	��y�Ӵ=Kc�7&���$���g�'�\Uh~·�yv�5�We0JB���0o]F��yo~��^ E��T�KP�%��^p����P�o��T�`�;�/8��B�rt�٣ۉ̀�����%��aZ+!�A����K�pRzi�0�E�\}L+Y����j��Ⱥ�R�wP��K7q���V�����5�k`Y���ܹxDmG����b�A���\&�(i� ��K�=�ӻ�����3�����$�Ŋ\m�;(��7��}P����z��"�\
���l&� ([��G�k����т�W�yB�ݣ��P�"��H�VEwq�E�f~�o,i�&�'��5v\���rյf�%���8<�vw�Z�OϢ��ݹ�b2Y7��`Pɟ���v�{��K�W�2��&�\��o�)r����'p��_��K�j5'#+�LV�q���F���M�pO�D7 ����k��\W�[�:S�����H%|���+�\�F�������=c�l-z��?��Ï�6&�ˬ]}����[�o,��`�D��َ�~�M��=B���tF�`Fg�AsD�!h�E{��`�~�Fy)ٹۣ9o�z�o�p���2S��-�x��|�"tm��� �G�	p��-��)v�r���_�I*6�@�	��ͼ �� j8�
vj8
���EI�+���?M!"��&$ 1���4K�_���Fl��g�	�T�lǉ�]?��h�Bp2h�Nh0�L��3�q�fe��1�~�D`C�Qht��[�)Ć�_�etB[��;��︸3��|w"�P���ʋKF��#��n����� X��M�-����a	M��)_M��+*�a����
H�����n���b�eG�7��7������Շ<�͙ FD*|�GoG{.D�D���+(���zҞT-Br���!��Gb �p�(ī��Oi�n�p�o�ŀ,~��T;�a\Ü �;a9	���9|ܙ)��xPl���Nb�*uu�=>Xg����1?	Q#��V���D���J������;����[hi��c�<�p�3����Y�Q�,�>�p3�7d���ܪ3U���i�Y�j� �x����<e���)�O�z��yrG~L	<��:�%���k��	�����±׋�=�5/X���+�������~�QJ���$�5(��g�G@l��w~� �iN��P����e��ihI�[�;�TϊG��l�D��p�l���%��s�8ϜK6�qH�q)\�D�ÿ]�s!���J6i4`ů�=�Έ��	���<���:���P3�nX
���%�H��os�m`
�lc�a�?tA��U3Bo��