��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �'�(�٦����6M^� y�N&�hM��\�[ʘS���Z���)/r݇�?*x˯F4<2>����NM��o��E�/Y�tBR�S��j՝�ڕ�!</
]ٷ⟯%��%Dq484)�gL�A�)L��@!h�xr�m����y��4�QM�DG�!S$?oH��;f Vl^7LK��rC�W���r�-d\�!��Ռ딂��?��m�-5�I����'sȘ��q�Gs`����c��� :dk#V9K
�D#�n���s!�W�V�#�>��Z2�c˃�{��d�XS_2��z1�x7�ζh��S������I0���<���o�
��Q��)���aZ&�A����x��Qn��ଔ��*N/-1�<""'��J��n�%��g��8�Z��пg���ڲ�h���
��D���V����x���zj_��DڲM�����s�GJ,��C�C�x;�M@.�xX����M�e�/2ƃ9Zp4����>;?G�S���:srV|ګ��_`M�����i�/1H�c��\�)����B�cc�^�DǪ���!}�!�R@/� �U�k�r%�`�"��$������x�L�}u�B=vyrA��U��W���o��Db\F�IR�G�i1&s��_�kXI&�����R��~ϵ����yPܫ#�R����o�y�Tކ�։�5v~�y�S��8�@���d�Z����777I�A�<0�m2�0�&��
����Hډ�/�:0Щ�ukj���奁_��c����9�����l?�7�0J����h�HV���%tQ-��jqmd]��*�����=��Bh�C��>G1����5'��X2N������xJ�N^��ڵ
 oB7qEzc�*jV���viP-9H�����j�e4� �d��?���O�~�R�y��>w}�zF��;_��mxd���h��ڐ%�r�����}mF/WhLĸ��K�,��Muz�5�b��Ӆ�G�4^ڳ4�bm6��$�J��������Qr�-��H��n۶2�7�e�I,�ަU�ۇ+B{1�"W�q?K�a�×�Нw�|&
"�ͮz�*k#R�����߅���cI�:�?�S"��v��U<�[Z��̈́<�͹f����'���f �چt%�p-��ID�K�)i�M��]�g��>�
�e+7�{�+��M��K�V���E}M'?Ʊޙ�Jl�q،��8P>�sj���J��y٥:'Qw�=%l����Z
 ٗ]�H��Dd V]�_�ދ���u,��7��t.go�� Ӥ��C�Oj�ɦ\���L�we\���|) ��֦Fg��E �$r��6-��L���{�X#/V�$ �Q���*��� �`x/Ǚ ��$�2f#z2^��K/��B*���� ��֢a�!D�v�����O��&�XB�4.V�{@A؏��,\�҆5�Z�iGL]�#���I�y����??����L�	QֲX���:A;�F���zLt�}����z�6��]�p��
��N�-h��3�r�����0��9\������f��4t��or��(�=NOM���|\�p��V,�{G9�����T�3�[��^#�蘑�ֽQ��=��ֈF�Z�D��Z%q��̙ ��.�1��˴�/	�Np��a��?����4��(s=���k?ް�R@�H��5%�Lm^�uA7�%?��k1���4���Г����H��� ��;S�Hn�8&�5���QLB�z���+��e�|���q_ʻV]����*pC��/
/�:s�O�}�'ԝw�UEq9��L��b�|C�%��to�d}����u���!�	H=�A�e� ���6�ɤbw�0p�V|Մv�}�;!��=xf@�4��o�:+h�g7�
ŭp�V�f���f���b2G��|�A��P�>����4����O���b��6�D�ђ2v�K��HJh7��^sV��C#�'�m���
�%����F�?ބ��L(�hU��;�ϧG�a���GAܳ^�)K,�O��C@��t�m��b���jZ\��XF<�a���Lc=}�)HҢO�H8:q�x�pL�P�~�����%�?�+��2����jYr0��)**,ߌa۳2C���+`�6�x�f}r�o���QԹ~��M�L('�G�}b�n:j	%�ФIG8$`�~]���t�8c��8S������"�N��n@Om� �<�4�Ұ��Y�	fL���,�cͅ�s��ɔ!n�a�P�H\����?9�IS�E���G�ir�	�U�.o�Dh: ��QS����:E�uUm�Lr��ǋ��*���<4C
�G�����#f�qd*�w�[M+c��Jb\	�&�� O����D6��#K`��1��V�e�A�߶Z�y��bdS������J|��fa�nOI�b�o>�i�A-���� ��V�9Y���x<�F��>P���'��?\��ke�l�=!~nK�47u@��D�����=�"a-�/��4"4��k�.�)���m�F��d�6�6"E*�RM��Z�)@	�����Ǫ�/ޏq�R&pz(�P9�o8)|���_C�P���W�:к;�ڷ�ӣ	���NY�]Q��;��3�6�ɵn��w����ʏ?9P���������\�#�w{�{3�q�-�$��
����gO���V����G�C~a&&�yg)Y�o%����?l�3=_Qd"��;����)��4E��q���R�/Z~�?m�~�ў��:�����C^�X/�����`	-�t9�c�-����%62"�	��/L��|,E	����<Gi�q���&1}���x�����J�I?�gہ���B���n/���h
��Y�2�Ա�ʡt�1t��Rj4&����`�"���ܥ�Jߥ�Hq��?0�C��|T�ա�"}/l �&�-X�1F�F�ŤD��&7��!�au������_������G��PF�қ
\ ���C3��:6�J@x4�,���׼�eڀ�ꁐ��",���h<:�J�Ş��=+a�WN�t��۴kW�ğCD� ���y3Tݥ���+R�Nʟ6�t���ka��j�v?���Gy�yR�<���f�f��>E���e$�����L�#'YR����Ƀ�q���B�������΁�:� ���&_ ��g	����=�O���)V��K�k��r}Y��&x�� Z�nv�a�%<Z�� g=*T��C�_0���Jn7 K��>���I5�,s� #Wp�a���h?�"N-�C�E`7������
Ф�n���g��0���uVg��hPz��v>?@���f�ei�5<���h��r�p��҅ڦ�C�ɵ��"^�� Wx��#U�E
M���?�R���I����I<"������7S�b�<.�B�87�8��ꭣK$>����Y�6�KW	0�7���/	��Ij~߸����f�F��u�b��+@'1�9�����#��#�}���j�ie� �GmoW��e�u��[�E�=9��o��g&G�+�;� ���2��y��	9�m.^ۂ�+2L���[��׮�^0�B4ܠ���%���t�m�lr5��P�� !��
��B�t��'�����u������ʟ� �"����TCt�%��_�ci�c�.�fRnw�=�bEx$�Z1�X�G�)��Lʘ�!m�/76y�a�8��K��IkT��������z�c�f�^�A�f�"�&�J-�5fH��ױ�d�#��8ky9���C��ʤ�)l��_���N�:��X���Ɯ��Nf��Cm[=�'�ϸ�*��0 ��M��Ŭ%��,�����ʂS�v�ĎƸ��'��h�v���x��CS�uD���
��8����D�����-�z�T;#r���g>-���\5[���|+��D��K46���ᐔ�0Q*�Wv�P��h9�l�J��UJ��?e&���h��b{�|�������`�ugRrT�,I�	���V�����5�j�Zb���.����WEF(�c7)0��P.P�&jOBڐ|��B�J�_�RS�/�gc���?s��vtI�6]���L�͝+�è�@
yA��WO�1�"X��s���߬\I��"G)�p�e=y��u�DC3{�Ǉ̠$�.���GM�14IM�VU2PпJn��[r��`/u�},�Bޢ���t��q�S�p�-���<<�'��Zu`})c��I�j0�{������5���UpΥ�i�+����6b�%'tdQ�%Ɉ� ��[
�Ȫ���nTH�<8pa�*@/�NFߊ�'�� ^�Z��;�#�52#(��00-Q��*𽇗|����ȍ�Q��z�)@y�! �Lc!��*�b�ms^�W���O����G��)��ڶc[j�y	W���py�&N���.���8I|���ݚ����_/�>ȳ�����]����
�9&����g�|!�Q':��q�D.�w�SM㓳�tC�����İ�T&нք�ά�H�	��_n��}~*�B���%�6P��ioe�Ն�2�u�2x")��b@�i&���N�=�P������L�p�mYxx��{C��$	^Z���d�l� �43�jt������ݥ�eK���t�3��2�sd�b�m�}�~R�(�1ӝ����,&�����\������J�p� �<º�X��� ��4�u%�Oj�|	��Y�D���V�?�������BBFo�(h���#V�{tNRH-��4���}��Í��'g�aޠ��fR��$�f�p/`(���r�,/���~��amP�+��j��w���'d�P`�a�������.s��峀��FSBDݰ��.��
�����SQx���ƾ�Q~w�+/�H�T�I`Ď��%E:�r���.=��=Y'� �*����}�+�j�a,�a�����2E�� KŎ�����/��Ҿ�_HXn/�n�����ϳDT�#x��^W�W�X�º�D��fٱ�� ���ҏ�#75����o[���(d@�N�z����Q"��:�\)���~3�Zͻ��JK:3�8�<R�Z,�tv**�����yOV�m�-��� &��p�XDP �:-�p{5�����X�Rpu`q 2���8��l|g� �|���؅��ň��(��t;ߨggI�߃�K/QR��
���61�3.����CT���$&d�v��^��:^�R��2LO�,��I��Sd���b��Q��,� <�H�|߉_鵾�^m+�%�+$O3|�РuL�e.Ҭ�c�DJ�o@'�ifh[��^�t7�xo�65$B��cA쾡8v��T�nztm�7t�k�3ܬ]��~���� n�������NV1��ݴF�"���8*;���0�~ۨ��=���rWQ%8t�G�������ksj��T��h�%n1����c?@n:$�V�[U1vi���c!��{նÊ�%s���Z���20�
�ҽ�G�d����q���E@&r��w��R%��	�3%8F�s�Y�u9�syW�t��9�h�ks�f�)j�t�Rk����18�:�)��m�(�C��P�d�����$$�=��s�T�#j�S��L-�y��+���l7�u�R&�a�@sﳉ�A�;���}E/�n�IJ����f�aŔhYA���^v����������J�1�c^X�_��l(�����8ɼN���` �B����8�Ҟ����L5���M�!M������˄{Jm�|ZubQ6�rZ�u2�����"�LYu�a��cѸ�c~-�<�P8`spy��~����F_;e?����A(�*/������������ѻ	p��Mg"OĠq$a|��:��iu��e�O~/��!aG�х�T��Ĕ7	W���Q�=B	$ ��PkՂȧ���Ǹ�MQ�w�)�C;7*�Ob#�Vhk�]����9�T��-P�"6�M0�WJS��m�r�:��i�Ӄ���a�T^�8���7yC[�^��d�W�X�,d@��Ũx��m��X� ����޿O�����+�e��waK���K�r�/S�q����
��޷Q�U=δ��l�uc}i]���'�1��I澂Ֆz�������j�ĝ�\� �
��o�A��Q��'�ݸoޛI�N+1�'i�|��-[E`ҁ��-���,BY̄���,T��{|�������K�bիtѪjJ�-��Ѵ"�� Z_�о�/�
���]7��c����n[�5Iʿ[�ԣ\�_���E��^O�0>��?�������o���*�\y��-��Y5��4W�~�PBz��T�|x]�"������Q��CxZ��-��C�ު� �e
F�v6�*�I�u%Ӌ�H���'m�H^�a߭�%
>%h6 �LG��`�u�$���]�D������HALsP��"���o��ɕ����Z�������B���q>����`�.ߢ[T��.�n�H/rZ�N�����O.�zG�f��Yo揑�SQ�]ݥ*o���v����j��B�=�\х
��ӷ���٠?q����IuJ��v��R�s��+ijBE��>�U�Mםjr��o�5,�/b3��J�x$GR+�J���,��ooT=��ҕ��r�����N�j'��U��j�p$b����(-z�&�Ɛ�$�d`���*b)ޘ_z�4I~F[�D��ƌN2d{h��-2�g7{��>�f�
���_�O�}��(	`:��Lk,ק;��NJs$���Q��n"�	�`G�|�K'TC�HΣ���}��A��/nd���6��ץs3�9�Xz%Ey��U܎Q�=~�����u��6�Y1����.>���� ��@�ϩ���%#4.���|/
;�fi��P���Wj8�+b�������{Ո-�t��nM��T��b��Z�%ABfs�+�y"Q�aـiP=K$p������^�q�o�?�%��Z"����r�B���2% �5L�Q��Ɏ_'���$[GZ�']���Es���;��WS�����.�1�a/�YȆ(��z)�Ú\]��(�=��Y�:[71��Ɣ��3�k���Eʂ6�1@��MCj%�x�L R%� �u8�L��˨,Ͳd����X�F� [7�T�%8=�}��Oh�Z����	�x���!
��ܬ��34��O���Z�/���`,Ah)� �Sأ(Be�*��Ň:�k0��+�����[�}�$aSN�6u�sʫ����Ez�ר���g�#�4�	�������xb+]��߫�{a���Y��(���8�{�H`8bJ}�#~�}�{zRT@���Y��t��Rj�#V��?B�@��	2��Kl
�*$��ov��%3Ib��D�d��UhP�B�571q� �G�4��&%�FV����7��9	̶v:DX��k�A��A��`�3^�9��F������V�٬�R~��a5�Sqp��$��C᠉y�O��P70�\j~�J�ؓ��>u9���t���UN먼d�L S���N����x�΀�}���|����6�i��}�Ec�Y�y�)��㛀�qj���:��k;	�V�v˵S(����K4�����Mm�$ޜ�@�� �>#���L|��j�ڦq��$l�s��HN>ر����_��3�R�OJ[D��|������R���]ΌP(����lq���nP�����ͧJ��]8��y�_p��,��z9�ں���P����^!7͖�!���G��PzdQ�%��t��ۙ�bR!"B���7p��G~�ҿq3C������X���4Ԗ�A[�z�F�Z�(ä��F��g�fY���:�����☎�_��Ic���[�� `��.��Y��R���~[�*�b�-�"EfUx�j�/ߌ��=�+��A��F�� ��
t�b2��z�)��7�T;�sv���e`�T�X�i��A���t�m�mkZ��!���8��zs���Ka�/4c:dW��hF�fʄ��t��Fe+�a˒`�lzV�c�Db�)��C��3�{+Yw�R��P�c-��z&�y�P?r ��b��V��wH-�z���Š��0A���b1�wI�I��٪Ւ�����K�t����h�a���f+�'4s" ���w}���Ȭ$�&3<�8,K&�"�y�}`�WC�ػ:��E�E�+(��q"�6���ʖ@�]ԄPv资m�����K�/�;����AvGg�y��$�����y�)Z�>��7l�����z���ņe��Z#�_��3/���Q��O}%	r�=�߱7/>�B?sJhm9�{�80fu�f?�� �T��DVUT���%9(�sh�M[�#�"�
@��~�U�ũ����9�o:�w�2}H��<&v��n��*�ڣ��^���6�(���D˖�A�g�@@\�˦����:�x����g�E�X�)��:�s��R~gse�D�W��C���H��O���n�k�U��\^	��L��~��ށ�u�ep�����$�j��>�]0\&f��GoJ7��>M�.��� c.�-���Lrw^ƥ
j�[/�� W	�=��}��2l#�h2I������]�u�V�"�dWT�	7�k�yN�lw*=����DϘZ�Hv���k�D��1�֓�������I���8m#C�*��bp����? ��~j�Y]#4A����p��cqV��� zʛ�����!���P)=�~_aj�;�����'7�e5�z{�h��Z_�S�b������0��f�{[GU��t�Y�O�����C����%Q�*w�e��x$M��4��!��%��zw�V��V�`+��
`.� bc�)�/R��" �M�ڄ��5H�b�4�&�J�Q$|�\���I�s��X�냰Px�l�޲��c�;Xt��M��]Nx~�0����yQ���\K&��͢�`�T�T;�I�d��a�16�xV�50o�x���T���.G�LB��u̳�Tl�VG�v�ʔ�u��>���0�7������[��}j�£h����E.ә�8�J�{�;���j/`}�gߊ�A0�n.����w�.�=N� �/����u�(�CAw���&�Y�O��PB�ϑ��м��}V��$s��5BF�8_���F�%G�H���x4�!�|��4�����<�?[z�*��5�J��AM�+t@�T�/����$B�������q�H�����hX N��ct��]�s��ܕ�=�U�87�*�v�;��[+�H�����"��Mkj���p����Z+�O�A�{�3%�:�A��r��{���M	�8�^�k�p�*�ꏐ����g��c��L��ܞ���p$ݯ�����o�	�y.:v��*[�yO|�0	�fv�����_��ܸ��W�k�.58�-zJe2$c���O/�s��78P2�i$L��o�	l�=?W�=�aK{����˶�U5�Aj�?���[�� c�p&7Q�2qW��'�#������rm7��{�呢ĉ��j��c@|�e�T}�یP��Azq���Qߏ��r���{� �:��d�g$�W�5��Ϝy�@갃H�Hb��^~��ko�>`�2�ce7�\�E.K�E�g���?U�q�EFF�1]��F(]`��?F=��$f�爚�.�U,֍*����e�������{b�7������i���n�	��%K�����ߵ��ߺ��(��� ����B�;h�E����HR����ёg��؝dl��JuQ�1�e�6M��U��#��s ��O�F���B݉��b �ݕNW�qI����Ϗ��7�C��p����O<���+��q��>�邨gn��k���6��N+�}�̑�q���;�@��E}��u�tP�w!��f�� �o=��QӨ^����Lҥu#�Եl����:oj�p��t�]�u��	�C���Q�?�2Q�����.C^�>�mXWOtKhTta{�*���b@��4D�vY7�����1��hy��ʦ1r}k����e�k�s�
!�X���1��O�{+��y�d��m��X�B�˵����Թz�$�/r��၅�l��BF1&/'�0r�7�q�82�#ב��uC���0݂Y?X�n����J�[�/���a�Z2#�����q����:%��d��Q'��Q��bX��۵�Ey�#��,�w�ws×����~Kΰ����$��_K@vO��_+��=$g�SW�fB���	�\��t��2\�}Y���tð;SC~��9��9�>�8|�$���a޻��ShK�/"+�*�F@�%���- �.P��G"K�n���D�<e:���+��Y�u/�HJ��J�Ƣ�1U�ʚy�,�y�ɨQXĠ:d��wk��*��ݑ8�b�b�N��Mj�S*�ŰN=��pu����
�^AXu�i �¯\���[Idi��I[2���g�������-�s��6i���I:k0+�mi�Bo�n��z �F	ַ��T����#Ea�ȩ��rl�(E�u`�.�N��l�>Lf�('�	P�C�g�Z�{�xHo���}�jd�<�S��`7��S�*������dV#t�g�%��ٻE��ƾ���H�.��u�3ae�7y,C��S��t�΂4��XXVH5���n��݀{���)g�:@-~8���?�p�����O��s֨h��� M�"+�����7�M�uH�Xx�E�#1�}M'$`L��?��R�tJ��T2�= ��t5/��ʒ*�XÎ���8L�Z�ܻ��Y��|�$�L[E׹^6�q��q{
h�~���"�FF����rKx[���͘MJ���`݉P���؜?3��Z�Ӫ��o!������3v�5�%��~�\��oFԟ�������z|�1�МJ��Gq>�m��n��X��a���b.S,������(}���
ԍ�01��A�ڣD�KF�	�1 Nt�P��-�9Y�Ò�J��۰��o�/�h�Yv
�Y��4a�`�3�����R ?�Ɗ���H?'?��!R +��G�Z���:�e ���02�v�����ETXIpe7+i����0g<����lq�r%����.8p'����6��ܵB�5�M�Ŭ�D(<���=�^��?w2��C��ar}�ݭ����� !�b��i��OبaUa�T{�&��e��$Pĥ$��Sҧu��lxqe��>�T�㴾�b):yvX+�]qmUt`J��s�W��a����=ֲ���ͺ(4�v^������R�pdd�d���>���\�A�(�eϮF�N��� ��٨M�����v�u�t��,�Y`,+���P�b`{�mvv�7�@��8F��1m�\�=�\�z�.k�!x�(�jp�����86j|��i��3��X����˼ !NlNj��=*�B�T�r�!�\g�e��M[!�w|�e?	�:�$����59�u�Ȫ�t�	f��u
��r1��������:��hwW��U��*톔  (~vB-��4^�Ѳ�5ض�ϊ��a^p��s
�!�M_N��ڈ��7����G�����1��16��
M��uM�N-�\�hΞ&��LtS�7�M�j��"˼���\jV��A�a�-���`�R�5�F�>1��P�Dg<܂�9Prt�LQ���G�C��'(�K>��jS�`7��:��
���AtB��A�U���K�UZ����mx�+{�.R[3��&�,F5���iy�<$!�����I�_s��<����!bR�ȕ����++���ɚk��x4��mM�ˌ�	�j��K�s}�� �h�/Aud�Ҟ���]����C_�1�����MN�z����m�����)z�5�ɠ!�:�>,� 	��&JU�U�T�UCd,�z���Wd3�fz��Z��B��YDJ���4� ���򶠗�덻���cV�L���X����7�O�`K4T�&���ݶ���t�dl3
-�|D��Ժ���񻹖L�>�B9Yw6�ُ�-V����L9�A�eX��o쨖
4@��`+2qԡ�e��@�l�Ǌ��{�k%���g[%�����y���56MY��+�NR-�h��.ʕ���ͦO�s�&�Q����3��D��qt�I{��-(�O�mqΑ~����ⷎ��:Qj��wB����9�'ˠ��J��CP�fX*��e�w'�"$�	k�(����8/;7�6ɪ��e�˼u�%
�e_��
o�gk
6a��qޥє_�D��9N�d�b}���@����t%-Mf�F�`q�#��"Y`�eV��xT?fm�oF�Ǫ!<9(Bk�|]��`l*��R�� dR��2�H��sC2�b��[�����`�����1��<�V!��IޯX#�	Bwi���r�ά��%�] |�U��c&���u�/]F�k��=d|�#o.�_�����vT��K}<¡�F�<�A���?;�$ue̕K��2�34H�����(�����"�
�*׻[�F羻�ւb���A8717E3��gU�
�:$	����S��� "�K�%�忏U�
����%�I�Y�-!��H��#��"��3wQb���_�
��Y��Q)�U���W����翅U�W)�fÕx�`�Ra�S�X-C&�wA����g���ߚ�@�,���D���،3"����]x�$���eQ��X�֔P�S����%=	�����E>�aBȤw��9N:��0|eyǊO͉z�Y��71���Z|���{����Xݹ����Yw]{�a�u�|�5	�$��
a~R����*0��Ҩh�D���e�)H9r�c7���"N���ʯ�ϕ�X�&���9&ۻs���.	���d��|������f��F��P?�e	��0EF���WvLo��p��x̄��	F�L��A��Ω+'�[	�% �|�[�bg0h�&�D�u0<%%e,w���� ��7�N�I�C�)*���=Q��t�1�m0�l�Q���B�%�Լ������~��6��zP�,-�r�Q��L��d��K�۹7����Cz
@�/s\�dO=�Ղ<�RT����p��My
@-��g�L\ң����V��>|~(P@�2@F���z	K��9mz�}��{!�H���f<�;K�B?�m�Q	�ak�n�A�*Пҡo����A����=eưf��+*��T�?48����u�Q��E�Uh Ek΀U�6�v`�����hH���-)���q5Na��ꢞ�v�����&yi����O)Df��1�Z��tY��>���[z]�#xuR#m ��+lDك�W�E�����|͖]�?2�t� ���*��j���)�4�U���2�a��;��Pu�X�2��c����u�=��$D4QG+.�:�ZC�ν��SC^��ىm��2�f� gF�̗�K��ty�}�������uWS�C�ő�� H�Ȝ\�9e;�f���d8���i<�֝VN��?��R�M���q,A\���f_u�$�XD��"cA��P���0%���C�
�o`z�Y�t���u�6���� lV����ue�\�+a�ۙe�^���s
�ێTzR2G:�\jB�a۶u���{(B�:	���ap�àSX]��h.x�؞��`9����y�\O��s8��v "�r��R��8�s7*"�D���$rx��s�5{��K�a�j�/��XZ,3?z�EK�3�a��ҳ�����	E[/��16l�R���u��,�8ם*��qc)Z:�1���h$�����7B1���F\�E��?�v�[|b�*�w�y`;��17�+;�������4����]�Ѽ��.G��ҥa�WFqW�N�ͩ:"Z�ud�(�.ϹH�m~M����F�@&�ŭ]v��57;p��JՆXvE*^�?^��^�q�cz��r��ڝo?c��pg�r�VT5��D��q�y���=S�D��%l�,4����L�A����w�^�W�h����2��f����^	`�9t�?$le�wo�Wr��F��/$����	��f�C���k�(>\�o�B�H8B6]a��������X��%�U�)�-wc��'���#�N"�*v��y�J&�(�=�2���n[AZ�)-���3�k����ŋ��
�n���F��9�װ���he�n��oК
[0�|>q�;�>Y:�4��a"�Ŀ36FB-�~��5����
t5ۈr
��s4�J�������5�:s���e2A׈k���@m��@ڴ�sq�%p��.O_��Hú�d�AQ,f���]0b���$�_��U�`bS�D+��b��������_�9���}%,⚤���;����}Esܤ��Ȉ�zv}C+`�R)K㢌���.j|��^j�F`�q^쟛�X&����.���G�BV��?��?���	�.����u�o������N� ���kZ���.��M�g�R�,/$�vt*y�<u��gz��6V�$�Ͱ�蟵b��А6�Ƨ�� VUɂ�P:DV� ���Q�ϒUZ"^��������g^l?��s>���~���TM�(^��%0��P�	r��Z/��� f~-���D)��؆����`KK�"pr\�����������bUn�
3�Ń-�"�}��I�ɤ��p/r�?��������ll����K%�F�ňW� ��$[����\6gy��!�L�)ϱl��P���m���|���4������Aw~��K��&t�����=�,�y���g�1l���0��UR/s @>[�zzr�?��w��ZߴZ�"�)��
3�o�.7l�Zh�7�vv��8��JN���X�5�!��XȘ3��[��{��#C%q'*�-&�-��U�O�6��=@J��AHk�Vׇ5�85*dD͹����:�S���B�ŋ��q���x&`�d�O��p�Z��K�b^lQ�R�a>w��5(�Aџnemg������@�l9�T��ɝX##�m$����z���Ⱥ�mDC`�
�!�U�]��X��4R.��4L�|C�ܺ�M�D�ž �D B\���Ҷ04����n/�[�I�%NL'X>f���|���˦ݬ�� G��V��Nfj8��˂�3b۩kH s���+��ݫ%Qpʋ��	kca�D8h���Y�Y.���@���ts�%���u�-�a�A��gqAR�BA (@�p��Rl�B�@�@<k�pAG`E���g�{.�[�%"	�f�I�+S0z��t���j^z튾��۵���ԥIJۯCe����1�Yh�$.v��+@)��-߰�EA*��xY^�}Es���"M�;5}QiE܈ŀ��w���Naa�
}�b>^�G]�X����S��]M���$�;]<�٩��y�y�r`��l�H�'WD~����
z��^b��zE�=�2��Y�R�D�:ZVX$?ޙ:�f\�pX��2���.�y,_�bk�:Ub����EY��µ����J�/�(014r���x��;�?B��1�!鎆À�)7,�V�H����;�U��������+�D.�����P�S��rЛ=���aG/Ą`�鵎�Z p�ڕ_
|&��
35n�2�o��Y���J��X�f� ���g;�iiF��((hţp#*=����Ii[T�M����Xv���L���Gs�8ф�LĄ��v�LS�҃�a��{ζ�E~аJ�~�\��Vم�����|��R$c�Pب��GP�)�?eUF�xkU��IM�׭I-fR�G��W񎫒,(	��>Rǂk]ǻ��>wZ]	���c��d&V��r:�_��[7]�Zb��>3� �a��u�vh��X�X��܁K��ǗP�Y:X6�<�DI�u�1jJK��X��a��B�z��MP�B$Q��B�5j�į4��O��X�I�85���hd����6Ѯ%X�r��D�o_�qAxA���4�u��v���x��Mc>~P����Vd�4�F��������k������u�@�� Ýp���(��3>��E���lQ�����e��b�o�AL.)]"bv�����
+���5�~Y�K2	kzRE�H�Pm�U�)*�'D2�}t����~��XH8���]�l1�߸�N������
��1��f���y��z�|{fj�q�ObD����^�aҀ�����%W�啥��֭S
B�p!�rŶѕ����Fii0=�R�Ц2�5�$�ص#�<�MӅl�>�#�`U��4cG�)��6�>�Ǧ/47͈'GGN6t�oĔ�8�F �(�E��̞лLn�T_Ĉ���j�iX��8��?�p��!�Ra]�Q�݉��pp�`�'���[M4���� ��;��4��wJ B�kBLX���>m7�����vO�Ry�\����[QFc)sk��>� �=\纳���mP��O�I�W�@�����T�٭s��F����|����Zp�X��,C�	9mR�ʨò�)~�T"h~+h�j,����Tw������\`cLV?E�݂\Й�+�f�<���7�! ��P�7�a݆&�Rˢ�/=^k�6���'��@��h�&�����¸���RكJ0��iRw��\�+�KR�؁ ��e��j�N{�K��"r�8;L�̈������o�K#��l:89H/��[���N>�6�ؘ�-�:�/z���s�?B��n�V���&<0�W�UX �Ԅ�9��W��R��1S�O���C�\4���)��}`v����������Y�x�@�5j��	:��6��O�4x�#�
˪��ռA;�N+�xjL�)�b���9�eb-�Xjѻ�z�5���o��Z!��"_����Oa���H�5C�������O�%�b)E��9k=��I�tבt� � \��hm6.O����X���_���A���F�!�.Y(�k��b��Is9�����~��1(�a�Z͗�����-LY���7
�~�qCD���j?��h�4�/�mt3�y%w�E��u�Qw�;Ey�pBE�\����	C�����d�!~�@٣D�� �}�э�vXP�w<3����04��3���r(��
^;��e�iu}��|�������CK�R��rz4*���r��>�3�(��?h���l�>(ڹ2�X������K�w8Q��+׎~K���aK�%kO�vΪ��C��s�����,�Q�2�O�����z���S���l`���HOq}�Ti�0�-����3X��wS���8�S��N@��*1��p�>�ق1���r��U���e7����P��2��\=���n�30�0b)���؅W�S�_���ܼ h��^[ł�)�O؄���Dq9�Ѓ��.��.r�����g�ۚ�����=�����˕��ȧ��������������0���u��.���Ҕ��$y}�䪇���?l��'�,'�\
"S�U4���G`���U��o�*3���#i��e��%�gvb����<���e&���_��+��GM�}�
;�o�5�hʍ�c�F!�!ᒍ�I{Y�1����{&�ܤ��^�s��'�)]�-��cI�������z�:[����|z����^�b.�ᕧ&V���R�7��a��`Wz==��Q�ރ���|���l��;w:�![?����_q�S�NUR�`Ow�%��{��2[�%@� p6��q-	�ҖI;�(�v��5.�*���viڠ�Lt^B�����.��@���`���͸����� �y�.�1CNNW������%���S
��15�f����^�n��j��=��w�%ܢ��PIy��?�?�_��bz�;��aCa��>�w�-���~:aC87C�r0>�&�� �=贠�)L�=�uct/?��ǋ� &Nֺ+0�����z����~(������#!���/R����q���3}��&AfkU��'�У,��2��M>���K)ED�7�7��?'o���v�$�.��&��σ�x_�`>]�ۺwp�yz%yvEC�݄diA�eBTH76� �	⥋(^�j�&Z(�},C/�S}�Y�	�6Jx�\���\�cY'ax�ع�����P�d�=&n���
9S�����Fk��ݎ/�q>=�������}��_1rx��(9��H�J���ݦ\2�P�W˾>ԩ�*�� l�*ݬ����-�d�9��EV">z�����)�}��8�_l��@��MN�Q`�'}ѐ����A
1:;\��?��a0*fR���o �a1�!�'[JJt*�v���(Ξ�h���물��_$ �YTWI@9�J�
�CvO�W�E�A�~��֬�i��DzVh ݸ�[B�o��; ���=I<�A׎���h9�K�S��h�_�f���&$$���>��uq.��a��f3�sM����2~�����s6H*{ۯoSzv��- ��h3�k51����e����P��srKm!�o�3��d'��B �NM)딺;��*{��|wlz�1W_�W(�\���i&�I!sܳγd�#A~q^Jx`k��������X����D��+X<zk��}]ͫ�M2cM�<��S�a�1��-u�co��|E�!;�"c'�I��$�K�����8,�9�Wgj���?���;ϣ(���;���d�� 疃�Q�,�̂.5��l��i�Y���"�0�,wv&4�#��!��F&��$�?5�c��^`O���0�\:C�94yn}>�MUSA ���u�#�2Ơ���@��ڠ׼g\ų�G�j<a�&����:��i�K�"�k�y���=�6=A�}V��Z�J�9�Y���b�
`�!1�f�`'-� 蓦�{��fBV�D(��OI�51��D�k9{�G~�-o|���g�k����d*�$�N� B).�9_�:��H�;b�o�?��>�P&2�?jq�,7rXV��ޖ"8*��Z���a�źW&K[�l�	����HHG���n�%�����1�$���w2Ot ��-�HG̫I�:|{��凜O�=�Of�%t�H��[LG �̻?H"�؜+��uOt���vas�@�Z��ԍ�
�~Q󗄺;��R�3h$ct�xjE`����_�҄����6˶l������y;�F����:
	��WNwl��C'=�Ц�<S^����u�p��M���1�:���u�nG%'�. �5f@p�i�43��fP� ,~b>����ɖ��R{_��]^/U�Y���`N	|V��TJ�I60��d��Õ�M�λ9A�/"�~�3��f��T{��D"�� ��j�jb���{���Gն����>s���ǍiG߬\��v�̀u�x�V�R����眀�;ɄKy�",2�[Y� ��2ڼMf��HP����,=�G���&��0�*d�.��o�W���e	W���ّz�M�>��ɏH�]�O�=�tn��^ �2b��paOM%�����Z�: ��\O�K!�V)
L��8pe{%�L�� 25o}�.q��]O�mgᧇӓ���W׼|OD�6ڒ�h��{˟�O�{�Ԩrq=�/�U��2Q����Ay.̗�V1f�9��a�f]	v��[�I��&�-��C5"�\#r*�G�e�Qi�R�l,oE��J�)��щ=�֌�qR���X���� .��
���!�{y���_|&�'��ۣ-�j<)�w�ּ�~�vV$W���Ħc�!���1{����#S�Ә�!�"5ͅ�q�r�g��$$u�����v$W�����˜�6���م.�[�鬬���yo��9��,@�]*[5�*l�����J�Aa>��dA|7k����DZ�.u��m�>r3�Wu�<����4���-��G�J����a��+,[0\��;��xaH���:���}�S���j'q��$DK���y�)� �j�Kv��df�5>b[*���f.��0+��C�l�.�!y ��(e�e���K}xz�O�GF�U4���=���1{�2��lt�m"���?�m��g��Q5���O[��cI$[7R�\f����V]h��"F�\�K �|eL��g%���95R~�*������||Ľl[e�"5
�a�1��M�:�2o�K��c��s=����=-��6?7\r�O����8J����{�.z#P@���G̎��q�^���*^#����0�C&(W��p���^�k��e��jıO��(�Vz�j���v�P�lQ�k,�N��-��Z��]>��J�A�1�{�0Fj2ǖ	�-b���K��]�>U�}V�!O��U3�s�p�sU���(��i�)�!���vJ���gk���E 0�+�G0Z�{~H�u
�Iu���jM�f�]yă�/z�����z�N�B�e��b|�1�Z@5Mٴ�~�r�AhW�`�ob�(�E{�mwk�	/lj�NbɎ�fU�z��K'hMt���U���-�G�3������"��}F&��m�+�+�~I�4TCP��Ҟ��c&ύ\���l3b�n���9)��j^���{u������rҶ�JA��"���"^@�wU�pܼ�hU�,�=����T4����,A�VU�/W<�K����\H׃p� 3����n�����q��~9���T�J���%�0ͅ��l	*�WDf!kq�]��Tk4R���u�?-'�rR��UC�>+�7�N���<�� ��x�2E%�QW�����}qd��Pۗ�$f��_`�������3��� ����
�|�+�+]g��5��`F����x��D�6��vK�

e�
	��T����넄��(�z�7�L�*KBo�WW�4�M{�U�R�_�:�����ơ�F�Ѿ��K�d��#c��CFXw���mUN��n��m�����(8�P�TN���:R貣+C��P�"I�L+���=r����Q�C �V�NC_�)��v���J<�{��������r,��%P�5��wT ��^#݆b\������S>�ԩvOѝDRmڂ�W-T|��v�v�9\b�ђ��Ŝ�R��z|m���x�M$
�&�G�Q�kyD�h�&Yi/[�ޭ��O�:�	��f�I�r0�o>�53�8�8����cjpl������3HE��&I\,�@*��|�=�f�<Hjw/�b�E�I���fĄx�]�]�9^��CM������ q^g����H�sW�gP.��~�����kB%IhF�w��cT����[���p�;�$�X6��L��qѫv����LlM#wd/�_���a�q)R���7`��ݤ��2GѨ�W0e͠�ϚKֈN{8��]�U��݃��s�;GO�h���M��i�{��G�������F�EnZ�npNi���r$t�6�h�/�� ��C��}���+�<�x�'{Djnc����L�	_����.��2���8�/y�k�H﬍��7������x�c�F���֪S�v��1�k�燤���g�1<6�V������|Y/�����E�� 54P��;c�v�
���T���`,��j��~�޻:�Fa���>�н�Lt%��|����
�A>���C\i�M+:���j�>�J��	u��v��{�s�a��jC��d[?E��B�F2Y�6�d��R��m E�8~m��C�7`f���ض%;����9������;�!Of�Y�K�m9
��0���a!��ƻ�v�b7��`$��֧>"7�5^^̿��j1Ԍ`;72�����{i�U2�! MԌ�+-/x6~z�?,ԦF"��>�(��H碳�͈��n'��X��l��ZD��p,M�.�(8�%,�z6iQ9&(�L	K++���!��}��Xx��~{4תv
TD#1k�!=���J0�
j�i��U��ĶI��i�#?e�7���`(a�����4s�=�� � �BhF6߉ *KP<0������Y�RJx�ş��#ș�e�v4W�e��C����Cjkk2ڌ�e[�j��ؠ�����*7�zms�J1�~B�(ʾ�A��Gb�kG,�j�qn9�&+ӗ���4�����v�4���(
�6A�PO�*w��Q0�,��2Ϟ�^�7��3ĵ��6�T�0M�z$�}�|rB��>tM�jMiD���&Xs	O����]�8�2�r��^{s�d�Ug~�������S�n�V��x�]ZOo6�+R@�'�9C���k5��+�����8"�@B�H��f�z�R �oܫ�5���1^/�2� b�-���Z�� w��<���$E5Un*��<�mVsç�#4"9�,N�nOhskYY�H)�^BF	KN��G�`M��JnP��&Uq���1�^��9�(����z�N�K�u�,8�0~;>Ы��7����z�誰��^;�����gV��ȞM@_�ZY�J��eh��G/���:*�7���U>vxK3RԨ�)�{8*XJ9k��`�V8���eĶbT�Hܱ��B �{���ւޞ�Y<���|��V����@�z�n��W� Ϋ���oԿ����oF�N;>��Dr�X�>!�{?ГD8���Kʴ9��������c�̧�c$�4btL�X���tC"���PT��Y-FyA-!�~Hr�
yE�!筲�C� �~��0�i�&[�.+m���6'L|���ƫ�Y��v:a�Uv�>�Nc.t'�� %F:ŖT��!�2=�)S�?���U�*�_���km�GF�G;�x[�ƭ[&}2�L<���X|�]f]���b2��f��E��B��JJ)��et��a�}��T�Q�;T/��O�1��R�R�����B��[n>�L����Sغ��#WN�a�ۧn�^�t�O�f�ʓ�C]��:t�k6�+��0�2P!�k^Q����ܥ���dp���;�ffc��'0e���k�	k��oQ��"�#``)�t
�� ^\5U��xV`�'*):��>�+�^�+���0����g���
�ki��9��:f%È==��&��v�'uq���0�!=)h����n��'{.΂ �����z08����8B�.U�1~��5E�k�gN��è�{z������9����p}�S������<JAn[4w�g$R���ƈ*K�*����Z���0�h�4̔k;�sW��Uƾڎ(%N��Tp��؞�z�0L۳0dyw*_�k��lN�{D:<�&��^��8}k�����
���G���ˡ��0����f�c�.�KӐ�Wo���Ψ,@��C�L�)d��Q��<������Sa3��m���`���q�X.%�����k�����h�bʰkdU�� `�د����o7�t*��:���x�u�ڊ��.�i�n��8Z%ʮz�F�C<詒�(f�g���rD�Z�'�B�I��ȳ��B�βN�`����O);ԋe��ȏ��E68nm��캄�(�!>���n9`y��!�H�6%L�(#�~n�Kx�-+2	W�ҁq!#//�b�G�������N��� f�+7i�����HK���4UK��^Ģ�Z_gE$�=��,�ql�����̽S��M�<D��u�W�asF����Yp���%5A~`��<��.�Ԛ�!b�s#�SH�"��
ĩ�⯎,d��ɥX��'��8H�?c��H�v�l�rS�k�{&�>�!4`�F�Xw�
����Yֈ�8����f��߲x��	5E�N���Rd����\�'t\D��^(-7�"˔?��#5�[W˸��?���	�KZ�׬tg!R^J�@�cԡ��_�N��%�H�����wqD:Y�_�%Em%x���m�jI:����ÒS<�y���TO��`�q��׭F��S����l�E*')"�C�qkix�)[R\��$p[ZS�qpBmF�9�HU��Zfcƍ ��8��6 {��#_PK�=�+q��@q�x�@�H4!�p9<b&�J��zB������4�S�Q�&-8f8�"���~ck>!�x��g��7��

���$>�� +�(�����u�a�j��_�v*/��rpY���sVH���r�9.�GA�H�;3�2d�a11�%�(�AW$�p8��)���4�$�8+�?�� ��񢱅",�OtH[�R?��WY�7��G�yH��34��B�XUd�ñ@�Y���&ƀ1���,�S�`�7��ŷ���u����/�o�&|�J��[2����J��!�G.l)P	ӆܚy�?\�`�[�`�&�c�S��Q��L&��Ԧ%S��ќO�?Il�ɮuS�UQ$�:���������\��Qm��Gոf�y�G�_����>��3���T"�O�{�_	?q�F+��S�M�����ZM]��8�yi�ȴ�^t����U��cѸ�E$�0�	� OmS�Pf��@��I%��*(�mvX�nؚ�\�x������>�A��Z_�KrM�G/��#ũ�M1�m��3lR���K��B�[����ʄ�Q��tݐr���g(�#߄2��X�4�ŽI�j"7׆�C� ���mv��R�#|_x�MbR{"^-�J7�����%��.�	)	�������"�K���"�P��z�R��gYM��
��8��S�&�߻9(�%��~�
2�x��+ 5C���q󽸆�p�8�ޅ��ՁI���A�����R)Z��7j%���g���@���|��g�bq�����7��d� �&	غ��'�_ȁ��5�W	:t�
.m�!���"6&:���X6�GM����82�� �{c��4u�G������j�>K�t����W���"l77@��<��҅��kq��
����\E�Jwyc�:R�r/ֲf룏��5)��6X�堚a*�"��kn�S'��u�2��[#ș !�<�a�WR�u���[�3A��|O/w�p~�����2�}WZ~�P�@X�T�a{J1��%Y/Չ���Q�,u����ɭ��M.�O�6��-P8���nX�x^u|}�� �+��R|T]%�A��!�&Zh�����=R؆W��0	������o�:�ݍh?�K"��ٺUȯ,r�	��_�aP���kT�F�+�).f���2O?0��=vm��{�R��8�1�q69~@rI��8��|ǳ�~wH?�Ml
	��&p��c�W�w_V\�@(�;꼽"C�>�T5��K��$a�e)I[�D�>�i��:��K�e켘J\� �}1g��*?޲6`X�f�sJ1�_ѫQH�[.��G��̘�:�����OpK����T
�Y��i�3�}	x@��*ωF��"���R��%��[�k?��{��9c�E[��萣;nXXrk�܁�/��^$�yK��A����;Br���/\6=��k0��kX1��j3GL Xȷ%i�1Z��˕X����ķTҋ����_���h���������z)"����!�k��.�l)51C��~�!۩3<�wc��+̊�`XT�=Xx�~��}TG���))_�����̩����9 8�=��=�U|iL��7��to�DM^WP6���)�o�5k]�*�9U�/��6�@�o�v�`�]J�6��A}������E��+�m���ڸǱ�|��V@����wT,�����D����³+�D� S��Ӕ@�4��u����֕h\+�*����^~uc��ky��f�}N7���o���K�b�"�H��Ӕ����M<�	l�D�nZ���A�C�	9rc�R�c�;�o�4��8�����q����{���v��v��ū>�VW�n�.iᛌ�t9Ip���`���'�ŭ60ZΠ�@Ü.��3���75�P��
�ڵ��
��iXZ��P��_��L�Ƕр�Uky�u/�1���?Ċ��^0�A���ˈskF��pR{� \uD����
�Π�8��YM��ఌ�z��	�!�������y��%<�};�$a�T7W�	v����ȗ�����!�o��5�f�$����P�tc�P�5`�ө�b,Ѝ�3�7�s�j��e8��M1#������2��sG�2�4��6�ȣ'܂A!�����z���_p=bR�p#�Lp߰RO���Oi�]���%��5h�}���1�!�N���r�{�h����j�9&RŁy�2bs^9l��j�嵜I��w��K�^�)�����V�Gr�Gq� ��L�b<l�@�H�ܫW.N�f��x�,��Sűq�	�M����i�Q����J��g	6����1�f� ��ܑ���������Mt+�P	b�)��)0MQ�c�]�I��8Y�_K�q�q3�7�1v.ɱ�����co����|;G�T5[��JV����dnr�.cӃ)�l��vݲ����hR�j�	<�ϸ�оy ��6Q����R�=:��|!��G�B��Kr_V���le��hF��J����LL����b��֭�H��O�[T���PzX�;��ˋ�"��?b�����J/B�`N�&'�o%���vB��ׂJ����TW��ax���q�T9&�b��&y����&-�C~�oe���9M�{��H��~uq�4uj���ڙ)F�2�Ic+��B�)_�zs��]��7�Kܗ�c9\�E�x:���e$� ���"��)41J�Qsi^��J��6��k�{�)?��m�nN'mM���p�.(�����YW���VT1�!�{s/�R� vza{Rli+���4��y�l�:/8�K
8+����k���ctH��W��g�!��$�����n�S�$;69��p��c%�d��$��bȸ�2���@��Idu|�X��a���h�����zϨ	��U'`�Ҧm��6e�d�U#tw	�fך���@�-��Lf=�7�6�F?nHʑ�I�e�[!�.�V�Jڊu#��i�,W��9�?$��0�#��~��ԭ!��.V`���וs�����@��9��ɹZ2��宅��UiC�. �i/�p�ۊ-0���C�����S���Ϻ�� ��Otv��ہǶi��*��qR�v���Z�M_�I�E���8/nӴ���^h*�HC��P�����&�u�Ҩ+�+�B%%�nMh��s4Ă���B�\dg�1%ퟨ���
�ɻG�!�8.	���yt�Mv�x��e�����Yt@)p����;j=?}]|ؽ��2`g.����?%�����%;P�m��կ�?Re�d>&7Y����^,זq& %sDW~w@{j/ˀ�|C�
ێ��SHv�N��xL�}�T~9�g!`��Ƃ�Q�J�#�\+�*l=f�հq�5Eൻ������k�X�����4sk�gj�XL
��	2�'�S~��U1S55�k

RҠ�@���y2��+ՒYPY�˴4ɱ���4��_��&�q��^`��\����s��D2e-G��(���_j�&�����T��!���6�o�Cl���*U��	H釬.e4�f���'��Q�)IjO�BWА"��*Y|�#�z�g���⸋�b��d̞�궛� S�䊀�41)]��u���^B��%�	a!`dN�������C�ҝfn�fby?
ԽN\�%�` {��BTx��ι
u@�{�xg�� ǈ�鍆&� 6+I经&�-_Lo��::�p�,`���ٍ��eР�[m����@�ʪ93y����w���j����I��:r]�g7���� ��@r�@����*�G�4��ӑx.�*u�{<>��w�4��̝��q����G/f�]N���Vj��{SP8�#�����l~[μ�Omڋ�^��Y�l\��\��2����)]ek�u�g���ʛ�����~�Wi-vX5S[މ��\6VDS�MF΂� 蒀r��&�,�2�sHL߿��ѹ�WƉ�lږ�g ��rW$3�'�i8�I�k���wr��M7:b&Cс�H���s� �᳇ae��������Q*8�~c�o�� �������ֱ4��3�YSl?�5�%{д��ĸC�@��.")n(IpN�p��z`3ay��ؑ��'aL";a"66஄�
	�eޯ�5\ם� #y!I���"囑c���R���qGiW��D� #b�'��C��,b���Z�n:�S���'(��Pc9�^`Gr6N''%�����)oxj�Ů��]��1S���j;7����'ŉN�[���Q���m���$]p�j@9!c�jV����M�v��Z"�P�����_�V"����u��B�2��*x����-�zN eii�1{�oX35H���/��a��{Aι�h3pS@)]#�i��&k�A���iO0(��叡�ֿ���Ă)�#Ɔ�VFY�J����o[�0��x��K���l�I��"ٹ_���#|{�?|꧘j@]��X���qo`[kh2��U�9��:�vlН�!����D�صΐ@Kp��AIF�o`L��$�C���D�M�'��0�y[k�:>�[p6@?���A�;�����+!x��;�w�M���l2��/�h26A���/����xs��p�}B�Dq���nh�ԭ<�"ɫu�i���� P�/9y+3f ���ŷ��>ר�&�xU1�����>�rW�	�'j�v��.M&^�$�x��Xܜ��:���\͇���2\|`S+VF0����+K��ʴ{�g�4@`�i�Y�ͫ:�@���}��)(�/�	�9rp3�W��\��������Z�6Q��V�9.([�0��b˳a�����l���Lw�e&/=��^TT�Xbٌ�O��V�οcfDL�����_L*	_�$Rb%�t�to�ޒ%ϯ��>C�dHFI�j~����J�.�ĵ�R>�+e�qC[�o��
Y�ue�I4T��1�(��k��CĂ^I5<������zQ�2�X��$g���&A�;0�,Â��>�2��Ж���S=��B81�b%仝�0g�x��%�� TŊkȷd��[�
zf��U�9 ��8X�et�L��u����������$�
k����i�'�_���s�����o�6y3��H;���]C��\0o�~��+X�P[d�<�#V���?���]�m��ws�$�Ԭ���&p��eru�"���I�S��ّl�Ž��"Z�^��4:�d�)G~��A��+ ��4KhN)�`�(���5��E�_�.�+)�����y��<p쯟�]��� ���~���l��A(Յ��W�\��5o�oX�/�6�2k$���Ź3|�-9=@n�$�L^�Ph���<�Az$ə7��jt�8�����o���	|�e�Ӥ����Wc*CB�@���\$���X��3����_�SY����4ޞ���A�"�^p������j�����6*�`��J��'�塂md���o�C��}�}�c��*lK�!�G;�?���:��#��O�F|�A��X������K�sU��)�_v�y�oQe�"3�j���oA�7�vGf;i#�$�%��n�1EK�-�]�}
Q�N�;-) -�|�W���"�[,O����NI&se�
!���w(l��M����F��U{x_�:���m���4�i��Ni�(znwsy ���d�>��oڪS�}�8�=FV��8[�u�>:Q���]��	N���~ݺ�ħC�k=�����'u�bw�6�Ĉ>�uw�eDÛ+oy�-
-Z/�W��U�XZN?��Yb��� E:$d@R&�v���\�|�c��s��>���e�N��EEW��M��8��m���~�	g�����5�5b3R�$���W�V2=i&���g�\{�?P��K^�!�۳qn�
>�q�9�0]���ZU�L�M���AC�� Ev�~,Md�8o6 ���#�r�#y�<x��]Jsrl�\�	Q�c�9'������'���Ş�����7�&ȩ�٩��
��Tv�&���ҠPl����!|�1,on���H�ʪN#�d��뗪���Τ�C�<|��Yڰ�Z�E�Z�pG�=��4�`'��Hv9톘5�6��a^��j��[V!��M:V�Gr:��Bn�V�,��D,�hC���k�?W^���G������:)Ѿ61@��b/�\���3P"�:E�ہl�u� �K��k�i�L��V���u҃�h��63����<l��r�����������?�y���ؾ� �-�]�;���/��e��!<m����a	a:�or<���d*/Vo[���]Uz@�3ìKVIF:>Fm�FI����b�2�M��?�Bqk�n���e����h�.�q2?ݿCѢ�8`R}��zp�bC}�D�y�dad�/�!|Z}\�/O�ػa��3^�zv���,[.c&>���9�2`G��@<���n��ҙ������h���=K��eeݡ@AM�.UB�\?��jA/�\�a�8���w)Ō�`J���<�m�d��UY��s�W�F���{\���B��c���;�eR��9����k�T�s/��f�f�G��t���Xv���'��whSt��A��E�=����Â9vE��;����+����E3�|:�d���bN��v���q&������T��R�+�������~,�_d +��+���^� �\��/3⁛�NT�|���E�&���q�cM��@ʂ��U�Q�^�����{�-�η&(���DC ��T&ô�b���"��F��iDGh�EW
M�IN���?+|(���w�`��S��`�(��̇#��Z遖a�[�.��k�k!�����Via7�����;������9*��&F.�w,-IԵ;IYO��Ů�8�s����#�"�j��N$)�sg��)`%���\Pa�i^��|<��TG&��y2l:��Hv��H�OkIVG9��b&�sL���刢{�#�F1�.�0`���@Х�Zi,>�9�������;���4�wNȦp��aŔr��#*�=O�.,[���\��N ߣ@�&�����r(�5���O�j����颕Շ��  �Ȑ���2|���C� ^��pN��28�<��h% �橞`>��/�~O-�znhp�+R��q�uK��s�e��%�5�#¤%�K����b����l%�s~dE�!��6�kM��a 0rYx"	H�O��P�o������T�(�P$�+
�r�w��A�x;»]�u>%�.�,���:^���۳�څf:(%�"RA���bs��� ��'���[��֍Z|��/�]�@VlI���6����d��Z�|��-;�\~�h��
��<��'u<,�q�5�M�5*=�6�5򲘓t�n��q�6��4��Yx$P%.����Hu��D9�dFϳr~��ڢ���䴻�FV���={z#P�8}�Z�� rm��z,E��"R}���C��S�;��x�[��;��2��'>?�3�%�S:�%^�vC �.C<��Qmk��!;�:r�+��	4F�{���㫐����,���6't��Fw �8���-�n�P��,(�Ө�{����	ބ�{�le|l�l^J�\��d�윶M�|Đ2}�&*��L��,H�L��T��|R		5�]<M�T����<9f��~e���6�FU0
Z���8E"���^`f�j�w0��ޤ�Kb�%L�Ŷ�~C�}��@��G3���<�����*����x�U��ݬ��5��jǔ�C���+l��K�z��˻Ǌ���WxIAf�*3u��+HӒO�'q��Ha�
��_�	*�[Wf�{\�*!��
���!&=d�~O���B�C-�<d��A�5�ɐ@��}Xͱ\k'��a�.�Y�����)Г���� a��Y�¡��ϊ;,H7�"Ş�b��gv��͟��15�K�Wd��5B�~�Z7]v_!mo��׺��^��K3��!
ā�����'�7���k��~Bz�@����ο�{�S7rᷩ��۳=�̈4��E:���T-���4�f�tfq
�5�c1+>_�s��2 *�����aE��=tk�@챯�u��,{�ɤ�C'B��=��o3�3�;Ą�B72�ߞf�qu��۝G���f���˪	�@!�BW�z2M�P�]&6��⍴zH�ʈ��ٹm�Fw؛����]��^�"%�ค	\�9g���$lʭ�<t���{��%{֮���MF=M,5�m��ҧ�V��%-	���\�+�.&2'HnwU�Y�s1,��M�U(��q�q�\)�c�D)��-����9�� ��cfj�W�c���'4MUG��=�/��B 0�G��V"�u��K>�R��H2����Ԩ���
�K����;:Ñ�k��l៛,�L�s�̔;�Fn�6�"d��y!�C��� ��離���٣�V���#��@T�S9.��ٳݭ�+i;2��0�f�,�k�0��
p~��U���CY<Rp�8Wb@��Q�����h��`ǹ^[�Xt�=_���+��y�3��s[n��gi��|ٙ��F�44c��,q�_S-H�>r	��SƓ7-�?/FT�(�;��]e�Ҩr�#
1k����b7�.U�۫��/J��8(���.��@��[*���:E�$���\�����+[-�_���p���L�B}���Sy)��f�9}�l����.R�,cbű�+����}�� m�R'�W4��
��&����0s�{� ���ja"Mͱ��H�VU��S�~��Z{�tGT��� ��o���iO�C�
s:l�7�:����[�^�5�۴.\�B�t��8^M�P'/{_��F���������� $:����s��[�A�c��'��%S=�����(�mӂ�bmㇼ�@�]s��kAEbC=��? ����'��\���w���%������,��x�U�j�w��J��/�2�Zi �����A�b>q����v�2�Ɩ�_��'�1U��l��aCU��M��������j2+������B7����\����߅N�p;��'+�w�������!{��rE��tx{��Xr��� E��ֹ�9�c�o���Sy� �[��9�F9��&��(�T�8@iۻ<��cH�zY�^B�29.����Uk,��n݁�Y{4�nyHg���8��/?C�ǘv}��_3�Q7F��a�3<��\u�0ApNj���ΰ+�{�.�F�����1���^�]��C������n�u�u��k%�u��˶Ֆ�l۝ ��X��n04pL�b�ڥ>+,�ު�
��i܉ҟ�TM`��&$�l@�N����[Mh?o����Z���|��w9K����)ɛ>���pf�W��P�~�>��"��ɉ᥿-K��7�HȚ�>��,�ao�4W�
"Oԏ2��Ňom@��n5���/��"-�mʄ��B�wé�(,�:�����,OϪ�=�Ȭ���>T���ϩEwbl谟 �'I��'I�o_Z����� �qC���'%����4G�3�z2N�l��d�������ZLԡR& (����֏^qS��-�����ڻ�^���C�z�}������,���Pe�̏�zc[F�t-�R���9WrѪ�1�#�T8HB��F�XԨ(>dN��m	t�!�1�>�Ā� n��I��/�47/[ ��Ga�X?��*;�@`[�\è��33v����"�qc`@wa�2�\�w���7�9U�tŘ{?�������'7���:Z�JxR�l���3Z�+���!��vW'ţޮ�9������-z-�HC�1�[u�Yu=�=0�<ϥ����ʪ�˞�:>��7�?��q�R�k�<A�
�i�����$�@�x��Nsu� �!G`���G;��{��w�Xs���P���_���-��%v�7,�v��w����v�s&��33����	��pX��V�x"��K���<R�V��J�e ��t\x�������3��%�jM3"��69��bO.0�����O�)d�<���<s�H�\`β��T"�iT�"�8aU^��Q��$�b
�
�b���`Â�:�iPV5�Ój�qCK[K��/��|N�V���`�y塍��ؓ঺�:N�Ε����[�ݙ���W��Sb� o��Pjҏ�ʘ&� �#	%����i�)JU���G��r&_�P��\��nV��^%�PG �ս�%�U&cS�N�ic2�s��lW1cb���l nF�� G"����Fn��>e^j3-]���>1nh^}8�t�{�� ߑl�, "n�?2T����dPK~)�;�&`�����*@3b>���'9]�4�͂��%�>fNZU�o����9�[���l@3����-^9������껾�KY��S��o�� ڷ�(&Ai��b���*���y��S���CC Ġu�I-t���>[���d".$���V~低��2�ij6QZ-��*�Z6ł+��/}tlS�
�_���{�x��_B�>���ZF ����XJ�৙m����)�eQu�B�d"2#�^�d�k_��3W���L����ni��{f �N�1����t�ÀIg���U^;�#�rz=�:FNm��~�+��#E�����H%�� �1���S�M|�Z�e#�I;dgvl;ʫ�� ���LO2�7s�o���K.u��h�Z:ċ���n�G��@�[Y���J�1��Y��
�Ak��}�i\ݑ�2���.�m�:{�.�t�^��:r�'�� a���Rʗ�v�\�!J6}ʛ8�\\i���IWqV����3���"s9u��hz��;�t�e�[,Y�,�n^�E��i5�r����9�WY�5PeE����s��g!LL$p.x<��,����M�?�UWDPs-�.��@�Ԅ��՝<3>b�JQu��|G ��	�7Z��Θ;!��"܀�����p�s���5����<��Jk:T��%7�D���O��B��8~B�ԡ/Re�.�)��͖�f]{s�KYf���ݡ�&�_�ݍ���$�p]�zA+O���V�-�!��o�i��JS�n�U2:����+�or⮣�15K�?�c�%�S�����s��eAb.�o[z�$��9��}���k
D�E�3A?���=lB6���5��WPle!}P�X1���s�ɨ�c�9�G���h�� T�I�z�� ��o
L�Q��-]�1�W61�^X�̽����I{��@�`?)$�����'*���,z��̶q���Q���^(�@1b��g�h.�ʕ�0���0�7?lt���cB{pM�.��Da3� b�|���o�<
�q�7ْ]���>s�{yO�1��^C��Lp�"�2P�F����3����]y7��g��E���_<a~r��i�?t{K8*0�RIJ[F9��u9]�{LlA���3I�����e�Z���u�E�^a1���JMF��wOqj�js��7_���k�-|: �+��'���uq����zW�K��$a�8����w=����iV�-���eC�+�$9�/�3��RSN�WS�'�5�S��PI�RK|�믦���Ws/Y�ƌ��$4�yTRwfF�\�MCR!�/���l[������7eW���UNFyPC۱X�!�.��0��4�z�Vg6C1TҊ���zt�(&`�b&PU���^����߈��&�$�]�2����\�2����>*�,6|��1�uȜ����_?��v1W�-W� �0�,.��+5��i��܃W/��/����?��	�~pa��ܫ;(G��O�/|�'�����"$����͆B
0�����Oj?�_%T��vLw�0�/��е>3��qCԓz��IU(�kߺ�Ț�sT�DH��ɼzI���M�q){�߹ê)r`0	߽~g�k�E�|������!���d���C|4s����ہm�9���8R�US���r�%M;�<(u��0+�Gy����Vʙ/�(���#�f�!(ܳj`�yI��j	mG$��<6bAn����!�+�B�0X�8��FЪ���;R��Z�H8�8̌�9�FX�������y\�ܤCF�V�M�-������j8��vG���&���!6o�F���f4�(2�$s���A�:;�9s�:x;h-R���o��Ӏ������r�<.T�����g'��#�[]�c2Jw����e�����P�q���^����f�ĺJ&^�dt\�lV�6�ܥYRng� ��E�=�m��Y��c_3�� %1�eg��T���ܓ�kxlܺ�$%�F�/��'!V\�A����"�7�-�?eJ�p���Jſz�^�{!䄦��\�*0��F����_�2�����p�ۯ~�L���*�2��t��Q����|�u]���� ;��s��t���k�:Ŋ��&�ɆƬ����e�ߵ�B;+և�(=$��P��-w,�C�K�Z�>hƓH#��J����>\������L.������a�ҝ?��f��d�aQ5��"�ۍ*��:�\�����3��`���n�+[���}45ga��Q�ٜ��4Lh��mo3�B'^?0��b�w1�A�XjB��2��|i������YIE��y#��f�6�GuR.��uP	t���Gcf�q��8.ym���27��AFɠ�^@�aQ<�?T�^��|�˷�sA�w��g��d��v���a2%�Ң���������J�c�]v�U���e���G�r��Y400��R����r��=��մ
��XFm�#g.I�	m[��-��*7P)-�`M/;�e�X�9fص.}�A�ۂW�[->�+�ہ�ݙ��Iu�[:�*���]$��?�p��Ԗ����>Od�SZVj7�+!NYҠ'G�ן��d�������g&B+���f�)ײ�<�?"��o���\�}p��PI���C��]4�t�zL�nJ���t�5v�&�D�yLԻ6h��ODO������b�|��i�c������\`�/2���X����XK�r/��Q2���ZH%�^u��/ý�k�Kif�H��۠)�I7��-��I���I+�c��b.�87����h�t�EN�4�fgX��}2	m�:�(���gR�0��|��/5
��kpI��5���f(� ���N���fq\o�|�ŧ���}3�xi6�"E�����G�֫�d���bq���	�p��e�$�X�J�ܪ��+�~���e	Ѭ�K�3k�y�^�Il-=F�w�(
���]ȕ._���BS%Wni���/X�8ȧ�xY(��8��?����5��i��|<���>��tԁ���#ݮ����=RՎ���\Յ<zj��-m����oR止/�(�3������g�MY0�v����ѐ�}�T}	�l�|���Ed��pVq/&�a�1p*����eEAR�r��[F���D�PU�lb�9��/>��]/,D!���b�_�)���h1#���f�w���U�$|�"�����r��`�	F#*'����)y(<�}�����Ūy:0!������R����*�Ú_I�L�E���b_pZqg�I��*7��A,�Ƽ&�ю���r���Q�Q6(�� ����pj擮����~
��[�	�G�����aS�S��i��6�&s�R���cu�����P��ph6�gl�,�6�y�R�{ݟ�>��4�$����U��e��
fWr既�g�2� ��&���~�G�l�¶JȚ�lU�ڇ�m�R�V5�'� �a�<�N���v4�y�1r+E��/y|u̗Í>�W1Ǟ�&��G�;���AZk��	�/�y��B`���8RvOp� N13�L���:���+Se#��L�s'�S���	����ka�5�X�m�ih"|?���"�%��Cŋ�&	�Wc�:��r�G|�{�,���6�Rd7.�GCRi�'�}Uf
Jh��y�_�	��W�%@h��Ib��)S0K�4&�fX��_z�[�@Z��b��%Y��7��� d�P]nQ�z�ӻSz�{-慻̌1�A48M�yv�p���j�
C��GP+-�ز�R����Ba���}��'. �{�g��n1��RL2n"�i���1z��6��%
N�`���z�;@���E�YW77���r�Jڧ �=;~��p��ߕ�h�-�,*d�XZ)�8b� �bZ�(Lu;��b4�F\���Ft_�{�mbL�Id7��H�w��^l-A��iת�+Vk�./3�i��ϖ<���㔽�?b�=����'W�t�t�u�bh�
�nEζC�=��0���� �ϻ����`P�O^U�/�I�I�X��~��Z��r����ŎQ����#��F�����V�W
S�N�8N�Q�+�1���?��@5|���|zG�L�XS��t�H�$���HEKF�5��3Mk�f���#�P��p��	�%'��/x���x�,������1��}pYׯ����0x���!�����ք�A�%!Y��aXГ�Px�D�C�y�#�����>��eoiy]�����7k�^o��"��W�	�I5]*V���nQ�5٠IZ�7��k��J�
R��w v
(9�W��p��R~�3�hR�4mG�"`9��ek÷`R�a��t8��`Ѝ��]_r����Og�����FUK�1�����h2�i����Ի����0�O��5o%��m~�ڕ��AC�� _�-���m�������y3]l��uϦ,n6c�\P�JP]�
	K�|�-$��ou	��N7�g�������ڼ�ޓ�P��-mt�.a�|�Ͷ^y�8�h�xQ�+N!���0�6�;k��-"&��-���`}�c�=��D �J������4~J&� z�/�������I��U-�i�J��F�g����i�L#�~�F�-+`	�oƙ���R��&/��tm	Zil�����>�3	ů��d1�.-�0�#7��(�HJ.�Yrɣ�Խ'
�&�G�!eΉd�y|q}[9���e�����h�ta����|�h�;��%Ds����Y��'�(�3Fk�zUd>�=Hm1���A���J���[�8m�EE-IXDC����i�&geI?��A�횂��VrοI4�J��%a�������O�bD'�4����(��yHl�:�K�6�z/��H؎�K����q塣Uٙ[�x8�8�r�6q��CXIK�?�Cu*��46&�ٌ|6�.�'U+�����?����{	hx�&2h|IQԺ;�vh0�c=9D�4Bɖ�%��b{V��Gh��j�4p�:� &��0�U�6�k���\��6L=��[P����K��"eC�R�"?S�WG���f��ߏY�4V5��9�&�Ln��5�.º�l�������l���֎"��X��C�L�Y�U*"��fG+H�� pnm:¬v��ف�N�k��b���(JW-M.bTb"�]Do�����@�#l[+y�;C��iN�=�&��9�*gz!��8n��4�S{�7>U\`�����ʉ+\�8&�O�ӿ9*�GZ����y���Ih}%D�+%h�[Q�ś,ﾒ��s�J���0�~��ߪJa�\'�}����R�^⹺�������u��W�$Q�FY]��0S(7�9q_��9_$R@�=�5?��K�� ׄ�����\�?Gܙ�S��F����)���T��̼��`��&2gQL=����<����w�ЦL��\��*d�Zjԍ$)�¡�4V�3|d���Βշ4ks�y:��ː�Y�q�8E�F�g��h�Ӡ1/#��qQ�z�q�S�Xo�2v:�ߖڽ
��&�U���#�������z���Uh�f������0�φ%;��k��X�x%��_�� 5^0�}�^q����a��Y����G\�sc��Ł�*&�:\ף�@T$��gk�u�P��ҠI�{�g5}
�"�G���[Ե�g����#c��P`�%������a�)�o,��M.���d��1��1�lC� I��y�,ڍy+Q�J��M������4�����U�=���nq�z��uiST��|!V�:��v���~W,�8�
�Y����/��p�q��S�Y�8/�ܝ� �ۻH�D:*�-Њw����7�s4E����q�-���ܳ�)
N������L�x�_uP�dQdwը"p���>�Ӑ���$�'6� �˝6��R����;��Y^�����T�`>7T�F�� �E W��)�!��?#9�]t�l���"�`�L"�P=��\�Rr�s=�qFp���ͼ#����#�a���ҌY��sϊ�z"��QRڐN�k�V-��c�*ʆ�w��$���[�����.P���t�z�6;2���k<\�ۺ|36t!�-�����Ya�����eG7���b�Qy����R�[��?y´�L�ð���k��7�%^� �V>�3		!�B��I�K������8Y���fL����o(y��Q��h�;��'GC�"
����$NWA 4��bO��KN�2��Qh�Ӛ/���8���翆O�mDw1���9�zg�RT�.�pΗ^���p���x�ި����nu�/P�J������fv25ß��Ps�(�jņ�P΂ b�.�c�������oҬ!x�j�/�|d��8�[29C����j�U�2�*�d��!����;KAs/�$򍪺�o��b��	��{���xZ���e\��>��?���~��r�9��2�3m<�ߍ�t.0Je��wV`����|�_..5oJ�Z?�b�cPQW+^"XN(�U�]���q]p���S+���6ɬ�ԟ&O����3J��bǼ���>�:ydOeG��bܽVSm��sʼV�B�#���s�w�����F\��4n��w�&iL�)Nﵝ��`"�{C̀�AA}����$����9�,�׊��,�c��W�	1�L��N���Q���6ƨ����.�L�<GYfR�0�=G>�޶��l	7�@b(
�(Rݍss��i�ߴ�.;�E3s�d�,���;�A���0iC�Ѫ���E���S(ۈ[�CrE8����Z;�v7X�����c���'K��u���"C���[`ۦ�ıt[�vkۓG�+F&H�4�;fG'Z\��{#�Mښ�Zߠ�1�,��L�R������#k����;��뎳�bu�*+G{��Su��oZ��#-���F��E�@�?��l�'��<ٗC'0�P�?�5�#�"�I���8��E���vo�����Wh�A�zhn~�����d~U�{�R��ĤM4���ֶ�Ə���tE�'�7 � �3�}���g��e����%��{�H�$�;�\ђ\w�	='��usE}��p�F����(�����J�$����a���B�7'��D<N
�mؗ�>�j[Fҟ@���j�p�j~Po�#��q*��gX��� �B�W�z7f���d�'DPZ�cI,��m�7�������b6���'�boIa3:��f���y�c,[�C̠��?7�mrs�-���*ՒV�j�p�+h��E�1K�(k� =����i�C�tN�F�U\��2��><v9�tS��p�2�&��J�M��g�i�O�iA�m(w��jqa!�����/�,�>�gL�F���{0��������� �go���퐬�h5L:�J��d���}��zCL�����1d���=-�r.�>�ɐ�y���>s����Y�hr�y;~W��M�w��?A,�r8��g��pMi	x{bїL�i���c�ʯ6�W�Xr�`򰹻���Hk�=yne,�r�ғ��x�þ�z��>��F�_xk1$z�J�wj�4�^i���+��m#h�艾����7�0���Z�ފ:�Cn���c�u��6� ��v�"P&W��8��%�Į���o�]?�l܌eb�,Cʉ���0%���GW�P2�.J��cc���"�3]�NW��O'�Ҫ�#��)��P!	*i�y�����L�����f�Z�w�K��4���O@B�j3����i�ܴ��������
G�fc����H52?Ȇ�=����(t$œ8 ��x���>�E��9�Y��� hF9}�s��`zH3+������,�1�|.��O��	 {��t�M�K�7�^���|�YBH�k�C�f��z��*U��@lD81�Q�Y%*G�:��(�H�D�'-ĶV��qr�#�<2**)sy���.r���(a��=wQ}��w�hfK�°�Zq���qO�ܯ*)��曒f��o�ӕ�TcwH��"��.��\���?�bЉ$L����4R��[��R�C�h�4��y`���cn���8�hg��@�A'��!���9�oH2"^߈$$N�刺���g�������6Z�(S��J��r�
{OO����t���fH0f���}�.�q=2��N�5 �;�foW�L�qh}�7E�XSO6i�]Ml1C�X6Ʌ#]6eY�*�j�l�-]�\�2	�6t�J8rG�"�p(����X���Lc�+��V�yG¥X�9ز�3�����<z�~U�>���%��^���e� H��b܆r��鯛z@%�Btl��0FԖ{�C��:oY�޽��"��4(hŃ��b5��m����1� y�Z1*���6?����Q�G��,}��H0��y-P�8�&��C@cI,?����#[*>p���8��,��J|V���V\�Y��[P�������6�8�ǻv���!ڿ����tG���n��9�ׅhY=c����i�4�����r���-�0�2����h���p4�~���$9���|�^2�I2���,5[���	O��ע��Zl�����l
d�L����H�t@���na����*����K�&*�t=c-�n�Xu��\�e<�X�Q�����З�%�x;���h��� �5?ƋS6�|���؝��uW�ƫgj��m*Cu�pqbE2��Z>�� (�#�#���N>�K4��oq�&6����t��%���Ϊ��`�Y��%|��0C�w ^����Y��}M�'�_�Ui�q ��I%Cy��+w�ӽ�}��|EZȠ1Hy,�tt���࡬n�t���HNV����Ц��eG9"{����Ͼ�q��WYT�ri0.��h�$�a6K�*��R1{"), @���K�8?j�`C�}��.W�S�E��[��P'� w:
3����"0EÉ~`�3L���(T�@WD(�)��T�Pw<cd�YKaޜ��m;<��;�}��*yi�Y'ny�B���ԃQ���U��bHu�K���{mg4eG$Lz�Fc�,��+�b��F��$���A���og��GN���vb=�v�1�ŵ����� =�\���R��6lJ�B���y�}�G6�O[-ptK��5�CH�ڪeE.N��h����Ӥ���C������׳���	|��D�:�q��M0����֗������)�;a����_ۜn��H��v�PM��r!��M�,v�9���G�<*�.C�[L%t��f��Q�i�FxTI���[��Da{���m���/�i��y����?�����#�T	�/p�_�}�l$#�D���Ω��!��!{���09S� �+��7\yw]w{��3��O�ڝk�$�QTͱ��sxU�܊e�}�\ ��p1THѳ--��8���+;����sKD���yG�&_�.F���a�Ҕ��� :��S�������F�P��TE[��W�X����<�5
���/���X��ܽc>2��>�6��()���N�!�D �+�
-/����o@�0�8"v�������\̍�}�@�7%�g���;����?ʇQ��`	�t�Q��=�+F �-��
m����a�z"Hp)r���g��r蕾��l�TFT+m�
�8B�-ٷߢ�m�[F���� *�� �R.M���.��5�c��tɹH��D��~c֖+bh���xC�`F<��{��v=�ȿ��ש ��pȕ��*��Qz�Ǡ �X%[$�`y��̨z'C�g�Qs�ž�2�Q}�0$ѻ�J0�vv�?� 
'������=��)�3t������Z�N�W. �k��f�y ���� 0��<��{:��_5�|�#k�\�;aq�^��C��ZlX\瓰�
�v%���h[D34�)�MmV���85�)��ulE�`��F�~\Q&�*ṿ�����|���=���Ux��<-�y�	�R������-�qx+��ȼXձD�`�-��X2�W裃��f1�qB�k ��g~�r&�����u	4��vj�H��jl���`��x/���dL֚F��u }5��(���fhC��Q����o��3y��;Y��Y�j7�[	XD�{eQ!���`y��Z�	��Lmu�8��^ [O��N�g��ΛC�	޾SeV��'�� �ފw�8�)2�[��e��N)���aLrG]�ψ�j��:.{g�0	FE6��>�Ǝ��O��E���~<L,70}&LK��_�)�f��~c7�	N��!&�[yJo�t�p1F�r�2}JC�� z�m@W�	{;���a�/ւ���U�F�4����q�
�X�Ij�U����zO,/��1�%^�{�������@�)?��C0Ω���U[u��~�Q*�6�E�$5/0_6<�nDs��iC�P�[ �(��U6R��i�ֶ�I��9�m�y&*�?���G�Z(2N�ީ�O}��v�H�7'��B}bm!�"�M�*ݳbY�/�(ݱֽ���ݦ�HM���,��<�~��ߙ���HL��遪��X^<I�h�
��N4�`CZ@���V�Wa+n�0k1�diP����[D���>5��*����&��>v�_��a�1��,E��d�E��8����N��]�����.n�2o ��5m��[52���{�%ڧ1@}���j<���A ��9rƽ{a�8u�����4�m���i�^��G�/Ƃ!]�	���5���7^�L���:���(-�.��m�^���%,Ӎ"r��,,,	�}W��S�� ����|��ﵴ���h�"��� �W�[��<\g���&������yI��͉�R�!�ť��XH�{Yߺ��o�ͽ͠���5K���?��I�d,�8�o'L}��p�X�������߶-��,qH>�����*�;�����z�W�g�&��#o����J7�m�����[����U$�Zp��
���'��Fƪ^��o�D����^��:e�'�op��wͳ[N&^���F���Lp|Ɖt|m��]�^�ݱ_��5�q�ܚ0[;u�A��wZo��k�Izf�Vvg�PϱN8���-�Ti�v�C�!B9[��`(SA���d�g����@�@���v��5�� u�����_�]���n� k��ei���<�55eR*��9,�2�qd|�L� Л�c����񴀓�Lt������L��]�i��)A���+X�17t��0�F���
� a�ё��{ڞ���ucZ�C�~��)j6J��Y� �?x�ޏx�;x��R�� 1��!�B2�tB(�9�Ill��ih��^w���ޜ��$v�N>͋�p��l,��v��5:o������1V��4�p���o��L�h#r]9�AI�;�/1���G�(��0ݷn����[���F.�6G��)��ߵow���B>�˧
�eZ�?�n6nN��A鄱�[lip#����A�s��K���!]���bG���Z�ؽ+�G��uݏ��#y�A���MM�J�$�r��
.T!{���������o썦�!��"O�y�PS�a�.J����[���]$+q��	:/��˛�����WMU�{Fe�ڔ��0*m��B��b�T���2���px�X��p8͐��� ��Q*��5��p
)\/ס�C�4�[ϸM�š8�%	�hA9�u¨{��3o�D̡��4��M%�-����*�ևx��p����<�R�F�'"E��0����.�q\{��ʴO�R=]:�\ɵL�CL�	�f�S��#��\��{�f�6�@���$�b+-�w��Q!���?b�]��5=ӹ�!7Ty��a�΀cEJ]�z��J�� ��)�`�?��cNB�f�d�=?�(kQ41C��LJP1��g�j)Fmy�rUA� k���+&�DHRSmw�1��@�Ylt(E�y�8M�����u�'B0rU�?b�{aXew�@��}��6����=�Z�tu��Ӓ��Z%%��Bv��|��/�KA�"S��f����[:?�y���K�Ynz�<dx��s1��	e�RDO�'�͂t�"���~�"5l.�,����Ŭ��$t�
��P�QD�gwp�-��h�ݴ�K�N"	%c�}ȊZQ�lG��6�*�/���B�,���N3>��tu�[ �,u��Ƹ |B��h`7�"�(Ų�R �'Un|�P����_�M|CWy�i��$WO��![�q!�В�%K���ú�-dd����ŧ�7S{��4�@�������+��f��6������4���L�p��2��!0wD+��fs�ww;�>߹��p�\�4:���+��D���"݋�f���I��v�;�&5F���y�-�[�^�bq�K<�����E��:n��)�gJKކ����1�� �*�̗�<p�x��a��FǆT�Pm��V#P�:o�c��\vH |�D��A�����ze�P��1�<�-k/1�A�ڙ��cY�����S�.
��4Ƹ�5��oZ)US�$w������B���{N�TF��Z���)|z����O���-��z^�\�i(���F�N�Q܃�KD�I1�1s_|*��<�ņ�l��m'1S�p��#v2�We�"�6	��4�\$S�j�?{>M��j�zӌ�K��!��S��g���`Wi�6���QX��tGg����4��nnl2�VW��!�b_6�[�B�7ݮ����}���a�=���7�=����S��x�/&��;I#�����woL/���8Ip,��}#�n߇���:��۲�����E����=��Hځ���-��	���bҪ0J����k�hb�g�)��Ѕ3	�p*F��>n��P�I����	�8+���-��*�|FQ�-���}�<�1�v[��N�e����o�u��;R���H�8�5��oB��V��~��]�M��K��|��n�+�x�*���Io��t�Ed���mL�i߽��icߍ�%@Q�{�x3Z�k�t�-��z#�8�)s�o5	
�c�O;/�7)�R.-"���u_S=�!��&�H������v���������ׂ0b���!��q2$�CϘ�M�Ԙ扫)6	����v=����`�-E�=6I��9նA���vV�?���7�5n	k	,W��6S��5u-���=!V�n�Ʀ�WC����s�J�{��"���>/T6���F��cO6h���^��U!_Uh�`��>*,��&u�p"1u&�W�)3�p��_<`N=m����8Ϝ�  "���r�C�e�Ҁ�W�.���lм1��8�	����A��.:DHӜEJ��9k�?�����#�e`b��S�ѡj�Q͒R�-��v2h�g����:�^�2x�pAL<�3ULmQ�i��Y�Ax΂����};�\qE!z�Q��4g���+�kc$o����"B�Wxm�����(��忬�	�H�DT)���(4��{O9��B���>88�d~8pٍu
Vs�p��P����5���vzy譌
���J��O����~���{$�T���K��^�!ʳ����X�2�	����)�rA����-����g�(DP+B��