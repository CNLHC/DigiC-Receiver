��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��cJ���@n�s�bshG#]��<p��*dP�fʣ ݕ=n֝�~z��P��b���
�j���	�oF�VVL��^MZtm��.~�n��M�rV��oe�.y?fbA0md�5����0X�13O�H^m��*$/NK8�� �ʙh�M�%���&����&cj���fXn�]Ѕ-�M+'����Ɣ7�P��߳�,� �/F���4���3,=��S�خh�KUI|+�XkJ�nIث�6��U�ֶ��b� 
��N[��pǳB�N���΁����F�	��r.7ҖЧľ	�O1b�k����\����'��F
1~GZE��T��>�5�q��!;4-y*L�wfs18&�xI��A2����A"EM�V^}|L:�6]�`ʢ��}��;Q�G��vy;vˑ�x<(�����06Q�U�fÐ��fh_cN�U�ӎ!�T���S:<'�{�A@v�]��ԃ�VqZ�� V�8���H�-.� ,�=�+e���嶇 �Z2)�q�L��.��b^�?L�c@Ii�	�;yH�\���������οpy�eD�2y�a�[2�RS2���Q���K"�N����^��U�K{�����r�Tȥ���V��ݛM^S7���L�0��4�[��� �%���ley����i�/��Er��.���ƹn�|^o\̕�,i���Q1]��B��8$�<C�e#4�qG���,�_��$�t�!�\u���r(�t��5��?�r0к����D�d���#���-CG���7�l��?0� #����<!bNd����O6�r���ժI�ǟ��|]l,�ES�3m*��Q�����Z�� Z���Qx��Ǯ����T�W���9N�>��g��TY{L�*�'�k���to)�]JP�,���D�
���9"���h�g�g�z�Ё����UD��������o�`Vκ}�&`mY�a���-�meb�wŧ����k~���P˄��V`���X�~����x���9����=�=+̝2��1d��ڥ}�Q�C��]��,9���x&�^N��,mf�<���	pP2F��`��l��$��	>7J�)o%؂�!��?	(�Ȇ͊<��V�5�/���̳�e�1��VH��*d��y���&��ڵ�!]׌L��l�wP#hj��\��Ħ{�d*њ��t(F 8k���뻖�:>!�~ovHaR`��^�Ad�|���V�:����M�_]�쉗G��+�'P��V�G��˟�FY~A�MN��l�U�U�iZo2_������S��[N�g�z�X#w��'��a��K���w���e�F%P���C�~�U����ފ��#���!�yW���Ζ/�c��JŜ���r�X�ߙ�Rh�y_�	w�w�H�i°
��1�ݿcxcaF"K���d�����ƲR�A�@�Ӣ�]p{`���"]��-�~ʤ�9��UW��wN$�*VѦ&��'¼�a�Dܚ8����5�N�6�M����xcZ����[��Rf;�����*�q`�c�뭣�����H׊��#`5�=@RX/���Ԑ�'�&- O))�����ȸޗ����0�����2.~��<_5%�0�B��7���U K��/Yj�������ej��~S6�� 1��!q:�W��n�,���+���v�~�1����
��f�/pƞgAA�ѮI�6A����;�l�#��-��]�i���d*Dє�2�ݺ$L�Dgd��t�������b��1��3sъ$N�[�����3w��-�23�&��Y󄅪��3W������2��sS�ֳ�i��dR�޿C��Ӷ�� ��f�[�&��\��y����V�_�+���W�wN�Z�uO���;��I�	�ݕ�-��[Z�������&Cl����O�纈Y ��U�t����:-� �W�MUܢH��*z��
˘6������;:ܴ�����y��� �$��'Y]�e3R�\u�
ڗD%?��b���t��-$p� l�14��hrZ�z'� P٨���ɣ�H@û���Zy!δg�)=���>�����
�\�Q�k[gy )�[�i�[^$ q���b����j����T��9�܈A�C�w�PL���S�\��k���b'��0�������Z�Դ�A�7q$#��£�o
���J"�rG:Fa�I�BS��;�?�`1sJ()��n/"uҺ���o���NX�؃������Q�t_y��%�(�G>OIc��9&�I��!���H����˧7���{���0��U�� <Z<���6\�P?���.��h�rPܻ}m��A�%U��d^"��۴Θ���7��k(Z�6��D�o3�_�����ƕ
P��Af�?[w�=l�:����iJqp�5�͎��Bz��
9��U&��ߥ�7N"��e�㎋|�$.͌��I�_ ��ĕ�57�|�i���p���u����&��7�8��.w:����d��0����(�`��g�)p�bR�i�zCh_;Q���(4��[�l�ʞ���5��uz�2����i�C�� |nNfZ���d�R}`/�%�&�O�k���Q��9.5�OA� D2�:oOh�Q3Մ,Xmb!���p5�TU�#���:�߈�<�b
�4�52A�����o���!{�ǻh*����V��&Eo��rh��)��AL�Ѝ����8��Z��t�[o�AQX%p�D��|G�r�OG��T�fhi��@�R�a��D�l�lOU�n`v�8ȕ�{���-
�El�s�V���o�y!L�ճ�`(%��qCAvK��P�GU��	�Wq�T���wsC��+���L4�n^#�C����<*�����۴�_��{th���]?l�.f��ea0�a.]�$CW��%ڐ
�0�����@��ä�<�\����r��+ֳ��Lފ�����v��K%��������ү&GfuP�7��ة}xD��� i�	��Fb�>+����n�J�+, S���l�R��(H��I�ϣ��B9�->�� c���+0�D:*MAI�H�� w��e�Y]av��iǫf$�^a��ԧ�W�H����R."T>�?����S��g��ǧyȃ��o�ܲ;�*^a �t�"z��CoЍd1��:�t���7eI�?Ib9��߭�vT#R���	"aj�E������h�0��>�h�e�/���ч��C�k�	���8.��7��|°��Ѐ��ȄEl�} ����f��T�eo�?\�����Ȟ�q��@��#���oc���g7eM%���kj�e�/,%�b\�R)�A��*�2�ɔ��>��Ґl�?�5*��,W�$��2�E�^���>
��6	OK*Bz�!A�-MԳ��>nc4/D0�7�Ҵ�9E�7����J;[y�u66�?�bb��z�޲�	�`�S���2��=��eM��Y�$��?�v���֙>=�K=Y��o/��� ���Ȧ��q(,Vx*�V���*!�b��4ҡіS�IK�����U�#~{���6�>�A�E�R[f�.�E�]K���4u\f
l�^��l�ج��!�,^���#W�trO�����nVJ)K�;�)�1���e��K�j�I��qʾ��`/�K�x酔a߾n���kf֟��pR���f�2(���V�mf{	$�U�cOA�ܬ��Y-��(3%bLW�	p=%\Ǟ0���ե:��M���Y�oЪdT���d
@=9��h~��d;בnN8>���_�>,�C�lƚHdgx~��A��<�g~��/��#<+��ٶ+*�n��N��������lC���N����Z���"���&9L�o��q���I�&�$J:���VW�4~ ��\3�����xR���=�yl�Խڝ}�f�)pB}�{b0+�f�
��P�Ll����P�.X�%�H,b�Wp�2��;��oƚ�|����=l@�5K��N��Dn����-����|>��u�kM�b��*����Q���,A�L0,�bk>0��I!?�2t���^��ɆW�����U�����N�1y-o��7U¨��.�~����	���6SQ9@����le	z��DlC.ڳ�[w��#�7cO|-�2�@��e�
����%L&3��x�F�T��gJ�eP§_�ս*9��m��m��s����K�C�������q��c����$^`����:���eC�߱�8�¬���� K4P�JGJ��!P>���1��$Z�?��n���`�G���$qP���fVf��4^*DR{��2������{���+���4~jt�I�5i�>f)~I�W���\�����i.�5R�M3߀|��ქU��mu��u��7�FV,N�`ZBQ�!�ِ��z×�.F��_5��@z����X��씘�_��i�� ���Nqz'��{�ȬQ�ͺ|@�h�?��T�Ւޮ�3���By��nJ���M����&��4<7}\�����Z(��fE	4E��gJڑ�A��:�2���\ �d�0��e�������f$.K��tT�D9�*�����xf0��D�Ҽ"��,?��x�=ZA����9uЯG�F�y�M�Dd�7�ȿ���ک�ے�H!�-P��pĳ���Peq��AcH�����������Pߝ"���{bJ�>&;U� хA�x��~/�cr4g~���>]�'5N�8��K��8�"��qpI��x��U8@��@��_�q5�2*ֱ 5#iA+���e������	�y�)�6��"K�������:V&�oP��$�Iq�h��\���u{���"�;�1p�Y;W���˞`l �A툿�/A�Ւ�B��^�&����<���:�qaL��#˅�[��L�w��*�A���qM�8ڵ�33XX���V�5������S�@߬���&H�ت�;!���D7U0���z_�1=���=|����FO)���7���t��x\A�ݮ7o�����J��ew��u�:E������̟nlT��^{�	�۴�D�f�PU|(o�}��vl�)�>䉩��!'ӟ���~SjT8i$|��}c/D��}��P�� �sa� u|�T�\����\��J'	h@ � ��=�zk�>��}*�~�{c���µ��fD���xS�Ǐ�ML��Y�Z��1Z�JhS�,�cO'ݴc*P��}i�/rFLO�l�.o���oBz������|�l딉������eSO�׉�~����|A>l�%,���ъ=��*�Jf�C΅q�v�*����̫�d�ۈ[-{�8����rĜo�W�n,Z#�#h%?�����^�B�2�4s3s� �%H�u��Y�v����
�'�c�A-���Tk��)3���﹦9GXťG�HKxvKF�݆I��p|m�y�N5�8ilR��X*M�IK
�Z}n��)1���!��z�-��!�{��*��@��6���D߆���@�RK3V�g���u����i��.���GP�D<���/--����*���>�M�8�ǲ����&�B�~�Oo_��CS@���hf%w\�z$;����`?��x��n�ŏ^bB�.T�fD�L��� Vr�&��}p
=zɤ���7�3�C�(3c�uEo8s�_���b���iJ�R~�0��؅�58tJ	�ժ�k��"^>�מ���k�e�xKs��T	��(�9�A��t���p�/�-&�M�şL�*L!��HE�t
�\�=Q��6�r �P�Ӏ�v�L%>g�J��b̖�wZ�u��K��y�N��{��Z)g�Y��.�7\c��&S$��.�%���� �ņ��I�\���k7��N}yX��YMXO�����T�>���¤��x���:!�Q�|��,���NB�5��8��	��?x";�;��VxZ�ط��[|e�vd	��qU�ȳ��P�ބ�7�(&Y���NQ�w:y���ؐ�腴�g!9<4�?P݁��$+�t54�AU2S��pJ�.��j�Y��T|�d"�;�J- �M�@�-�Mf�mi6(���	�v$+n*f�=�r1�	���EQyp�f�#����	���0e%+K#�X&� �u\�=��2ߝq[���H�p�/k"�ueڌ����^>`;p'��ְ=2@��y�U?�B��辁ZuB5ػA���Y������ �ao���lOKۤ	�~�]��^���7D�,)q�H��)���l�}�~�"��I���UO	w�:~ˏ���A��e��QBEH��{���J�ֆ���^_ԓ�No�L���3��k�;��0�2�yh��YCb���3Z@�X�;�"9	?���j�}T	b��ghL�D�ص����E<ЭR`�T���O/`�O�}"�����`U8Y[|��H�124�1����G܁CJ`^����49���ܸ5��O��[A���X��Aj��N��{d9ڮ�����]�,wtwQ���B'�w	;Y6�'��WV���_�T�R���8�g��AN"��*.z��d9�,M�#�cDϦ�����C\u��l˯���T9B�bX���a��E4�0�{D�vucv�V�4��.�\�P�]��3y����p��A��/F��ߌc*ڔ�VE�`Ƒ&�U�)����L��88=�t�s�(�n�j�����G��W��eeB���$��"�B`�RL�����P��/���\���א�*�dn�%}!C.2� �q.�.��]��"9+o7�8  in��bEػ�:��ڪ� �p���op���E�0!66�4bA�c���x���O���ah��R�I�lMЉ���.���Z�y��@L.�yae�I�}��&[��G�$枋4�ؕ��q�ău���q��2�\
O�>��i�͑g�(��(���l������^
�J��'@�{�\d1ਨ��*h��4�;�b:g��|K��R����͂�z�M����22).�c�8��M%5)M��c-�W�rV0 L�*���v��<_Bڪe��,$W�w��e=����Tk�'�*��Vj��5SS�T��2���m�N�Ɏq~����8-r�`��X5A$?2e�$8��G�<3�g�`�فEQ����5�&��}θ�m��f����J�-8bPR��	�n>XC��_��9U��4TQh��s}�ě	}Z�B�ܠ����<%O���`�y`���݆6^\fViu:$tْpw����F�"Kv�7�\���+��
����6rW�jt�r?+�+io�������=l�.�=�}���ص�0��es	���e�g�M�I�?M��߻��Lʍ����f��[���{�4��W/��5(��3��C�b`ܪ6�S1y1����*/�`~����7�nDopp��Q�uy���J؛H�bRm��>4�F,�faj�c2�	ÿ�V��{�f��vƟ��H��r*�{��;U�BYt���3����_���f��8�/P>�O�e�֘��m@C�ӼLN0�*>Bb�WL1�T^�U��Ea�u#�M%���19�~����u$��v��	p0��(jeڀ
�/����rbb�K�G��Cǐ#ŻJe��pC���Ì�]	)�[�
/R�d�re^z�Yݯ�mTF��W7鳭G~�M�}�WN #mo���§�)7́�}Eq�WL1'w�ʛ?w�&g�&��
OT�yAdWE@�Ý).DpD�k��8H�)ȓ�g�W�K��Zȍ�y�Ėr�������[mI�s~Պ!��5��&�#��O�~?�k-��/Ga'F��|#�j�������_t�9�˜{yT4�����rl����b[Z��>u?h�M��W;�0F�n}C�,#��˝�G��	X�C��5�뮚߀�d�[A����Z�<�twE@l�B��H~�a��t����'���z1���D脈YJ��=���iXb7\D��M݀��Гrd:d�bE0�s��M��Jc�d���<��Hq����?��A]H��"t�|إ�n%\����|�HPr������������/m���5�6�6ַ3^ī�Xm����_Vop=��(6�Y�|��H�^,�Uǵ���fʚ��5ʼ�kY%�̓#�B���N+1�vm�2�7P��r�Y�s�b@a��
A�47�H/,�`���^�5��H��#Ky�|�E��-��w�p��P�p�H��y5��nj�����u���Hڜb����u�#��Ow��d��7�9��G�b�(�B�&�"���;O�A�W��M�Ά5��@��_������V�]r�֦f�`uW6P��nߎ��{��5@�8Aƃ%/��c�Zo[�t��'�ʤ��R:A��D��9~o��ƅ`i�"�>��.Bs�Gj�Q%����g�Q�u"Ԣ��H�W�4cԇ�}E{-�qvSk��3�A�QߟFE����Y�^,�������C�4v�ɡm�u���H�$/0:�(7����N�6�$=5:Ό�-���h8J��C�^+����S(���1{�S�1��݅gb�#�F\% ��u�
`�;��p��Y�6o�*&�t�� 	�1�V��{�T�(���W���=6��w�����J3p�f�夛����;d��a�a_�v�b�J�f<�һ �+��%k7O@���T�\�^m�h�����ꦜH�Y\u�@�}8&^��vB�%R�U^�N��/�d6�H�w�V�g#4z1KX�u��6�-ے�G\tY�_��uz��8a5�A��%��[inZ����f�䁊7��*���N8*U�ޭ}\>i�a+&p7aopca�)sd�6_�]<�r%Z�:#�����+�����v}3���c��s��7�i�����hȨ��ZKo,Xy�*u�)��J�3^��͈�? ny�.�����0u����Re��u��^(�GK��1������*���>� C�6 �}Ԁ�l�GPeJ��� ��u]��X#C�����2%��نլ�4d6F�
S9�4�� ?1���q�=
�>p8,��w�a0�u&3�l��8�m�� �ײ��6P��N�XQ$����^�.��@�dW=N����Q9kSV�y����k����>�#*��!Q�D�D-��u�e�R��}���������O�d���7��<����~�O�(_6hDi�F��_qD�N��;h )hw`�����"��ad������oh������X��Sm�4O�K�N�~f{D�;:sU�N(k32;��M����Ӯ�h�F<���%L�=�HȰ���l�Ą��0~��;IFfi0&f�T�9��f���&��u��ol8,��s����!<�B !@AU�t��mt�:�#y<w�����R��gK��*p@�s��5��P		�2�f���{z�X�}f׌��@�1Qt2E��R�ܟ�<�<��b��v��E�U�T�$7xpn�0�.Ȃ���u�!�S��1ЌJ�o�˲A��t�pز��&5:q,��h�@��!��w�;��0^�ha! &&��P��㿡�Y���Te/�n���@k4|?@upGL��x���
n�6T_�0~��	-7��|a��o`���J�	�����<=.�5��BDF�h����lh���3r�*�$�ZI�0s,���ſOt�{��27z�������U�n��Ǹ�⫉-�{�g<0�Y֛)&��,4��A�g������'*8�hr���7��Hr4����uߊ�w�sDN�3Q����83=4��+�_(Z�cj��)쨻��A���n�)��6�S-`��xO��M	a>r���awE�
��5�$��Y6ޟk���E1�A3�N�M����^�<we�����o�����U�����ŽR�k�����1�V%���]9+�p
l{a��^m��R�25��p\�s�)��tN��ĵ�i.h'u<ZiY��S$�~	M�������2'�ff|�-����`�Q�TA�.G0����Q�b�kn��*�q&�o`@� isAY8�$��A�`KT�����Q�x_5+�"�jc;=K����0!H��c)���F�)�.]j���u�Y�����Q�;b`������v9��х{]�y��G�8�S�_f�ғ?�}f�_�~�m�CQ�A�,�('���FL0�0�n2釞�t���x�U/�ۦ_Z�U������g��9�|�V������M}���S��8�-N)����{Wau�-�5�95)_s��/JL�*�0��Cu-迨ٟv0#^�L����]�K�!��3�QZd�6�GQ����,��j�G&f�%e �q2�'�}t=���$��l���� ��&�\�U���\"��EVkV���<5���F^;voI!��f�R�,/h�� >��H�p�܈O&[y��M�(�ID��:c���Ojm��Y`��Rۃ�F�*j�;gN��qco>Jd�:$�LT��#���i���a3#^.$����Te��"�O�"��	贃�u{���r���D8�4&yi�z\��K����CE)=�l��bkV���*�h��+�N�,X�73�b����BJv2�h˄H�5�2)%����۹Z	6��ԊL1G���d#���	��:�t��d��VA�-F �Ϝ���ۆR�c%�+7��*q.vn��}�J�y. �|��9g(^��EtL�[ò���Z��� +�g���bvgdJ�yIzC��;�(��:&)'up��fJi����� ���2k'8�JJ���P~�U�_i:잤�_b�Ng�1Ԯ��'I�I���B���v�� ��B�g{���R[q{}֨}5��9��v��Q���-�c��5�Ǜ�k������v�6��rh.�3�C ~)�qoI��g�JM!�!Q��{��5�z
Ξs����(����SS�=�r#i4}P�[a��a�Q}�������a��.V��/~�,V�}}z�|�h/��:w�gM;<^r},�%��yhbU)
��u�<B�w=�,�g��j���.�_?�m_ �g�Tg�H�4p�0XذJY��Sl�]-O�碝��!m��9��P�t�&�_�s�0�;�tc{���S]+�����ܻ7�L��:��]_�9����`���IT5�WU�w
��az�fF�A/gT��N����������P��-��@{�b�I�L�yG�����_�L��cY\�r����o��R����C-��=���V�RZ���fp��	PL{���㬀 ��t&!�>�o c�X�99�4�P��������7	Měԟ=%���q�'����kE?^(]�Eb��ج���t.�Ѭnr�[�w��4N0�\K���E�4OaXC|����O����� �8��s@->ks�k!�z�\K(�{��=}�ʘ$���HuͺՀ��`�+r}f�j��`�B��9ŧ�YẐ�w��i�B�d
x�Z��I�? �.����UD|T���� I���G���M[@UF������s�eM��0 +�6���l����~~+|�.&YUǙ˵K�'$@�ꉋ\d�[9[�͖����zR[)!�+R�2�v�]#�$��N5aWy�����֬d��T��Zq����9ZѯQftW�;�"2)��D�-��*L�!F�ɵ��Z��Ũ��C��?1]6�\?���$:��|�2F	��}�_�ށ�SBO4�7Y�8�j@���,ys������(s06�W۶�aE�k�G4~�G�8�f����fV�����p�մ��*��wfI�M��F���4h�E-~:��[}�k�H�H�"s9C<G8�3�J47F�3� �-z:��zt��jkjj��3ӗ����:�I����rQ��A�6��ԄQǡ��K*ӝ�"\��W�A� LSyh��lΏP����=͆sw#.K�X�Im��>z=�KǺ9f�Q���b��kedҺi����j�k�o����7�s�_X�Un��
&��u��FѲQ�mM�mc����t�W��o��������M����yuvԲ�b7)�>tr��h�:��ǌ��JCѨe&�2Z��K,�<=��̣�M /jjR����c�L�jû(t[�3f��f�ң�C����ͷ,gT��e�.�^m/��}�d}�"|�1�ԥFE���������
�'R�P�;���eJ}���:����zV�����������S�|y��;����y��f��Eg�3W�Tl�E���b��v/r_����{H��F�P�B��H:��^e�hp�e�'M�*J&������-�Q}}O�b׉���z��&�!�G����6O�7�9	��1h�5���~�Q�J�PJ�/����}�����e��1à)	M��ڂ�X��s�X�ӢOP"��,�=��o�f�i��a�U�q�M���:;�P#�#������:E��o���L�zOϢ9��[|!�Eִ5	,q~l�C��3m��Y\�ٺHs�!���HPQ�>aXF<6K7O�P���(淟AQ��!6���x��8�_�%Ď���t��ƴ��R�!�~	y��*��7�cR��B�v��r��<AN����Ǭ��0	˔�SĄ�u��0�Ǽ���6�V�#`��IEQ��tY���¼����I'���4\���@�_��b�W�7=�0����km�s}����t�0Az�}if��|k&r��#H�	 *����]�ۄ���^�������' ����%M������J�K��"`�x2��`��y��!=;m�,��а0��E¢z|*�;��=u�4���9����\; ���D�/���M����0z��#H1M.�(�C!0�e(�-fHu�����!�y��9/o���q�DԱ�OE=�ܱxZ���K��Q~�3`�p�W��Y�����d�U̦�D���i�/ko�$z������
���E�_����n��.�h�%f"|�6M�\� L#�\#�#��|G�+���Xǎ���Q�b�:���
5���]�����6��x���уT�ka�Ȃ�h�\��z�] !'������W�"��Fm��'��C#�U��6K+&"Pa6���l�:��!���8�ԏǶ]m	�#�\�����Q��/LS�������2�'R[o2�L������k�����[������WՉl�-a3�٬��:pY�|���Q�?}-��ei�%UGF�u5�N,3�qO��q���x�M�n��;�)��~������K�6[=��5�F�2���M���GL�\�qO\�'L��nY��p8
��S�3�����yrmC���we�_v�(BG2ɢ	�5ՠ� ��VO��q�Z?y�h��6��E�����	a��������$�_y�Ô�>�4�ؤ��l#�"q�Xy��wC��{:*���5y�f��1� �ٽ0�w���a��]��1��PZAaIk���y;W*�p>����qӈ���?Hez�c��5Y�G���x~�ϙj�]�Iw9G�/�,�P�	�[˽9Y���$ϑd��ū�f�YB�{��>��L�t
'@���\�����LtǮ�*2����8`l�/�x.F�����e�k��.^gY�StI�XF�OvM��T�%�Bn�\�P���z����F�g�2��Ms%�dqRϽWur�a��ӻ�؄'���# (� ;�>.`����H�{�ش�9�8�Z6��jr��RV��F�w���X����c;"g��5�I�A<��j��11ᡢ��Ay�O�ELwXN�Ex�ȓ��X� jQ�:�m�5_�-��,)�V���4��t�z�<69��R���=*�Z5F``�a�fk�'����XP��+�٤F�����8l�?E���񷝷�����2�{,Z���ʟ�u�.���&��?��v��}JKe��K�V��u]rF=tm�Ȩ�4x*x}H�I�lr� �*y�"2�6_.=���r�0�2����8v���½ �(��7P��������2|���=��m~
���\::��Ćz�@���;�N�2S	"�Q�CwHH2R�[�kc�Is�ّ�*|��xu�0�C��f
v�O�����y Kp�?c;���h�䣤���fӹ)��}NG
��	k���I��b��&�q����Ѳ�n=��?&���$��N��XAp����[�{8�#hˁ�6?��qt<853,dc��$2'd��Ԙ��0���?��R*�ܜ}/p��3�([k0��a��ǖ�u�b�E`)��}̻��A̥��%hCK%ګJ�E7�.��Ի`F��˟ރ��陋7��LajbB+K�/4��	M����% �"�dT��%�f����c{J]���(��̺���t�w�5_q�H�s*��9�Ұފ��'[t���-n��9�mu��+⥧�^;hR���]qh&�iTĂ4ef�Xv��n�n�n�uCj���G]��y%�/K�G�T@�k��b���}] ���$m���[�|G��/4^}��p���d�M_[Δ"��`z�*җ$�,�C��]������D�ϣ���C
�!3��.,��nM��<�w�r�]^ܤt��5Wg�驘!���I6tfad>:���/e�B��Rfd˵�H�yJ"��쉦R�ւ�]~m�9�4�V��Ӵ`�C�-t���OYd�x��������Yf���|
��$��E�q�F�m�i��=��G�����X��:��/%|Bp�*�y�4~SI��1�W���Z�6�<�I����e71m�DA���\D]��!���ii��L����+8�o<x!<�ӗT�Y�fY�lD?�O���7u4�+�2�Gϱ�J'�I����sp�bg�|�{l2y���3�lTG�E � �RCZ��Lә����n��acn�A�Z�R��@]"�h���>|��k��?�����y��0��WCj��-�@eY�#�����d9�u�x�b"�O)�A��XR��h���W=`�BR�wEJAKɃ���ݝ.�Gc7�� ����r�Τ7�y�l\"�����-��g�+'�7:ˁ�_��y��s[�IN�_"�U2�]��{����rR��gVJm���zc,H?��/E�[�C�UR�5o%�?��Oț�.E����~�Z��,<�<T3�x| �k��|���:vC�)�\�L�nϡZW��3F!���g�O󜦩K��H�/(FQ�F�w�S���uIZ��<뼣<2s,7�o〈��� 80%��C�	DIM7��W!�TC�x�"P�!�%I[��${��y����,F�s�	�C~��˪���,q�����r���Uʼ�����A�����3��٦}��r�����+k��=h����UDr3���ELzV�'<h�g����'�ǰv�Ȼ��IS	�%fC���i���b�R�F�#�����s��C9�?֍��H��7�w���7D%��Vr�)�4�AoO����3�̅0�^n��Õ^~',�v�F���am��0+��
۸8!��S�F��왕�������K�.�	�����y��Z ��O��}sJX�E���3M��}œ�]�ZΑN>n�G��:[���x����fU�*(����FŰ���Cc�I#V1�2�*+2����� r�X��m�7k������|��%: ���~��Ub��ل��9�{�D+/M�t��.XO���v3I8�J������M'*] ���q0����/����_�N���,��L̀|Di������х52�T����֝g|D�)�u��0��*$��W�����QW6]o7�4��,������YS>�|n	La
R�sB��Y�JM݄�ˤ=��f9�u�c7�D݈�ǹ��VfCt��Q���&��Mf����I�qP��3��d�����L�KɌm��Q��!���_��ʷ�� &��5;V��
�Nju;9Gh��dQ�o����'��X��DK��iTxZ+Lz��MT5#��D�M���S:��W���P/}[�U@���v���5����)�>������n�&�|S��#� +%m����8A��7�èR&c�9v0ڳ�L��U���΄N��L������ז �-��>&~<fE. J��+���T�����뢪g=�j�fe�_���eR
��ޑۘ�z���]hO�贏Y[���*w@�9��s#�v���	s�;2���0H��2�ͅ�<ߏ�@��Y�i/U��GC,��&I�P�&o�ϊu= ����e�h\,u�d�ڂB3�l+2��Vy�EX.��Ow,	�ͅ��J�R��SOr�Ċ�1D��/�CwRp�6�/�O���ؑH���-�w�#32���A}��4�tg�\<+� (_ ����;�Z��:A"W=i0x�kaC���M�ɜE�l�-��v�VyT�T�q2MUZ�9}���ùoa��p��xZ�j��0U�$"e��t��:"_�ɑjp`7<q7���K'ׂ̞A����?�ol����^�A� ����Re�4��C�Z�6%�4�]��ع�8r��륃��d��
�'��4�����v��ex����r��yS�v���*�A�����=�C��[F��H� ɦi���P�����L
`��u��8�ɞ�,�V�/�#�=��DJU���>�&�/��D����ּ��Z���'I���)Q��Ӏ�������5 �Y!4NB����.������߲��}��	����V~uM݇�X�����6	G�Y{ˬ����%sJ�X��GU�o���s�]S��M^g'�7���Ù�F`a���r����I��#cW}17W��kV:H�=⑊���j��=:-N��0�f�;�w�Ũ�"t�鼢�~b!'��w�����ET� l�#��Ջ1_
`�$7��.2>�[0֝��ˆ��U�J[�zpkr�6��Lcҳ�pBk��J̵�΍�Μ�����ffH�i�%j���=��[A,�����'�~	*Y��� Mk�5��ǳJ�H�,P����Z$����1+�6&������8�`�k8���n?�)�1�2���5 �a��0\B����}3JP��i�����Փ{փ�(���tgb���iK!��.�i&�^L�K��4#�+��ܿ�8	���9+���d����r�g��s��d)<�r늰s�}�\������gy���/�f!�B!$���n&c�M��4TL����r��i<!xƮ2ޗ-~����Z0��fs`0�j^�j_�z�ŭ"!�u�T��b	����~�k��,/��ƭN�A��T�5��}�)괍MO;'�����z���(d�A�fo��eѭ7Hu��������Z�NMŹ�#M��T�g�C�/�����c���&�B��;ዳ��1z�la�M�����Q0�@�}�e$�(9r�J:iÀM2)��e�q���N3b���o ��l��H�����ʠ�ǬO���V[��b� M�H�(֖k�O��=b�`Rr�%*P�QK�ɭ ̋�A��p�T]���'!��@VV�Q��V�Q�k�n�edXvK���%�j���5�(����'"����"ů�@����*�@H�o��V�h��4��j�~,f-y^P[�G~@9㻢�=	�!H�������W0Z��J�-�I�c�/����>��U��Y0�sS�z8�Kd��M/�Og���H+.��	�*���������Q��Z�u� �Q%'�;xė{���C�,��rT���X��prn	����� Hx�Ŧ�0N�*ԮK-ȿ�\Еa8����_�Fm��+<� s����F,I��h�F�쀨^�i~!���� }��1����-��,��U�J�l���'.���T�#B@	�y�&�\�y���|�65��+vL4,���k(E�������K�و������� �Ubm̭�ۈr����oz���$�;ޯ�gO��8��>����4�D����҂���F���X��)�:��[+�c�8�A��o�"&@�%�D����^S<<�oIM_4V�Z�f� ��H%\7O��&�-�;�w��Ud��.�)��8�I��I"���������!W��c�Zn a�52X���>T�%�]���Ҏ�q���՚����o���7��� �,!��1��� t�m���J�c7Uqs��=��i�Gc̓��~�}zh�ppP��d_�Yw�,h%���J|��V�����:
�I�"�=v�q�B�;���=��O��wZ�崉g�M�IhD�"&:�@W�Vi�=�ai����t���qEՎ�I�V���8'a����ǒ�Q\�kㄥ{���~�����ݡXI,�8����F+[��zG�mAz�;��۴�m�s_��`�Xn4�s�P�E��jIA�V��-�s �V�e:�I}U��o� W	k�rtD&�o;/_���A}��vQ]�B���l���Ǔ���#�O*���ij�X�]��i�b���n�g� I����ʕ�1��s#� P�Df�-c�W�C5lXw$iN��q����T���ȕ���,�U�W�B��tA��Nz�|�B뜺��<?�Roi������F19-��Ys�G� �W�4�o�a����A�&�ig��x����+�X23H 0s�߉s2@�W1}����Qi�j���Q� �H~�O�Oc��* R�M�5��T�`��^�'����eN�uC�����o��'����V����~޸Wn�v�� �U�T���#yʗ��fD�����YY���i)�����z���B3(/��'�[g�����&�����ț�3\��;��+W��y:3���$����"� P��1��T�B�ە�KZ�K�;�s�u�{B�c"dg�w�(��63N{Or׉�p��Je%�͵X�މj���w��i-z��wPߜz�.VCC}Iբ?���ƍ㪈PI�V�l��&'�������MQɧ�ř{w��MN.�3^�;��͋������T��vyju���O�
�5����т������졈�*&�m�C~�ͳۤ��-���?�܉w#�G@CY�*<I����"���`N�z�]��?pA��5���VD|$}o��u�S�d������~}ߔ�F��N�#�R,�������=w	��~i�V���y��t�FGl��S̤�oS����4��L�܎���쬤�rM���SSB�����@�@=��K�������z8�P���P���Y��{iW��j���n�w���Ꮂ��Ӏ�v!_�k�z�y+��p�d�I�No�Z�._E<��Q�;��!�2~j��H��8/�Ir[��#�k�q-���Ȅ,�%3�μ� ��Eq�u)'{�|�y\�( �-�f���\��¥�IÄ�TZ�,|$�Λ��F����m�,0$Bbk�$Ǚ�1���5�Aȍ[ۃ���҉����%F��cZ��Ƹ��*7Y�ލ{�6"��$�«����Fc$��������F48sZP�f�:CV0�Ԋ���0p�h��'��B��F<�/�D8�|Ẉ�w��}ߟ"N�_R���nT%�$|m�5?�O�y~R�BJn	��wD�F�N1���ɴn�m^��}���,f�)b��鍍�ܛ!��e{7%SK4_��/��_�yU��(�T�>�[ْ�W���o�/8TE��[z�%��xʃE��xa��)	ޡ]���sr�abV�ï���gl��D$t\��WH��Q����Qa�4�,�d����ӻ���o��s�$c�a�=�˥��=�����}c�v��3I��+��n ����*�,���g�&�H�?��K�����鼯�@��u`���r[�2�E��v��sv�J$��51�j�-T	\��^���9g3���̯̝����Y�k'78W����H��8T�M��zr�|�o��FB����w9�n��g��n�a���V;u3�y���fd�'��a�d`֑.��Ͼax9e�`R���T6�����xÔ��d�Rk?\&���h{���+���]���^�4���艁X9���a�������bWn�-6�ٙ����Q����sc�''�,^6���:7�?zh�kUn�,�����8��}��V�+]�D`�fX7W��P�OY��!n�0A0��ɶ�I�x��T�X?G��6P�[B�n����	lק���\3I7�%�8�z�%4� �wMKI��8�r��&챕N�=H���O���b��r�+9�T�|+�q�̃˘wT�E-�$�ޘ�n��''���Y��x�R?��0�.t��'�^���u�I�HX�,�K}���Z��_��Qת��6�|;=!;<r,!q"A_���E��S-�[�#$#đrA���� e4KC�D���zU&3�f��1����RA<#3�3Z�?�Io�3�:�&(Q{�,^}ە�)|S�n���>0�2尌&�M����Vk�,�,@��`H��	�q��q��!w5�c�)��ӱWJ1��द��֋O�Nd��`����MQ>��5,l�e����3�t�P�A��"ܖv2�
c��ԭX"i�� ���Q��O�#>��A�U$⾙0;ޕÄ`v)⎭���<a�S��>Z`Ӧ��3��4�-����W�c���d���/�Ԍ`LJg�H�����H;c��n<�<潁��6E�Ɯ�:ͱ�Y�B`薠��ܑ�,�x��{�
��S���Α)��gF0`����l]�8"J*��+�ie٨�[�`��֠y�[������}�p�r>*��Ť�=��8\(��Gh1�/�'�f>.�"C�,# �*�̞����,5Ԋ�˯�Œc!b+��e!+��W��Fp%]�>��l���p�)��UAFV2L�{�#(>�	� H��j�/���Sl��g{�RK��W��]NǃU�� �C���<�/*���tz˛�i7�d�	SI�̼CŸ���=���*Ǝ�>Fn#�	��r��'��4	���2L����)���3�1�e�3��!�ٱ�y��<�#-XL�};%�����>�&ǌ���`��$�	]�.�U��;皽J��a��Py8������o�~͡����;vqmRy���"��z0\�c����Ǹ�J5�S[�Ϊ�"L�p��Vco��M��=�>�9��I���6�"��J���
/4B�Pr�=�N\3�j�I�a`�����P��"�����[ %��3� ���\w^���c��2�D�
]���r���������΍=BK�G膔EE'��2�u����I�'��1���gv2?<f9H���,��x�T���sFj: G?��Ie�U�.h��7=՟��Y'L��W}��ϔ4=�~�3 �zk�1/��o�MT�X��<�}�C�8���q�ɼG�|�M�"�};��.3x{�����HE�� V�ż��S4'�]�yE7�����;�c)���?&b��jy�۞��&�����}��*ŏ �\��;*��{�g�v�o�5ԛ�̔�z��kw�@G���@�t,���fN���3U�s͋��^�Z����PS�L.�H7~�*h��J���
	 g�I[�/�9R�C
��(lXu��~�e+E6��>7Q�b����\��r��l��a�"Rn�h�&L�^&LH-��p3@�̷�ĝ��J����Q
��V:-��3�ZC�B��;7A�&P�Q����wd#sn�,���v~O��)'$,���g��9��L�i�Z@��9lxPD��5g�`>��w��{/]/��5�_o�!��#�k���ȁ;ނW1�1�v!�tpz�9ԏA�)��'���A��ƛ����Ϗ��9���W
񰡚n1D@�,��4���Gp�i�p�ݜ|[�9��h�}�����;�KV������H0�Ң���w]/��zG�า�l��!S�]��a0,��i����$6�G�OGܫ�/��{�)[���d��53��;�����zJ>e����Ok��4.���0[��踞C�u�<B1�`��f|&���s�eJi5�r�$������=��\� bWt��̊�����+~*!����ȩ����Z�B����t�A���v�P�ӄRnl�̩���H�=r�ts�X����"���=�<c��ĉ�&ͫ���Q����^��>�J^�Hx*�-�����I �[IMo���aT���ܫ�{9!�K	�ȋ*3��i�*�x�����<�V� �O z=�B:�ݙ���x����s�b*}�,Y͊cX��l���������`���*O.�Z��f��H�F3Q��S7r�H:,{v�I�>�7�lwf7&>[�F;��I��Bkk85,��L`�fN���c���Ky�eu�L��2h�Y�$fj��ތ�lc���t��,�Jx� ����k�"L��������]�]W�Y���x�3K����i=Ґsޕ��g��q{.��n�t���KM�H��7���e���o�e�]��h����葌e���|�MW���@��1lq/ͫ��,�i��>�L��3}�Q�z�8�I{9&R��!k�U�;��������YS�]TK�^W�TΦ&o�=����H�!R��m���B^��\�b�f�;#���F=[Jv/:�c��}�׹��)����S̃ۊ��Hf�v��`s�!H���0�|���#�)a�}.H�`Ѵ��� KΙK��W��E��/є܁�[����K�h%.K�=OvP;���֮�g�4w�W�3*�x>�$�?�4'��RtL቉�@�����_�d�z��}��O���r��v��1�[�0`s����A1�?���*�a�{ղ����'�2 ?�v��nλ�h�]�EMP(�d��dMH��.}Nu��%-� �i+^s�`U�a��e����\s����o�@�O��+��i m�&��^�9��C@��G�bN)2c�$�m��l�D\vq��Q��]��U^��C�곘�K�/���J�!gS�B{�Z�Z��K���1v(yu	�,b���=U5���]�.�O���n��5u��ܩ�U�ŐZ��7�|3@�>�g�%pa���n�
�$!ځ��(2/��%�h��:����ބ���{�DI�s`*�!l+=7v�T۾��A�B���Ic]��]?������)��+�c�&.y�.�����������
�PFPF
W �)����:��3�7bo����YS	6s'���I��\�����8�� �|Z�t>ϛ�.�"�ŋ��1G.���.�ʕȜ+�#=0� K�@Gǘ���{wS�Kw�;+�T�97���^ș�qaN'��^�},�"P���)�=��8Id��˚�e���vT�lnh��(��+��hk˳���qfcz�J	��N�3�:P���86�A��kN�� ���D	�mV���u@/���1���<��$`Se��L, h�����SO𱭭_Nz
�\��N)�eE��Tp�]}:��Wq�(�J@��Ɣ+�#���}�X[��N)D1&4���b\�ն�E��$���e�q�o����>���h�㪑�0��7\Z47��]�/Jg�h"�3n
��U��/V~�{͆P�\#i�i�ב��:�V�lh�w�qm�Q ���Ѭ��S���5R������;/4�yk�&1z�j眄���;�^n�@�O6���=�r5�a��_`M�]<�T����G�@n{�W�3xJt�����?����u��|�� Ĉ�*H��_X�[Us ܗ�2��Mmv~�3�(�{�����)}��/�í{�|h5s��_m�M=��B�9b�Io��w�rx�`*�����F8�qcO(;�^����Q�*�,�U�>(���lP�Eȳ�}�,��^V�D����5��&U�q�q:U���Oo.�di��m�[f)Ӻ���R�4�ү�j�Ǌ�6i��4P��g��\��㭕dX���Z{�	��VW���T��"E��b��i�½��Y0XB}�4-a�<	���6@�(������0N�U�c�,2��C��>�5��7��A}�}�U!�x>e�����e;e5�Q��~�̮��ꗙ� ,K^^���+:y�T�~�1�Ѿ�R}���"�Տ|��j�M�~�o��(8�ze!X7"��LZS�e�p>��7;QL�P5�lK�����ñ�/A]�������67�Z�F��$�>Nph�4�3�1"u�vޭ` wȁ��9���!aVIV��k��S�ɹ �<� �@x?n S�u������Ć�wy����f�j�G��O����\����W߬�|P�n��ن�
��x�g�~SC��I�c�T>Y�g��j���/8)I!@�#�^j�3�׹¤����X>@N��k��(
T��ϡ��?MZ�;*ƶ�}k��;�+B�/����_�o�}-F�P̧S�/(����D��]����L��5=#��Nw��N��32��Í�2}ΰO��r�0>�m�f?�\^�Vf7��	���Td��f�}��V?r��������`mݫ|+	�
�j�:�9h���n�Y��;��Eٌ��]	Z�]�KX�����Ģ��$.��b�mRŭ�e6�Nk� <��3�]37c�:�� \*���q3sq{�I��G�ڛ�jNn��9���&H- �8��O�:��Xn�Œ|rI��]��e� �xZ"DU���y�3��GLN+�r�(`����r��̔zW����-;��	wX\4�%�"'��sR>���t}˰Ն$K�AP_>�U�����B3TΑ�J`�ؾ��Ü,�xd+דX[Xv������7�֥�6k9�B����}R����J�M//H�+�@�	Z_s��	�Ej��������Ag�&��(��MQ��,�������!*1l�b����5|=�lG�|�W@�+����p��4�Z�?��A�������?JS�{�rB��7�b�����2d�Q���I��}�YE�z�b��l���4Q�>?� 7�w�)=�)V��e�/3ۛ�7R���T�+W�F��� �!ޠ)os�lZ��o�tO�aO0�7�b�o$	m�jb�l�7%��uo/Y�}&�����&�t�k��FZWn��"/�'Exz�Sl�܂{���L�z"C��D(X�S�k�e��tcР���J���*;�kۚ.�b���'��]�5���L����s(-$���+X^%U7E�d�Gc����(�6!>"o"��(�7�R�Z��U.�û��9�!��F�>!�:fk,���X ���ӵf����j$Kb;m�AW���t�n������?�Z��Qkco8&E�l�����"��\�x�kn,�!��6H,M+�m[f(�0�#���?��Vǘ�^�i?�Fi&֗ey�O�:����j"5/�y�`�����rz�� rk%�;��ʹtR+�6b�837���ˡ��_��0Q �'Yq�h�o_�v���NV���� �Ƭ���m=����=�S�\��"B=P��/M��/��O�o�|["=Юԏ�����ҭ�km��G@.���m���X�?�Z��7FN=��;�L��*%W�����|QܺG*�����	�ݪ�*y뉍D�l�X�J�%��>H�>H!�/(��je�:��[���� v�K�ԏoWekG�onJ"�V��ߏ\�f��?
��<��� %T�T��-�g�v��׻$������(~ᔔxV���F)F��S�E���<1[.�]�1SC�N��3����|���##�1~��[���
�yH A����U+fq+����i���Z���C����� g�s���O�6up��&�O��ʬ>��0�FG�Q�̪�2�M{Jx�����C+ڇmښ`h�c�q)��]�n�d��-c�k�_��ح�������_d
����?�o=C�Nn$���7|e�>GGn��2%�Zb�Bz�[��A�E��"w�0���4��3j�����v�U�_���y��7����+�Dv���F�i���H-Τ�>��:`��J�r٨��J�Jo����wRq�KKԟlS<
z��	���UN��ڈ�W�����S��y����A{��ۧ ���S�}H����r@ޔ�X�ں�0C,�\��u�ȍ[=xim�d���%���o�"I����&�(��ڭ�.��R@Qu�Jm
�W!G3nYb' ��FE۵rj`�{ ���_�V,+�H�T�]�������x����@�ɱ���}�Է#&^�ZUKc�}�)$k���"���n��皔��>G�-��m�"Kw~�x�7Ο^�����P�7�����ei��W�JoŁGf0O;��m�>��R+߇!��P�<�VJڏp �/sc{����.�@��F���K�416�aӅ�#��eh�!�z��r�n�;��Lm����&fו�Ta|�5��jx��u���m��*ŷ�f��12�<��lv��F�(8O��Y^�?�)'��l����}�q��镆u?`�c&��0~�ʧ���$�?�Q&|����>-
A_[=yj3��(�n��w���{ze�%���K�������y++��CӒX�-@����h����myw';�f'~^�������)�x��ȥS��x��3�{��`n�e&����P�=�eqZt�(Ku�Y�s�9�
ogZݵv�O�iu!��̱��i�I�Z�z�Z���`��S>������,�h�?,�K�B�&t���Q����A8������t��~��W��Qt�3�f�!�֜�ò)#��q��-��U^7a��=�U�_;��A�>H-G M�\�~⮇y.��u�Í(��X�.��C�mqB+�|�/�����ҕlE;^��/�P�.]~V���a'71�+b�!���$��e�K�՘m ��d?�*%�M��Z��@
}�c�M����x��ԁ?t��#�*��S��d��G�_`�5�a��& J��6�(�Xk��`�d�E�"Έ�\��l|��H�EQ>�^"��
W�e"���>+l[���w��4�f"�Ċ=�)��֠�$hT(��P�a˚�)1�DS��3�^[)8X��������fY3�z�-�X#���Q�&��|u���Ռ���Kb�
c���"�N�Y2i
f��oo����TR�P��N�EJ+ZZ�� !]���;  vN��<ߑ^��6���jtYC`�=���9o�8��.���5=H:Y�G�M�j�:�J�PB���d����X�4��s�H�v���U�� �ߟm�+��:Ec�n6>��CAT���JoZ��4��I�MX�2_5���fe��l�7��4�Q��"�	2Be,�Ϸ7W���k,a͝3n@!��]F�U��˽���3����Kpe�/���}K��D��8�U�>#j�J��<��k�2X9��p���.�ȁ;<Ey��Fe|/y�^�� �Q��0ڈ3ѾK%��!��%�2�� Jw9�0�$��]{�{4^�qt��S��x͡QU��E�G�8{I�bX��c#���S���O�P���+�
*���kɡJ~�k�<T��E�����k��q%��<�K�)+U�6���J�[]��þ�ac�	
�
�,��.?��k�DVQqQH��{�5n���e�f��hT�`�����	�����OF�~H嚓�(lA���_Yr�:�a^>���f_Z��ąJ�Gg�M�!%�|LV�|L���٬���� ��ȴ��;������Ug"���׺
�[� ����d,��xTN�-���[B7���v�#�1lV2 Vu�8��$oYqB�b���.36�So2'�`KH~��~f�?�ɻ~B��G�S������n�> ����=tU!���<no�]�eܕ��*�'J�R�i�s�ґ+��Z�����,�����;�$�95,s:x�
��9E0�fu��$�O=���N����KEZ�J��i�vGy���U	Q\'��R5�T�����m�-0��Ǡ���/����䷌2x����6 ���f ��/�g֍*Drg� Α*�;�|��"��4�Y�&���µ��&��$Fn8�E�֔��r�~ �gwDT4qq�Fq<X�G����2�!�yM����IB[f����r=��y-�!ainٻu�Б$�v	�6��0[�^�,�Ȥr�խPUt�]��\q����D�{/9�o�n_�2ù�w7��Q0O�eS��������җX&q����h��xp0h�Z���7�`Ϟ;�8�V����zď��:ɶ�!�IE�Y���]}v�p��F��L���F`�|�6%2Ld�ܩ! ��"U% 逹J��A�j�7�CsHkO���gN�u��j?�c���4����n�\T�����Æ�x�1��s-B>���&�	[=���F[樌R���U/�y���m:���k�k��AT�(4wJ���P��XP�(����ɗc�(���)��S���l�)D]�z@�)bų�UO�Q����jZ+�;3�����#�1L`p
jEmλE��m�Q�������n֊̬�b��O{�X�`,�۲THk?�����B�fk������C´ϵ $���<�Ü̧��q��=�$AM�0�g��t�ό�G���c�th�@�}'ߝ�(��K�{K9�B�ݤ���Q�����w���kKV����ER�,#{E��#�\ ��Z#�Z�2U�T;�
��|���gS��b��	���m�CR'E"��h��-Rb�8v#�G�n�*:	c�|!콇b6 �	���{վ.��U�7�:�����@:�ñ�:�;��.�h������ ������A�~(�%Q�����YMev� b�bש*��d���q*+��̈́��D�٬���II�*�Mx���܃�_Y�{���W��ΘǷV�O�$�޷S{�c�9hB�9�<�[G�SM\�D�=�U�
�1P��CTdeos�3�o#j�k��p#5OZ��;`����M���aU��"�cv#�	5�TТ3��Fq�}!�w�o��"��Ӓ ,�A���1F.-���A�f�����[��� MNv�^w���pd
?oY7�d�[����w%'�:�1R"� wǅ�]��G���b/@'Ǉ$�f���R�!X
C�73�	�¹������'�kK!�(;^y�B��kAU6�Q����ʎʍOL�Y>h�.���%T�V��sy�߆I��̩uX>�Q��mq��R�z:)d��58O��+�F?��IȨ�>�ݳe�Z:��w��T�V¨�qÑ��:������P��z< S)f���}�hs��R�c����]�d�Q%�c�V�*!�<������;F4��fNdՆ��?�ނ�_�/����l�bݹp5S���D��ځC��u�0��fcȷ{�vT�vI�6{X��N'@&
�W��K�^��-�W�H5G?�R&я�)��#VVi	9�ս�HϏ���E�wa���N��E*�,?��RȈ^ZmOFQ�wx�����_	"���S�����	����e��?�aդ@�cQW \�	���ǬnO����0E8���x����tR��Vp#la���U�s��y���yP������c�i����I3��A��'lڳ�yK�dOE����Q�L��#D�5U��C���`�:���B�3���t���NB�{�f||�+�Z|,�5r�';ԑ
L@����+��Z��i��l��S뮵W�����P�XjX�H��8|_�gi��� ���a�}�}��x@�s�c�����i���bBfB��#���{I#GD߷}X��>��U�Rv��1�J���]��9l$J�X�6a�?)n0&cIK��d�
~ ȣ?�V���
���\�-舥��P����]6"�"s�Ş�|ב �W�k��#vu�[���L�qاߗ�4[�|���"5"��R�'�]��A�Z�e2�Y�ڬ3\�����$�Y����m�u�΋_�l����+��#��o>,�XS������S�����p:�B�Ҵ�=�����n�.u��8�w�H�N)�I��7XN[�-�i����B��h��+�\���C�|p�����;ǭ�S`m8��!�����F�0� ������~Gt5�qw^�Z������d�&e0��v4Mۚ��f�������Zc�ʑ��v5|[�h��L=�m�U��J�qt�ٸ�g�����zlE��i0�z���y*m��Â��8�f�N
�"l񝲕�U�9%��2&��g���mױ:)��ʝ_ ¥;�*#@|:�0y�$��d��}��k���AK�=��Cm
�$� ̻�!;������]bMVS"�xܶs*�.�����W��'��i�� ����$�t��i�x"��	c�۽�Ĝȷ��S= czݿ���Z��q�������`��M/f0ނ����9��}���xqu�s����fW�@���6!��P��7�s~vF�4|*O��X�P*%��_m�E~�]V�8α{�0j����-��2�_��E8��ۑ(ޏ5Ʀ!r�HW°�!z���L)h��L_�zͺ{F/�2�)��⯾�d���4�����4�B���ʁlX�	�Mg���X�}��NB��.��*�z䌞�[��˻�ݨ-�k���o7 bC��l#���2s�b�M���a��׉��U�s�$jz�B-���uJ���.�J�A^��*�����9�Q=1�]|�������&ʘ]���BN�^OA��D��X~���u�b=&�a3 ,�d�ё�[�}��#�Èܐ�=����~�zbf)c�T�u'�})�E��)Yhr���ۼ�<�V2M7�{I��3�-�R�H�x`��ǝF�Z�������wXܪ9�A�w��y]b���ݛ6����z*m���Q_�����V��̽�g(~07`�^��ڿ뜅� �#S�B�H�wI���jֲ�MQb�+�Ď2�	��C�^d�
�2%�o�s��p#�j�O_g�ܝD�<�%^3��MD�fo��De|�[{]M��t��ʿ &1Su�щj�x����\N�]v��ö:�	�?n��X]�Õ�Т�o��V�Н�+0C�Om$*��	��:�rFŐ��(�P�\�;�B��L�p��{y��}E�?Vvn�#Q���e8�V�dG4��W��ٲ�_Y��\�©�`?��<2*�$���8��ۜH��=���N��4�c�tb�k^mY�G`�+�@�.m��f�y_�������c�J�%������<>�I$$�s���?���",�Z%���~�h�*D�g��$�ӚIƁ�ҀeV�r��/��?��S&r��|f���5�52;Q��v�"
�P0�~��S�{�_;��+^�Y�^�m(f�-瓢�ģ��rϋ��6����<����͉��/'�����bg@x�n�G�7�ҏ�I;�t�y��1��T��?OP���p��U�Ә��}���>�;�2��Cǎ"B�S��"zc'O���T���z�>JvN�t[���F� 	�u�m�4 Q�x��JXO+�E���\��s���7�R�qRfQS���-��xt��}�ڢ�>#��C�
������V k�v(��,l?�k�@�O�῾�։���
l(9X��X�:1Af^}��5�h���rW��ـ�[�1.�9y5��݋�>�i����4��3�_�4�h��]e�jTx�Rͯw����*g^pτA�%g�j?FR����",�Hv̡n$�g�;s�d� ��yw��{^�.D�/7q놅%땖��Q�*r��)֔I@�w���Y����Μg�f��M����Nz���Z��m`ƴ��D�h�~��=J�NK�T��ע�"�ȑ,�R9��rBȴ5��S]
�n+����a�!V��?
�����K88@�@�"��Y&~�
��gà�Vٴ�5๰'��� �8^������L5p엁�W�JZێ�мV;հ ��69֍Bۑ�5z��C���E�����P��p)9�kjֱ��A��YQ�� |���\P�b$c����T����2>u�*��Y�k���W�q3�/�"K�޿��S��O�Q
'Ɲ���%��R�ʛ��$�����g$?z�*`Vx>.�Vi���[ϼ���	��cM���0��FL'zYR3�Y(B|e��K9B��;�����H����X[,9��?�ü�r�x�+��~W������֕L|*�4Nр"�|�LqkR����{���A{��Fo��'6xw`�&��J#D�t|a���G^��#㤱��|���J�,��(�:÷�Ǳj�Uy
��=¬h��h���֤�ͫJ���1I����Ҁ����Bܸ��R�b����f��u��BWV����zj��P�r�=����=�XϕeL-��!Y����<U����R�￫Pmv��[o��a�'��"v\����P��
mC-��Ox��O`��<,뢑ՕF�:K��O�^Pw��X���w,��zEHc�u�G��ў���<��ϒu\�x�D�ڧ��Z�<��7�	�QL�C�Ɗ����*�y���N&�h�a�����u�B�n�2�n.���c<�v��A�{�@�I��r�v��ׁ���	Q[Ѓ����s�]���r���E���1</�
D��H�����9�6bU��')��R��4q�4�,� �f��`?�Ϊq[��� �$����fQ>���|�c��;Չ�AO���n�+����2-]�$��v���K >J5(��^�J��
fj��O����]��T�D)ڛ�+��}M�j�ZD�����G�����g�es��7��d��@g��N	h���3�߾]���.C�#]:�к���pǘ�N��؞�6Q�1���YW�ղ��?�"�}��M�J�{.#�Ă|�n@X��1�gE�_�b� �;8�&�_�m�y������b�?ų�S��/�k�����=��<ᾫ�e�cJAb�wS�n�<�'�ɒ8�gμ2Ox[O
�DSݫ�D�������cٶ߁-l��54�/W]5����넝�T���n��Sϛ`K`�|�a1�6?9X)H�v�%�%�
�Ɍ7�zE:eYwKFc�$7J��eB��d=��VmE�����Bؔ��i<��O�dv�[��� �qv���z�d��كȟ���Q{[����.W:���-9�TM*���A�pD�/.���$E`Rd<�y�g^��۟-��i����>	ǲ�y��U�_c �����_o;����Ԃ�~M>�	
�ߥzA8���Hb>���i��"q�1�?O�~?'ㄠ9$L];&S�1� �^�xW�0��qC�g���v�$�rW�Q}5/�A%�um��{�sE�M�z*Gy����=pMk	�:�U9Qh
�Gc�N0+�\���N����[���a �M�~	���T�Hn�Nl�
:Nj��_į�P6B:�#���ǳ���{��p�>!�,��̃�o�:��d>Y^��Z���@�v��-8�%E����p����1�z�%3��e(Z��Ѥ�Q�����Y���$���v&���2 \q$�g�|���9�8V�vp�����Kc�{3��� ,,^�cd�$��v`�}��W����-��b��YP��sa��at�f��������V�L b���7�7���[B�ŉ[�ű��z\t�
�T,��g��e��7Ԡ�٦
��]�Pn��^��{�^���י��Q�+�)S�:��Nh�ξy�W���-�H�6��Q-4YzOG�·գ����B]'5"�nO.���Hr;�ln � �w����o�����w|_Ɯ���&$7���S��HCV����(1�E. ?G3��h�9Bt� �=���NV=u��c\~yׂ�/���.h��]��\7�M04��wd>V�u�GA����q7��h�d��J|nA�!���'�м�~:
p�Ռ��� �e�������U�o��*pP��~��o���A"/�(C0,�aA:���
ǵ�5����)A)�2WE����+R-��w%�p�P�W�`�M�Q8솾�e�~�}��Si'2ҽ�t�#��ZK���'"�9�Z^<J�5T�@����Y!��`�&%n��nAfN�[c"ɖ#��*- ����J&|g�f�Ҽj�6���7b�o�PԻz��ld�&t�]���$�IX2��Hd�]1Wk�Ɉ�6�-��XC
pR_���T�N�yz/#�q���n�}�	qF��0.L�gW�9�ɷ�O@����e(e�F�+nyx�w�g����w�w����wt�$�+�J y� E�dղ�k��J@]k�J��ǩ�	]e��<5(_ʋ�8x�=Ѫ�L�ĉT!���
QPP��-}��D�=>�5�p�.;��Y���4o�U��-�I����f��`�yJ����G�Lz	����F��Z���`Ȅm�#���
>����]&�D�XU*�3X�v��h��jCWc��$D����{��	�cb���D)�������p�?�h�_��]zCy��j���U�3�ǝ�k��� fu
4g�tR��$w}��t��[�8cu+y�����F�F�Lġ�KC�3�][���f`�N�$��G�S"6V
�h>�_�`m��Ņ]X&�4y�#���-��
=��ݪ��:�g���H~�8�\=D��t~�׎����Q�@���;�!B��D«����Gh���B��T0y���Ox�o޵��:V�yH�Sm���-��tC��?Q`��������q��"��=Fm��)��gu����W�$o��KG58�X�*DK-�Qep��;c�j���9��nU߃���Lz?�2�[Ŗ�/��^z�&d�JA�M�'W����@t�H�V�hä�m�9 �`T�9�M�i��
�g�!A�������S2�T�)#�����CP�����r���ca�T����u��N� ��=���MѾ��F,A��2��%g���M.XD뽆nTpĜW�E9l��v/ox��(�@�;���v����}��I�+�������|�h��88z���$�nx�[F���A[F �G$�T�{�g5R�T���_���c������{���4����X�4����N,%1cf��a k"��)p�(q/{9�v������S>�/��
m���/�|	���@ɋρ���+L��zN��t}�G�Ư}LG���������c�`]�ѧ�S�����P�6���U�Y�R���8����������\/m����ʚ���G��~�>$&�&3Ճ<�[������BH��@a�+�מ+��	�Z�9c}��H�6����3U ��JG;�E�R���̩I���oLi(.�I7�ܫ�lW��`�vi��O\2q�jR�"o�l��z��b���L����=��:��ŦLЧ�v>3��V��L�C�ꋬ����BNG*�өy��F���e{�\�M��\�o�c����	�+ӏ�}����u䤺���t�� ��/^Q��o`��֮�x~�q[D�4CT5ny�.�I^�m��PaFZQP�lmH�lϛ_��hХ̧Dj\TS�ٳ��j��D6�����	�F��V��Wg\#��	��öj�c��N�r%)�6k���7�L�]��}�}�q�մ�"*�`T���ÿ�F�h�ס�a���7	�ae
�
�:�-1�s�!!U�9��<��3�RB4�sC�b��ڐ�E���֌�񉶶g�G^;��&��h�Ll���4Y/]��2�'��6cG6��)kҘ��ߣv4�� ���F_;�޵M�>�R���imۛT�i�K����Df�1�2Ů�oi~p���[�K�dXGq����cf�L���ة��G�1D��F�3^�R_�:�^c)I$%��O��g�a+�CJwV�c�C��b)7��wj3���-�#k��I�P��B(W��Q����$�S��NsBt�odd�B��T�5��7��_�ᜯQ��Y8�ZƗ�X�X*���D_�F<ɥ�O��wgFP*J��Q�Tt��o ��z��]Jz3q>IA�>X��Ѯ�%0�PX��E;��!��)�a[`;���tc�M���"ԟXt������6��̖��_�&Q��:fP�����~�����Lht��Ix�5d�\�QEG�e��M�^%VMR�������?=e%	Y*�*&3Zp�ãx�Gv ��w�ؙۥ��Bk�w!��C�Ը���m�G9O垎��%,i���(�� &6�`�j"h�	��A�k��t�:�	�[�w��y����2gR�DG�qMl�+W�#�
;2OR:�7�o��6�Z��s2��HV��Dji�:w�~����e][�[�ԲV&��B����@}k�O���F����Ao(ӤիG�A<֥Om��vY�`A$z����8�yw̩�U���,k<����M��z�,�N1�h#���5�D��1��sBT�3�;7���0hۊ�ܵ�[��x��A]E�x��$ z*.(F�g����'a,�fL�x	�`F��� S:w(.��f���kv�AM�1)�J3�s���;6#5������?��lҽ�
X��a�ͦYr�1�gM_s��Q�?[a��� 0����f{���86�N��Z[hH�Tw�H[�>�*ɬ>�$ݙ�%pĀs��BR��:R����I�"��Lu6�v[#SKu]�lU>�v��' ]^�҂���[Y47�Ч=��E���,p19��2Ӝ��A:Q,dk�f6X>��n�~�����Q+�1�������x~!&��έV�k��x�� %q���!7z���+�M�S�+.�WY���'�D�P,�T]��[��3't���c��J�����e��CQxW	�M���4w����Ѵ��&�I��T�Wso�'&l��ʝ���� ����62.�z���b��ܮV��q/#`�&�@ľV�=�D�)Tů�dU�l��}��E:��6��%��7�V�:l���u�pd�Ȇo��Y`��h[ͨ����n��S����~�c�`F�:���5��`�>�2�a�,bc]���2��t;��>>��G�c,�Q)m��@��nܛ�q��=������� ���G��I�$��3�&��o�G�}�zV���Q\P )N�vt��ב�U�Ȩ�I�dXk�{B��-���:(0���Ә��>�N	$m�%Ft�ޒ�&EC�k�]T����j3r��ݺ��\�v`9c����}4��#�B���g�K5�����
��l�7↨7|!����#f��y��xژ��~���}��q���0��@�W�.����R0�����s�@�x�@�~&:��r�ql��u�K�_��6��'P�|�w���_T�B�X��|�(ة�Eф?�R���:� �?�t�T	1���p<��0%�or�_�&��X�����"����/O�_�Q��x��0$6m����ـ������ڳj1�JK����4��&S�x�J$xΑ�i(��M��8:����(B�V9J��_�k�rŐW+!i4�mMW�z���ذ�?��"Q���b�������p[�I~aZ�b��߉��z�)���-��z�Vh8����ji�\�#R_R9]GMy�xĺF��+$�9�Y�С���D-M>�z�8yV�|AW/K�	g DN��Qc%X�s��9iQ�h��KI����M���)a��3����q}���N�x���e뉃y�p8^��]��o�����>'�۲x�k��ܦ�.��QOLInP};(����EF�v/I?̾9�I�%d��㿟�F�ЫOg��%���UT#����o��9q���[S�w؊���B�ssD�I��GF�a:uҵ5bV�2�I������3I5���_�{亸��� 򬶠z�>�v��n��
f��M�R���gj��`cbH�H�,z�"�7C��lO����%W�ӊ�j�["���et�����-ʻ��W\�;8h��OLU��^����!��+T��a���f�l !�]4ԉ�����HC]`����-z��(`��V�������x9�{!�]�h��;��ljk�Ɩr���aYZU�Y=����@krm�n��=�n��$�6��L��T�����*J�{�KxkULM``�2��i�� y�P8�~������d��JI���0Gʏe1U(�m�+�۰!Ͻ����Bl�6������g��8��*�n��7e"r�".V���7)��
h��t�9�b�y�Ga���`d`Y.:�CvN2�x��)���l;K���Z<+m!��o�Q�o����zQ���ҶY�t��Z�1�/9>Ĉ�=�[;� ��mR�q��Y���_�۰&�A`����P��x׼���~>軛�.�o}�F�� Q���֟�UN{��[�=��ͬB^7�����K�Z��$H/��b����pDN�sۊR�^&c�H��|�������&��0���L��hDN��V�.g.�P�Zz�UK��=0�����3��*x�c�N"��}�����,�r;y�B��}��EDGjh.�y��K���k90�Pb�`��1�mLm�g�޹��:|M)����T ��E_�� �����>H9[1���Q��D|/�p��ݑ�/;��T(��Oe�y��»�,���RSȂ`1H8�^��3������Z[���8�D�'Yk(ݷ-�����иg�˘ͱ��
�)���(;���ޱ�����&�%uY�2��
�{�d^�Ѫ�Y���rQ�{@�9@okq3�'���ݜ�����a�Ջ���H����x'�� ���&I)��Ԁ�o�BY�*�ʚ�w��!���]	4;�o�,�*ċ�	������`���=B���T��]��b3m�T�~�н	0v~^IET���+��ӈJ�D\(�6n�Z�l�`�ɰ�Q��6�*ڔ몏�]�)� �zÐ��}��h�yO��	��w70��y�^"���o�iq-�gd��
�ԏ��Y:�^7�:�M�0R�l"�u�lщaq�G�Mq�-���fO�����ؼ�a�v��pq�~e Q��r_�1zI����nCm"o�e;|��(�(>=���p���<����|!��(���⸾؊��g�z�o�>Qβ�q)F;S��<Pu�a�l�Q�N��?z�R��>Q|���P*:��Q%l�������������c���T��A��ɜ�3|(��?���hWr�l�U�UƎ���a~�}-����nP�1�ވ횸�͎P3�DOo�ϊT��q�Z�)&�?l}��%�����ٖ���&X����5�r����"KbU��>�`!S���5�����6�$c�&1uv�ݒB&EtZ�:ct�xc���Q�l�~�&��R�*�Q����2S����]��h��G����]|��uI��χ/8�`��U�y��,u��`�����?+1�ފ[X&v�� �T$��	Lϰ�["�W���l�P�J�����7\�y�#�%YA��B�'�"Z�Ȣ_!�M��Cj���uջ����L��n�[6YS��e>{R*�B�\ uFs��*�[�xP8$���!�����^Շw�JJJ��{D��h=���|pΨ�S)�q��4<���Y��TcjP����?�lx�� . -s6V�Ñ�.�o�.�U��<�;�oh�Ps���_p�Z	�|������b�s;�2�Q����0��)�x}�t��	|9�HfRr��BUA¨���P�{rs��S�U�����h`�Xo�6���2��"k�p�<Qe2����%�g1
���~����ȷ/�Z�Ӹ�		:!�k(5����１L�ҵ�,��h4p���$�Py���fy��f03M\���7т�l�-bIc�Q/Y�Z4we��>�p�/�r��G�l���i����	\m���4!_�L)Ė�:��*r� 5l�\}�<��VZ���ߎED' �{�{�u	h&��~2V
�a-|߱�D����?t���:O����c��N=��x�r*�,��n��l�Z������4C�r�ȋ��?K$�@@�`@I���u�fi�V�U��|�;,#o�w#ˆ҆Sʋ�3H��;�������u��s)g(ѳ���2�Y�E�򡕋P��yё�A��ĩ?H8�[��D��zզ:r�c�M�=�R"*e"7�����d3�֠�K�OS*�4�I��6�E=:}�B���H?R��T��Q1�ߍ�F��&���N���á<�0�0�0����s8��9���f�M�&�.�V�6��"�2�3��[���<�8���$�&�~�75�mʾ��r�f!E�RuK�����2���a�δ�-K�>S��=���7�ܓ!Ï�q�X��ᆓ9�0��}�^G�?�i�	����r�}�ֱDu�2`���k#��3Lڝ�Θ/�r�+� �l���J(@��{z�X����We��'3��/6��O�WJX��4���nv@�瞈#Q2��N����x�*u�<R�\{D��ǭ k�S5rh��m�szf�D}E���$�*������~EJ���f�LF�S����W�(��Xh ��?��	}�Hr���!���t][�L� 0	�I�f�W��îV��,"&��Jո�1�=0N�G�v�^.������[�#�>J��u�	� ��I�������~:��h�C*�%�lq>gyE��|���h�](	î)g��F6SB�ۧ��@�`�m,@�=,+Il#���E��hI���<�d�d��Lo�Z�R�s��VR�H�R$*��Y�/Q�a��L���2J�@B��9����?0k�X��s�_sn��RS����6AJYm]m���e��aߖ�_C�2�@0�ŝt�_��zc#�4!��\��'��'��F���U��C�0����� �hQ�sN�y�Wj�XS�t�3#8�8��f��8��D߁b�$��v��n�뎝"�A�Ȟ�Bm�inbZ 	���F�*3*q}S�&jD(\d�N���c�	P��5�;��oP\���3�"\w�_u�;RբȦ��G�03��e�� ��N��8�{�h��ЖAE��5�h h��>j���H��Of�D��ʿ����"��X%���2�E���W=$Z�!-��Dף���}���|<vR��q�kR�6N�MzQ�/k���ex%�َ��*V�:'��zV�j�ӌqhc�������=9�o�p)8�Q2t6dc�6�mc��8�+@c}�R`�?�Ld�������S���R4]P��WԻ����c9-�P�?�ԐJ@�ȅM�h�_�Mca��,9�n!4b���n�0�C/�H?L��%�COЕQ���%K�G�-�x63'�?���HЌ<�E��"3����xs[���N��A�0�<j5������Ʃ.-�(�Uh�%���*�%X�v?GÊP��'/w�G����!�67^�h�^�	��&&b�6�,Ph"@m�=��LOfR��փ�X��\.c�N�y��G��B�"R��3��~��|:Ͼ:�?#K��W�ק�yp�s���������[�(ꑭ ����R'�����_�J�(�#[w7e��j*�w�����B�Y�����͎����\�5�i�?Q�Mr=tu1���o ���cP�M����%�?�h"a�S	U���`�EA��ͭ"9��4�BA1=�s2F�P��\�[*�HÖ�6~lΟf_ɠ�Z6� �����{/"���Q�6�g�����.h�X�l�z0L̅�ӣ:. 3�P��ܗz]sk�n�u�Az��H�Iā��̧��@,�Ř������3؅F#�$�BhGm�5S�DYW$ *�;$5��Lɞ8�}��Q��E�ޟ��bK���V�>d�ئ�2ALtVK��D:�s.a��ľ��JN^z��s�$"]W�Nh�5��s!�-�F�Rٿ�k�1�������SNBq��ڒZ�����¬G����� �M�Je�QN#	�`H�BZY� �{=T<Iб"4b��fIu�lc�֥=u����q���L���5������f�I}�g�9ԭy^���V,C˵�y<��s�ix�=\��+%;?Q6s��Lizxi�M�'��S�f˺��n�����@��H�f%4���+���tCs�����a���R@��F����ʣ�+nVjd$�.�4��o���D���u=�V0@�iA�'�n<*^X�I����2���Y�ǅ���P%�ho��{��1�`g���Hi����#����+)�ɏ2E��� �_��tӨ?�{y姠�|۱�Q�	��n�Ӎ�
#�s����m~X��ak�6v��<(�!�Ī�Eֵ�SX�_�L<�P��*��*�
N���{�!��a���2Q����Ϝ�{��������m�w]#��#_���C�#�L�9d�����j�����4�Ǒ8��H�8@쇣�+T�����G�7�j�0�����DF�I�]���פ�eq�J��ގ��/'�\$iN��)U�%E�1� .����֧�I�O�i�L��$Tb>������
�K=ʳcv^���@��T�s�p������x8Ν`9Q4̍��4a��L�2�!�U���,��v��1*�`�b(�
���Pcv�J 8��p�@��/#�bŭEtVe�]p���7Y��ff���Gg�b�G�6�SNg�X��6G�8������:.�i��2J���]������n.R2�~1xɼ�d)�>�����H�E��dI�3�p���ɹb��$8��إ�ǗW~,�!��TRo���#4���hֱ~
��!��{4�jn���V�ꆇޡkl!�2�J�E�Q�?�PDyZ�+�'a��_�kV�Ws���EO�$� ��& F҅#b˶=��ֲ;n!F�C���M��~f���%=m�h=u��b�1I�Ru�!�&�ĉd�����(�i�Q��O��yƝ��OVH����
����!4u�0ea��~�A�2���f�>��_=�Wvp�lDH@�Hу+q�1�u�`>D�9A(��SJ,�}<��"2�Yiv�it`C������x<
'��] �X�������
��=F�����j.9�27�c}�Pp��-p�t�k�l�UL��無���e��$�4��}f��
���g�UevD�WP�2K\uF��y3n &E��pf�L��]��� �{�J㇁6�1yB��9N�F>[X�T������I��. 2K��.��^d8�Sv�mn8i��aF���K��Q,k)k���WO�Bx�R�_�aT���Z���!_��r՘��;W܂u��+�ʶ>3K��>G�F$�=����D�3��3�K����<�Yv�-��gd�
qj��� +��H��kwY��:�U��X��hM�����ܙ���y_Nc�yS9��|�,�5�?�='��T�oQ|���L���P�:^�i�����g0:8f��������r%R���v�s�=��]�ǆ;�O�F��q�
߼�z��-�S��� d��V57!�lV�ʟ̕lsu��]!�?�����˫��$��lc/zϾ� ݅#=Z>�f�\8��N���o�����#�\�s�^�=�����)p��v� �@/�V`�$A�p���U�)�Jw��Mb|i{���� E�-�J��ୱ�NBR��ѿݺ�p�[\Q]Tc��K*	�'��Y�x�q�l�ޠ�4��1PS��1J?�2��b��Ǳo�*s(�^�$lv��Af��2�a�EuN�<�_����<���_$ۅ̀����^���j~����y�L��3G��p�aʑ5y�eW|Sxt�U١�!xz���Q���T[�O��I�3U��[��f�=Cw�/WZ���c���۬��������K��iS��j#T~To{s���`F���5a����ך('�ҥ��!�	s8xr�%}�'���~A*x=>��	�@Qfʏh5�{����V��F�2g�I��p����'��� 
��" /m�v� =Dt�D�����6+aG���$�߫��5�6��>Yw��?�O6��[N[P�1&
�.!�|�n���=�h��݁,�G��cz0]saV~Gt����+�O�(o���RU��RI��,�|��9�|2u@��X�o���i�T�p*�m�@V��7�i��@��DF��X��ЅyP���ppUq�S��+Z�D��ӌ!7�>�#�s��c�8��t�ǗA���A
�a�:���?�(�3"�]�N�
���$thK�eV�/0�h�0j:�-�S'޲����.���p�$�1�����=�B��J�QN��E�;����n����(�s�N�l� DHoC��X7P�\U�o��:Q��`�+-m/�5f�|c��W�?�D{ܼW�;���56�����0l��"L�|����y��I�D��|�4�&kh�SJ7y0W#z�5��r� w~��[��pT�����Y-�<��f�ﵭ+ ��
�T�;��*l�!Mo��������؋�#�ukҬ�I���mW���Rw�ꬑ�i��6;�)�8p~Jj�َ��u�����Y���U;�F�w0kj-��s��_�g�(kAύnB{S��V[~"�B�\c^<]�Τ&,fȯ �B�v�c��r]��&��?��r�:,�Jũ3>3dH�+^�#?���;��-��|�P�:��t�	C���!������K^IA�>���ƥ��ꏡ�od^4�GlƋ"�͊���۵8ΝZ�YeB�����M!����(����>��9a��@Њ}���C)l�g�ᬞU����^�o�!�ۆ{Zh�҄��m�����`�}�y�n�=WN�cl�W�3�ݛ�6�A����5@��X
�7��յ��By�������/ᄗ
�xN]�p3��ϹV\&�$�����I��>Y���Ha�%Q��\nd�p��pM��.{��c�'D�*�	mN�9rbh��~�~��!F�(�����1́澠_�H��2��A��E��9�S���h>6�'�H}�y(D۬���i"al�H�Mm��Ja��5�=�'m�8/�e�0��N8�,��<M��D|�֬W}')>b��@i;�vr-V+h�Qk?E��:nY��p�7�`��i����ƫ��ۿ�����Ul7l�h@Yڰ��y?�ڴ�0�0a*�o��5D2����X��߭TQ׊�[]�h����R�����%8�Z�e�N�;5�G���?�tέ����fM\֡��2w�[Q�]�(a���~5�p-V�#�<mé|Ȟ� �P&7���̷A�;���]�j�O˺�h���Uph|�6i?S'�Is�p��d�MY����T��}rL�1���$0>�����HO�@��.�B�|n������?2x��ڕ�E\ �:�Wi��~Pd�w�}� ���G4��۸M�Q��r?t����B�=.'�$"?H�;6:2�^�%�u�C|�4t�E��o8&e-��n����^�_����]}ҳ�%?S���Ln��C��[�Ҹ�Eq^� 1��%�u0�1�C�:Q���+���Q������";k��
�p_3m[Y/�l�3T�X���9�k`T�MP�(�"g0��發m��������_��>�Y0j�a�U����L�����#;��c��8�tfkgog��I+q٥8�S��%v�ts����We}_2?ψMd��Az�EbZg���6�,�e|�w�6���
���?K�4QHK������P�К�o"$m(?�t&}�<�e��S�Hv�/dEm��0����un�`f�?��<ʗ�P�,?g�9͟���婔���RY�R��M�^JZ,�S���03��!T�����`�y�b1/O��09}!�_5����Gؘ7�2�1A�"��S.B`N<?i���ԪC28_�`�����ϖ���������n<l�g��0�#����Jx�N�%Wt'T�0T��V�Ճ�]D�IV�� H�)���9_�7)��h��� =���k��3�������&.�U{Tݒ�~���ه:�#A���|Z��n�����P�0�����J�F\������j�S�� N'�Ia�"�3��a�Y&4ҽ��bz��cK>Ox6�@�i��u�Vzy��@�2�������� ��$��8�6}��3l��-��+�X�hb
�"���I�R�>wi]�ͬ�������8�F�w�%�b�vM�@����>	&4n�XN�0_�Y~%ⴈ�e�8��fRO�����[��0�9y��Ɏc�f�m5��V/ߐ��U�(�`���K����SH�e�k��[FO��Tm�f��{<y������Å�i�������H_��4"`���K��JӀN��3��cO^2��^��ŷB�É�cX����|9U"��0��4+�� � �ņu�B:>�Mw>\A)�.ƹ��TF�[�Ľ�4��2�L���Ӿ�	����HP�vR�@5!�bYo�/�vs�Ϳ�%��m,������*��H�YG%N����)ڦr���O�\Ϝks{x��w驺(��~�H�Z��J��Nr
��M�A2#��5T�'0\�����O��2���@���`�1�9��{y�u݋�[�o��{Rr��D\�b��O�ۚ Ԅ�ڎ,��
 T�����������3�A�"ؘ`6��5[�70��S�*� ��ƔV�"�;���o���F��i��=���P�@��H9)�EZC�c�PQ�����l��,�.���;S�O.��y��(�pΩJ��M#� Y�S2�#�Mi0
/Z}W�M{5��!'t�N�a:���|%
���;寧�iC��;����KE�RU���;�n ��ә޵�
/�g�����io��N���&:��g��W8����PI��ݶp+@*\T�i��L�Y!x���aW���%M.��fRďY�����B�z@e���@�;*�3�6(��t����	�7�o5O��&�nT��vY?B��f�Y"� ��(�?�Ky:�P��t\Ę�e��7؏�4LU���Y^'��3��uc�H����W�N�gƯ����InGZ�s��)�v<K�ذɯ���;��{�3'Xa[��4's?N�"ra�!=����O��g�������U����˩���A��/�o��s���;L�,��٫��"�x�KL�kn�α]�r��?.f���e�̄1Hr7RRR�F~�Je��"+��s]���lxެ�\V�����f��:nCĄ�O[_���<Pgn#�n9�M���{�/�m�gז[�_�x��4�9�i*�+��)�;s����hݍB�0�E���nBv����"����������=���C$����X��d�N�(�ꋤ�cr◸L�<pZ�[�6��%Ad;	g�|ӈ!���>�2M�c���:�l�B��[��x�r�ք� ��*,Bi$�d�΃1������x�֯R%�?)^;1Tk�u�%K ڊKu]���s�	����ڙ�ڴ�b%-���í�,}yYg���צI��6́c��ׁz6W����*�FQ�OebZ]��&���kUU�i���t�o�� U�=���q�b�z(���O��k����Hl5ɬwlh��)2�C�l���V����3�mS�[B:������=f�`f]\K����L�7���Ԩ�C�%����$rtC�?��z�A\�+��5_�u� ��16�Wa'�>�x�t`M�:�ݖ���u��Yl��7uP1�"�3B���5UC��WQt��ϙ%u��d�y�T�xܐ����8,��p��ȵ�*h�g`_�Y�Qe��?�n@����đ'��~�q ��R�@��a��ʨ1|c����;�]5j��,�vN_�a����t$��@���ֱ��?���3�nO��Fg>��8�H�f�Y��c	��r�c�"
RԊ��8�_NC��	;w��Ե���:)��^T��&Gvv�\�Ӓk�zȊgtDe�w����m�S6��mN)(Ya��͙��n��@u���V�������Υ[�f���+��cM5�h��ry���ѶR�%��C���<FzF��F�&���[\�E�x���P�6��0��v��JI�4�)��Z�A�� ��uDUU�J�I�Mtj��{�6Qn�#b��ͅvv�y+x�.�j��p��78��Ҥ!>@0^�Һ["��Z�`*e̊6�;��)�A���a���T�7����������)�I��?��.T���88�op�rk~��/����b��;�i���۽�No�y�8}�BS�_��	� m��)=�)�����	��rJ4�,3N+ r{�̮��|E wW�0��z����WH;{\�ڈ�QV4��� �%�k��c�)���P�fw��#��j�2�b(�C%��s��J��p7��@���gy�#Gm���� KS9�S6�N�!������y�ʴ)3ϟ�V�0�TTp�?�V��O�%-�vY�N�����g�jY�3����<'�O��ұ���z�Ь*Ts���ޜܭ,6}Wآ#�/��	��!v�)�U:Ԅ�K=�l�a%o9s�_Jɝ����l7���a���e���P�����vd�}-���\�r�PZ鞕�.�T��/X����A�D�*��#&� b�܍���P���y����7�͜]E�7c��|�MXt� u��3�����Ԥ����<���
N��+�Ȭ��g�D�dU~ApAd�����cl��T��%�4����=`���yλR#�Ω|Z�hTyܦl^�
)^�3V��`���m�z ��M���L?���6�n���/�r.�6�Y��"ńhm�<�����;eN?C��w�r'��+��r��[�O��<��$Kbu�^n�����OT��z�<T�!��J	�HY�ײ��5\Y%;vC��?YW½U��5��ֳ��N�́�OQl�vN\!���u��z�[n�@�����j�sf�m��"��m��ZH��q���ߣN-��e��
��2-��*�;��RZs�ω�g.��z�r��. ���ף��0�oSF�k�	!x���ް.;�ň�����~ɾL�+��Y6���+~������y�����Tå�#T]a �͹l_���>�f�f0b���Ȳ�1sG�q�߅w��a�zy�<���ܢT�����v>^X�����UN�^��%:+����S��6�i�}���V��$g����^��Ǯ+Mn��|��G/���cs�T���&i��=%s
\�v�8�A��xN�yu�r�N��{�}�[!���M�`킟�!�9]��h�K+ZrU��=M�U[�iί]��@�-s�4�Z��
�k5X�:�8&PfL�*�'uĊ̫��-UTG�G�x�i�ju2�_Z����\1��:���c�\�*x)��(���*��ZLw��
����OL��@��r.}Vg`Pq�~�>�]`�G�[�ҭ�X�b�H������X�/���9oJ�l�B\q9u��ɤth�q��q"Cw48syy~)�@�5B���s�a�u��0:���G�{��A�����>:E̽g)=ZjY}p��/�E`/&�����D�>2�
w��K�$���(�$p/���V����V� �A7�4ˎ��Q�TB]8�Ỳ/�_��X\ChMFም~�o���-�g�`�����y��q
#��z��N�q���{Ac�D" :k�ʝi[�R$pB8|(��V�D�#.U�4�Fm�\�r�#+��K�Ts�����U(�wjB��5����;D�
�P:02�j��+G���tk��
�&��T f��������D�� ���K�9�\B�1�J��J�Q��y��_�9�
�jj�|�!W��4"z�S��ᚙ�S4G��X�w�z�
[�d���P���Qv/��3�`b��L�@Y����~��Z�	�j`������ K�8g8<�Ӆ� S%cf�
��+��9`���V����<��#bط��i�[�d�\�����������ej�Bv���	�}Z�==�CW���]5T�s��	pר��ke��P9~�c=�[�*k��r��&�"���%�vNE#�j6�r�����쿵K+�y�.�;�?}A^ ��� G8�ȧћ�@�% �{��н;Z��K������R֟b�Ԕy�5�.�f5���h���.a����v
�݄s��(��'.�\b�����~H��iVϗXL.���=�s�����B򃷝����RH�Q����u��P�,
��셝�����)k��d]τ��,����b;�\=s9��ǧ���=��>^���co��$���m���#����66R@�&���5��Zg��� ��~;C�ܦܧ7*�=���Lm1�z��@���L����W���9�$Gs��MA��s�V�E�A��2NP�����T�)����l�R�2��	��b���I�Ff�I4(5���*����@�Q�3^3-1p�
���Z��/�]z���@��kfbɎ]�s���" m�=0N�/����� ���V����@�)?�tj�_'��٣�ÙV�7�p�˅,{�1�w�ߩ�]�2�1��X�nV-�IPb���m|��K,�l;���T��bR/�3
�5+ڛ�t3.��F�4��V>��VK�{��#�����o�:��#������ʚ�B�u���9j�6?�1��Fv�k������<��
�Ⱥ
&�}��O]�+����h\�9�K��N�}��M�j�G�E�F������&P�Cü~���(|�^�`�er�Ҧ�J���t�4�T���-�R���'H���QvG�����i���#����e�r^��^j# �i�'�qc:NE2���U=��3�יmS-���Ө�eo*���շ�`Sg~����}��]悍ϗ�/ĳ��
�j�=UI��"��8>�{� w�{��c[�F_!��VK'i�fۈʦ�w��¼��|)㴛h��۱���wđ�:�� VVF�I��)NdJ��W��{$��q�j$9S����ǧ�Բg{����3�0�+)����/�1�2Ed���̉�nH�<� ��=W`Ｂ�\��-j�U�vC��R��븲Z���mĞk���-\K(o��*���ؘ�U~�����㎞F3�2�t�v�\��fM��c8*��j�,��)5Cu�F����g3 O�yч��X����,�6��g�y� ���_�H�R/_K*�2{��
1Ve�w*�@���T�Df��,��-� ��8�����!�]ah��L�\)�}�(J�|58���$�"��l���q�TT�:l�������4�b�%�y�Ԓl�YH{C�lQ��׸k��[T!��OW�Ϭ��2y�?Dy�� �/a�E�&�����������c�5S��C~�:��_�U*��__��?O_��A�s��7B�u��E�Y�iA��ͼ`\�wQ�d���hCq+9��qa�_�.G���y�#[ޒF�h�-����a��[���]��֊7���y��މɀL��bR��bŷW������)���Sx��c�ZQ����͙�j���h�<�d%�^A-�]�7��'������{�L[*�~6�`��dbk��/Κng���_BхM�r��E��I-�I��<P���{,Z�0^,=��h�o�n���b���J�&`0����}��(���K#ק��UT����;�E������D�E>���k�#��}���A|�v)���@gA��1!�L��Y�IB�̾;�j������Γ��O��4!�b�^���ǺϺwj�R��I�R��=����<�qinԠ.˯��	�!�P||����!�8@��x���l���u�?�ǵY�-D縁��؉�*[k2}�\����67�����߄��N���5��9,֥����ѹk��~��ʛ�r+�}���*J�z������8O�ev��E��_��>ag�V��ɐZz�|���5+��U�����XMb�{)��#�� �긤�8yqF6RƏ�,�o2gpJۤ��˦YQ���)����d�r?1��ir�bh�>��T��Id�8O	$l󰆂���Z`;Cr�'E��ө�6	���L�q�ُ�K��:��` %o��v5���Ϧ��KK�Yc�9�����E�D��b	�1G���Xmk� �ᩤx �ܬ͉
�}��E_��Q�я�.��,2POEU��[[�}�L�
~�-vk�k�(�]����㝜WTn΀S%�B��_�:����_���+C���W�c����P�|�<���Oěm	���O�Ǐ�0)Y������ޔOk��3Ie�'���\羽��(>��jkC��a�����],%����=,�Z}�j���8����y�fp�ݰ�{�J0�]n/�X���0n��-� p��V�삩��΁�S�y��x>\�J�s�I/1�p���ř��Wu�v��g/Ӝ��/�T��1�P�M.�t5��oAA���C_�E<Wo�G�Dc����a�+7>-:��Yw�u���"-��Oam֑t�8ī�P���pӗ;'��`��fBˑt^�Ua�.}��Q`� ���$*��y��M�!0SW���^�#��jm*+E��jr3�/�K��zl�q���A1�]ѿ8fݮ6�[b7Z�ǐy�b�~��� �>Q�ɘ�t��h.�IE�3�TIe[��=y#�b܊<DѬ�S��|=�oP�LM�X4�H��m�+}�����K��%3L�e�#i�o�f��U'�3���р�����Bg�L�I�ʧB�b��k�H�TuQ�)*ҔV�ɼWn=�`�z�y�G���%��O5�]`'��� ��W�X���X��Jfe��d�n�h��� 4�ᬙ}��w��������s'�����',�[�j���Ρ���ZY��X+�Mm"�h�;)��ZZ�t(�\U���R�#���i�K"�g\����fid�$��缟�8��:������D�����
�0�ptm�'�t��>~w�?d�83L�O�)p1��'�I�S�a*�̹��f�_j�p|7�*�z��UG���`��Z;	.~� b��񲐾n'��O�-Kbh��D7T}-�z���Q�2��}��WQ�)�zI��>���|�����w��It���ZBͣ�O�x����]\o�¼$;��X���+V�*0<�8,4���ݏD��If
�?�ͺ�n+���Wt�e���t �J�FK����;~/����{��%�,[9gf��DMn8
��3hqU�V�r�G��
"�ϟ2�b05�Y�Enqd��3m����9���B��$&����,8�xH�%�1�MC�a��0�w��|�4��H�{���N�FE�T�0����.;������%2�@G���n�|�O_��k���)�[+܏��	p?��!�>z�E�z����9��A�|iB*N
6���Z��^����5� �����X�r�C:�t��lQ͵@�ڶSS�3���%M��h����}��1�t��W�[��E��M���c|Q����X�m��z�OQ��UψO"1cG[y��鷤{�W��b"�]NZ��������[�ȵ?�aj@�up��W����Uv��.��"��8�(S��,�♱]$��L�:����a��>�����xg��~���r A��P
�ɅX:�	��|g�$*�,Ω��j��×��pŉ
�(������R@Ѓ�hB=*����IA{��ԯvV`k����S8����8�<��\:�V�����s����J~".�ϳ���(R�Ǖ�e� �g�N0�Z�I�wc�Gx�F=��5�!}��4�ø��v,L�d�K�1�㻯�����Ckug�_(�����l���B�`	�_Aa�L᧐[����C���Q=VJH��?�{�^���߮���}k��˻D��I�F?b��s�i�=�Xՙ�%�3@[�<�	�:<*0���ʫO�}If�=(A�w�}���U?%dؕ�[)����=r	����n��0t�nZ�{��XA/ZK1�V�G����������M"��E�ݍ�p��, �&E�n?\B^tF����=,^���8�T~��������!;��`Y�]��tQD��^��-J5VT��> V���Ӆ�JC=�C���Jn'AS�ҕ^{�΀α��kE���Rkä)�E#	�Bζey�R��KoMq��l��7��`�,g�I���C
ʅ���?A+�8Uq�aCs������E��GS4��,�<��J��$��p;ܶ����ղ�b�`�Z*&]/�8�;=T�5�G��l�F�C��`�b|�ZD�o^
�e���=	k3'aI;����R��2�0�7���ub����Nl�q=�"�c�i�+	.�anK��Zv���\�������i��|�܎�ָ�>dk��ʸ���,��~}!F 7mпL�4F�k&i�N��q�O�`m��%kQ���͛V�L�+.j�.�}�n�Ƕ@��y�@�8�8MI�C��)0��^����+�@�8 ��|�J=ۑӫqyk�	�t�����=�x��=� . 5c�uWd^�
{\�
RɤƎ��&W`j�9~�Z��F�4�@V�>�\��<*«�xu~G��N��sWC��������ַ�d���n����h��f�ɜ��ZD�X�6�q�l@�Q]�v��Ds�N�MH�J�0��ޑn�z.����;���BO����K����;V��h�
o�L����h/+�$�'�I��H���$щk����/S��ƌ7��0���(_
w�`H`4Uw�X�̺��V����ݲ�r�6�,�N)�XD��S�O�W	��(��f�"� [�I�S�,_�dG�����_�șwE����XƋ���������3q���&z�<q�u��ߋG6a�҆�PS#���I��X�K�>�`�z�5�:?�c)�w��ǔm3���f����qM����b�jXH��%$�4=�q�#1�*'9ƶ�ɈVY���&��Rk��}~�I>.�H5I�ǚ֥t�V���dmP�|���(�x&�Q!Kw�[Rl!Ylp��4���H��):�@� g�Hu�oo��~�5��SQJ�K$~H�x�Z��*6�-r�×"2�6���A��������^�{��Q�5}����k�a����m���D�w%� ���`L��%'A��JO���ɶc� ���C�E��_�VA9L#v,wV������������˶�.����|��`��d%�aCb>��i!��B	"D~z��>J�(BR=4�^�"cc�0��R���np�}�Wo�W��W3�	v7������Px����3FXX��u��X�������M���A7`�=>N.�X��]:��̱��9���@i�[����>F�iFjXM��P�;�yG���S�af�W6t%$ �>k�G������gpjlK�6���.���=MD`X̳HL���DҘ��\6M�
 S���#�E>l?�ց���_cCPb��J�]-Ӹ��J�f.BI���g�����Xx��7��?0�D�&8����-i>���&�ss%4�r*�[�ne�x�U�i��w����3�%��]�y9B��������v8����q�־>=�����ֶ�)<���~ j����Le0e93Gϼ��}�v�_Y��Q�Z?��I�d[j�*�r?�����ę����x:p\�d&����(}�U�����r�^0J��َ��Z	b"p���v$����3�&��c��0p�6�����(�5�3�n"���F�W�)i�_%�ü�/��Y�����.�p	[|�־$8��o�_-i���h��J����N1v�>�f}J\�?�(���/�����Y��~�k�ݶ\�SA���K�w����L}��1�r'�l��q�����Xc�5�募�_�!��~N�4��v��-�����`1|RB\vb w��M��<]��L^�E*�i����Ywy�R��
�)����'4�g�"�Z:ȣ��*D���H���[S5��>ņ�x�l���m��Q��J�k�l;�8��u!Tp6��ˏ&ػ��c�$�ʺ�FWd� ?�qT���	�?I�@0�,�,�����/YX�`�#�F��+�x��Ԉ]�k����@ʤ�O�U%%,Y� j�9i�Z(��J��,�LJ{��;塗d ��e}F 2;��_�5��MtO��%~&6b�|�8�o��Y����d$*�$-#�� ���[�;���#%��r[ 8A.�W�����EL�+o��x��N�2]�D%��5�%�ƻ<�d�g�b��89�?�8��n^�q���uF6�G ���������O?b^�P��#��6���:^?�<�.��tS��۲k��Nwg�>m�"r��-�"鲣ڃ+�����Lc�(p<�=�
��w���2�zg�lsC�])�Ha�����<��`c��[c���Dz0w{�::�2_ӧ�iF�Bi��[�#�SЊm�O�`;	9��W�NN���AW5���LB(z����d*I�˥���dQB�����3�*�kwRz�b'��\PZ��'p� �0[�cp��]ˇ�W�M��_P��j�(PM�{�������ɖ�p�84P���)ǥ{OH�λ�L����;-?>����Z�|��'�Q���-�d^������I������/R|}�B�(��#a_b������w�^>(�m��� N �&w�tٴ9����J��t!8ȣi�P�5�r�@^�֢#c�a��Nv{��`�s��3J;�L�2��1Ԙ)+�Ȑǃ$���vn>U�T��e|���{����_`>o`ƍ;��?'L�q�N�QOS=���?���2�:#5$o��v�oȭ	^5N;�4U�Z�E"ZA��X�Ilu��mϼ�Ѿ�:Wk´��:mp���C��M���fN�
�']�^ɟH�R������'�6W���Ԡ;���L�HP#��=�c���<����-�'I�� b9��!*��U8|?|�� d7�f�2���.w8M�˖��Y��*g�<O`�ej�*��E�d��۝�x������oI��w���QU5]�D=��L��x�.�#� E,\Q}D9?7<����4(kD���W=$ъ9B��k��})h0���X��f�i���|(���	�*�W���p@ :�S��2@ʲ��@i
ͮl�>��d�O�eU�*z �vl�եT��v��A'�8�?�A�o=��.�ta��٪��|IC�>v�59���`��a�S�1|">Q����a����|�cCg����F��e��^�">�a��:[���X>�)TL��mT�Kr7U�g�j|H@�y~�����0�N"i��@��U����f�\L�ad�ҟý�v6��$w�:|��j����0�Ώ &�4��ֱ$�о�06J��(T��������$dU��w	Y-�vfM�-�4��r,O�A���I��Ϸ^(Ø���֐{Z���Iq�ǟ�z�?hGp-@fi�Zb����Z�D���\���ʡ~���[��`Ot�F�i4���߀��!O����gᩱډU����KUZ�Q�u��'?��03)Z��6�z�Į�]�}>t�DG`�$+�T��&n�>'�tAs�r�I�o����/��W+��q��5��:�����'�5�"յ�L�
�ű~���)����[���<�[��R�$�>ͧHD����gG�Mh�7!ժSB�<$�����'���R��_\�
#]�R��cheI" ��5�������F┪�Ɯ�ʼ`��x���F��F��)��; ���#K�[&H@L�t���i��1Z<��uz�O�꼉�!w.�d�����芞��_��a.`HϘ��G��E�y1�E����9��2��?��%k���a����H$�%��Xu�&�Y�%mY��H�'B5{�R�b�Og�+��uC&�㬌r/R�?��:|��o�퀱��B�h����p~��ԑ�qm]�Uip�ج٬vw�Qpj��8{� Q�S���=�wi�~/�緾C��Ѡ�2���x��O��
c%=G�O&~�ڃp�L�6:r��E�z�Z�n�`5�넺H��+3��8��BT?ou"�7e
E(�j�U��q��u߾�p�Q*�����H�\�jȪ�L�.�v�(��������I��q�j_P�յ�t�͉O�khr��)0�P�|�@�+�.C!���n	�6+�qU%��FS+W3�7=vw?Z-zܾ1���e�-�؛�Gw ����z����u�����I�I��?�易My7��{hC@"Y8$��2���5���?K���zհ#@3�h[|��G�Ɍ�iR�j�� �ԸM��_�����)�����,o����Z��I#=�4��;6����}�jxԫ�'���3�q	�J2�"V�=_b2
fe7�HujD����ZKڄ�Ջ"�?r*��T��{ng�E��wXG�iR�ʾ�W/g	y="򶈬�@x�����m=x�hv�\��]�u^}���65;0k�M"�E�G�B��y�M��&��rzd�[�Rf����f0t�2���R�ᄜ�k�7�c=�z�R�#2���r�?��lG�78�p.>jE�@a�$�m5u+�XO��.���g��F�+X�a8.K��S��9�U�,P19@9*m����*ϴ#Z�
w��PtJ-��5��.o���'@���/m�˝lH��3,+�k?�@S��|<j].�y����I٢�\^��7yV���ʼ��d촫ȷ�����%M�V���q�m<�vڞ�Vu���&pl{�]�[�״��`'J���q�B�{T�O��;q/�=��<�v�a��]2.��8�Up
�M�����Dg�G�
����<`�f�c����(�W_�0ݾB��%�߭��X��\��h���B��:�ݥ5�m��*�L��]�9�Vm�Oh���� WCd����.򉴶o`T* ������"��bߪg���d�R��j�Y}�f0a9���߮�B�*;UE��ef���HX��K"}�:|zq�s<*{��9�f��8*�m����~��=6f5�i���;��(`%�:ئ��f��,)_'oF�ֳ��H}����@Jk�x��=��u�Mc�4=�(xXAR�$�9o/���5j/
q��e�= =f:�&@��L�E�J��6ݑ�%��g�ݴ^R7��Ea�5C���k<�\Ҽ*f Ӝc��zy>�%]'�����r+�Be�hf?fw���Z�a���R�72nb���/��[�"�=�='TWb'ت�04K�!�q�O�i���e�0�2 ��3�K��/�x������WWb�Χ��O�t�e�� ����D[��	 �:��73�I�ɕ�FF@�*�����\��~���ʧn�U�5;.���#Rמ�C���O�Ң�'`�N ��q�[Hn�
�ˣ$�0N��u�7�;��S����K]F�+Y�� �m�!M$���tĻdb,Z,��(#J�Ψ�D���]y�W^K��4�jx
=���T�96�G�ą�i8C�YhL�Ɂ.�7����W���$W�>i>���I֞4��o��>e�P�\ܜ~��L��i�o�'�ϱ@�_�V�G�z���d�\}��lSX
�!2�Q�:�u���Ͼ~ϰ�#rԸ�����|���o� ������(1��m��VGNn��'jE53�)oO˺u;ߊϺPI"4S���8�ד.R=�W����F�u6�=��mW/� 0�4��jY�L��)]i��E�������l#���=6�ϖ�U�o��Լ�{,�|U��h��,]�p�\L��Q���Z���Ro~Jʾ����ch�cKS�sR��ޔ�(��V������7NF�����l���VWo����ܵE���.F��bKHtd���`X��3�Ybs/i�,B�4(d~B+sB|�?����V���޷��*ċt�V�7.�g^�>�w�uk���$<䡀�?L����v�_N��]����*� &J�u�c^��Hӓ��⌺ߑ1L>�d^K�)�ZH�m�ߪ!ZG�A¯A�1t�-�G��Cp�H�	�K�%g��29��H��CV�DL���2Ɵ�1�VeA���*uI��`4��jY�C;�p�[	j�E�œg�~����^���uuq�]7#o�{ ���f?Uy]9M)��}��~Kָ�2�[�FZ_0>�ÅS$G㌶��������3s���������	��z}���{4�'�p�f�v�Ś	���;��+�!�1x�s��G@�C
��.��@q]���'g<{���%����D��z�K���	���/\p��(Su7��e�)͈5�wV���st�Ӏ��"�.0�zV'��+Ӥ���di�����O'�M����%h���@�k<7Ne�M����^r@��&�v����*���h*���&�3_�^�8�!c� 0�}��,�F��0~m�P�0g@Ģ�<d,٢ȣ�)'jg]
�HI;]���غ�	wÝ�ޕS{O�C�|�7�ޘ��3��������5ǭ����џ���T���q�NlA˕�V�=^��qY�+�um�������iҴ~'A�+�p��M�ܗ�Þ^eƧA�NRF$�c�ӳ�<��	Vg��Qw��&�.�����7E���O���8��s��m*~�8���3�#	�Zߍ.�E7��&��D/�
�CJ�q�x�u���n���!��Tv�u��:7�og�>�9�Q����Ro+lqw$�]�(Q�B㪭N�K�ZE��~̒��.�U�E3(��d��e�!ά��N�z�ԑ�N�F����Ic�X0O�X0Ѽ���-�G�j���%q�I�s�y���g�ס���d��D�QR ��W�۟sAp3ocrp��&�$��]�?�
u�,$ռ�v�UbX橚�.m?�Vjy�t�ؘPh�X�!\��4�d�ˤ�yqB�B��ƤN�Zj�u�H�K9�%L#��	c�o됗j���'n�T��t~\9����~Y�:�����ə� 9�j�M�˗	e�p@�E��F!B$���==ii�*��X�r��-P9g=�ARz%�v��H���h��1��$�p��}� S�óv���C��?ߝr�?]\��hFȊ�+G B�n�%��	M,�kW���@���'�i4|21�u�jv��@��ƭ���-1�䃎!.L�"�<P ���d�A��)Q��?�:c����/}�j���#�A�\)
|�1ɢ��)��7���ZƱ�����3�Z�5i��D�V2�F���A�T�^��v�{E�֔�{�[[�������ߨP��c�����5��9��m�����.���3L�d5���-��ppp�6�2`r�p��MtVO�����դ��]*�~�s���0C5S�T�Cb�UK]w5,�����m��B��8@=�p���YrJ27��x+�l3{��R���R5�r��T������ď��|���h�qC������Z���0&��G00�!�Uϴ��F�>pDԐ��Ѝ=����u
��7-�E���f8�'���X=󾠑=:%=�$]f���r�K�����1..RyO2r���d��a3p�T}��RՎ˱H��6d�٣,�+f+pQ�_��IH�ػ����Ŝۼ�"l{<�K ��n�ߗm��0����x�z=~��@�J�N��|���6v����4g�#G�U�^�����p�?u�:X�����c�R��� l"�T,�ƒ5�8����v_�([�_��G֫^X�3�N���$d�O������+�7Vt�%�٣B���i��-�S�g.�qFHB䀠���)����Ep�3)�r:����cT��q�\�nF9r�>�L��ﾶ��h��aY�D�(����#&T��ci"��(ͺ���B��j��r��%U}��4�iT�	/wG���dp��Hx���V�!��J�
Y�o�����R+�^�q#B��Y��\�߄�|�%�a[guV�w�ׄ9W�C��v��ʂ�%�48k=�JY�>��x��WG>wa�Uk[)���}H�To]$,甙��GC!��03B�+$5)��4�*@�Ȫ[`UB�zoeU]D�%��U���4�t�IW<��K~���?�b/7:�]�'����n�,��L�l�3ΔDVa:+�v����� � u�PB���=
��+e�5,�w�ě3�β�Vs'�<� ̓�c��b�֓�K��oe�"2�d*lLD�b����d�Vg.��`��_���}�t]�	�4�i=l��^����`�TГl�b�ݲ�W�4�e[ $Lo�T�
=����u?�ؐ�a��,Qj�{�5�"V����/q�K�Gb��~�@�=f�6 ��������^8�inwk���/��@�+K�~�JH�N�3��
^O; }TtW�|mi�B�Pz�M���P(�n�5S+$�	�Hb�[��\&�θ�B2ډ� �[���o�����?l�0�Z��a7/7 ��?Tq����rS�J��?���MI%Ҩ��	 �\���:�a/��SZ3l_ �٩���(^�WfriÐ� V"��H��zIeM����TTʟ���FO0����BE:�Xe1�>y��a#��T8 }�E���!I�o�㯢b�sfK�.
��+���W&C�K�M��`��7�<�.W�
�����o���S�8Z;�����r����2m#Jf]=qJG�D9��	wv�6�)O�_h�����?1�vh�j����z�+�;��;6�2 mg��w����6����c�wSdb�m��I�b#��4�\l����{w�^4\�M)�ʧ��O`��=��EC٭��h�7Z����g�[<;�,PV���Gw�`W��������5�iIt�A�s����GP�U���A�	0_/�'H.�L뜈.�9���V�&�V!bKU/`��#�@�������6�*���t�4m�"��I�Ur>��	tò�I^�[w�]����x+���f�y�T���S�m#�F�D�]�]9�L�<�=%(.l�$K(f��V4�*k�$e�yJRh�i+��� ���a5J��!�"�D3��:���Ĕֈ����<�2bg�H�o�����,�򋱵��,�(�.؀�G������|(*P8|㼁EC��)3��tt�����,��[�?	V����� ��@`e��L�Ͷ̨�rZ�3'�lyt��K�t�e�
l��dbdd�ɀ�d�՞�V\�� ��dWq�ά�e�\RZ��?����)}u���U�ғG��ˉ#F�J�6v�9�I�	#N�"���qo�`[����I��%Ƞ	�9��ҩ\��3R�w���)�,4��!j��F9#բ�9�M]��!�x��@u����8X���.x�7C�:&�tI	v�����v���@�E��}�PC���� &��Z'V���.���v.Ic
R*A��&�N�ޡ2�yt���a�h����ˌ�PR'�zD{�6� ��6d��i}�/f�_�C��.�쿧��k�H <�J�#j���U.;�������!����Y�Y<�8��.�w'`����*D�$83:S�0sh�g�F{�{e�M�F��#^�m��U^�Τ��9��v��r�~�+#G\��KwG�@>�Mȡ�UhoE���n_EhR94)H���|��د��ɴ�o������r�5��8��m�81��D�z�� �-�ȿ�pP�pDdcu�&^��і.�α.�@�7vދM�����܅|:+�,���y�yF�WV�l(,�yt�!�8b�(8iHmJz�EE
F�ң?l�3��k�k2�z�F�UqZU����U�A�[NF���a�7�>T�!�B+��SV"0��\�FB�e@M�Z����>�Rz$�]��Ó����A5����R'�[�vU���^�x_If�&Kd������4����%UsYwUb�#���`Mg�Ve�y��qu�߈�T��ڇ�䬁U����iS�{�|�Yb�[� �]ځ�?���!F��^��>^��ST+XMy�"��/��XBy�
��^;cʾ��ޯ���2�R5���,\L���v"�X����|��²�OB�����?j��Վ7����`�X)�ov�Y��X�Ο��W_���gJ����*�4 ��&o���hW�,$����_Nu��q��^��+�G>3fa6ç�@��s�(r�*�w��?����^�"�i�-1$�h$Nl튺O�欉�<�Y*:�,��@z�^�����?f��S���k�H"�T�9K^M��?:"�(u���A���Z���ɺ\��w$�O�=�Ot�U���Z^�:��
2��M���\�����ua&�2�x	P<�����f���T���8��d�C��'gV��#�~�-4����a`��n�,�9
Lg����@�ǐ2�T�y��3/U��k��w�<�C
	dB���yD:��6�㬞���r��9�.�͹�c\�]�q}��'���fO������E�ªʣ �;\S-#�_�������&�Ĝ�9�a[���k����d�Ӻ�;�Q����U��/��tHKýǅ��"�2�k ��@������B�PmqE��?���A��+�VHK�iD!�Oj��=@��f�s�"*�
�f]Hh�����h_K�^GАG"�	D�]�M���K��(2�vN��� -q�����aT�F���G��<[���<�p�[ �dA������57�^�P�L���v� �M\��IP��$;���u�Үv��+L��|�0���eǜs ������7!�y]�Ge��02�gL:�H�0�]tw."���d��j# ��>���3��y���S�H��*�y/�w����I�0C����o�4P�p7W�H��b�|{&/�e�#�0:fkj8n��).��v�Q5�p8�u6�\����uP@�:XQ�̀a4�p_m����: �L,,\��le�j�1�գU�0�W�jַ
��A�6�\�7�ҝ> ����A$�ާ��{��%�ӫ�"��uQ����ju��1��=_>2�cԍcֆ,�pH���8SNAD$ 2H� ��Ҷ��y�o�W�����F�����>�Ϸ�&������S�W*ř3W���>B����OR1w�ǩ\i�|Bj�V]г�2J�D7�@��۳��N@w�����%�t��n��3����lzi�׳�,���S��ir��ү�f�K0Ω��:T��6��qF�EROȐ�%i��k���-�fpRRB�b0,�$�wXȂ�d�(�I�L$Y��!��W��wE�].����a�9���t�{b��y��m�ݕ�1B�m-e�b�_˪*�Rg���+�׮����dDs�@Dv��N{��.c�jr.�1]��[����zE�u�$�,���M�����j�3�£I���(Kr�TK��ӵ����׾�B���Y�8x`��5����>���k���O�=;�žE���89��Y�4Z�Y8��tS�=5���;М��{�;��Q�:@��s��fN ����~�G��VF���
e��Y�uY���ʃ���
�Q_�(���]m\���<�W�Ĝ�HG	��{	��K�.Z�	@��!��Ζ3kq�~	�MAN�:�H���ϟ/��N5Si�����k�xn0CL��]�d4�B�#89�|84d�i��p+R2����g��}�ґiZ.�!���.q�p�D��������Gn��H� _	��Mج�Xڎ�	Ix�����^���yvNھ�^�]9�y-*>%:��"Z[�S��~���`�((T�R#��5��#��6<7��㲘T�b�H�'��x~�b6���>�#�-�!�D=�h#�����Y4���~E�hqjG�r< �A�¨'J���v�i����7S6�LX]��'V��|��zz�"���ق�0�U��|��)�=�A}=���{�xg�S
�|QY�[����$+�Y{�]�D-��A��
 )�	�0�S�Z)������nŚ�,���Q���PĠ�z�J�RK%�&�v������{[^
�EYsZB��F���y<\�P����0����/��4�4d����e���^v��_�����-Ӹ� �!Uf��u�F��g�N�Tt�(��'H	l�և���ۏ���t�h�,����n�y0�L퟇�2�����i]B�d[��G�?����dsW%���]�<��8�;���]S�Fs��k�{]>s���r��������;��^�O��3
i�@V6dӝ����Ȏ�SԦQ�f։9r���ll(qn<̀���-��:����X4�C剢����%	6[��3X���s3�0Z����~���ig��ʹ?	������6^�;� ��SG�gs,�3�2u�a�1��Z[�����B�6�|s�f�����푾�7�/�
�~�t�h��D�(�KRoP1�[���k"�h託�
�g��e�n��6�-�\>FI���E̧���u'�����-���H�ە)�LRgj#��g��<E���D�U��}�jϭ����=r6\�)w��j�"����!z,<f(쮀�$^/2�����ðďM��x��}�ʡ��E���t?��� ���n����ߕq_�*[8S��)k�A���&Bo��6X8<�,�Ʌv:^�|L�av�����_q�U��"�KN��
����nL�����e�8�'4[�������=�Q�)>eL�,wd�\� �O�R�ŸF�l��(��{��$[t�9A^�T�+]n�F�U|`�o��M�	��a��d�{x���f�לh���*�C5^�=V�św���BϚ�y�%H���t`�IjT#�^���(ף�y��Ō��_m�.�[�)�d/C��\��q�ۣ�B�
F���f��[	�������?�:4�'�2 7����m��:)"��M���|f��[��4�l/�B9�	�_�ë�L��}�|W3�)�����P�f6�����Ms[�\�Z
��K5����:�ʙ���ҩ"��z�G���_�ԏ/L�~�%]zT���o���GҨV����ΒԹ�ـXpU��H�v��*U������R^o��UQ�R�����+N~EXk�e�f�����ĳ��>qcc���Z{!�0S������Us�!�_��������v^ �%1����cY��E0���k�#�`n���m�`z�R;Os����Nf���lmN�\�K~#���do�|v�M�����N��W�4�Wv�����%�6C�"4����d�)�К`�Z�GO9�j)Iyhŏ�2��N���y�U3�ڿ*������8�����sA��������;�('�9�S�9�
��y�Ǥ���p�����c��?�a�όX�z���	枂c�8�G�b��9��c��
�N\�82ɉ ��5�j��I�?X��.��׵߮�]����Q��S������3�=;��Iە#����U���=-��D+7�������^-@��"����z�����7�)Q������*|�-����J�M��~,��)ۛ���/�8��<Of�$Es�̯e��T�vZx��5�?R��w����ڤ՞��L� 	���/�z�I�I%�ٽ+��(�cB��8�s=N»FM��ڋ��w����ޖ�U�uJ��0dx�zz��A�֥A�������qgW���%�����b*Ȅ{+�˄X��G��\$��H����{L���;p��H7�m�e���ri�w�@O�`NV�FKW]��m1�O~7Tq�%�ڡώ�JA�9.4�\�@Xk�����d�Cf:UN|����z.��wz��������uӑ3s�������2�ߊ�-p��ȿ7�u�JG�g����8I�<-1��Em��g
��k�t^��nn� �*���5���y5W�:(eb�-�O�&���x����}z�4��h���x��w%�k�"����w��j��OZdkv{��転KPc!(����Q��=��0�g~j����[$ [wP%0������g���^w�ʅ4 ������T�.ɭ����@$��W���fk������w������skM���f!�Ww.�t=u<��J�J���-RL~"���=,�s{@�!�	�b��� >��~�©��ѧql{٪�����
�5�# �X�䝻���Y%�_�f욥�d�(g�D;�<xChG���+د�Xd�/�j^`d�K$צ��s!�-	�TL;r=�����N#���j3��0_7?�o��"���!͋��J(R)b�����=)vɥ�����ڮ<CE��c�����S��:+�%p>r�j㵭����֊���Rb�=*���][Pb��=Ȗ (li�\o0���d(F\-�~V��.��:�ç@P�v���u��>Ք����_�9Y1$��)C�����zƎe���!��]�t��μ�Тz��E#	���cm;����u���o��??Dm�n��.�:ۮ�� "Z�^��ȹJ�n�+���S+�["����ƿ����J��y���K��TEg4�Y�p{���A��z�<@���䀁�JA�8�e�V�h��͞�z��	�:2���2��Q̋7�cX��o�+'��>*T��������n�G��t"�N�;�'w���.�Vf�u����z��Jw|���fӉfl�� }��q�/��U���0�`'/5��4�g��w�A��RLƧ��m�~����k�� ��{�eE����ei��4�;ZE����hW��z���7g�
3+��ʲAN��7m�`�v	�*P�>��^�т>M@�aCY���5��~�U��y�_�cʭ!�׃_ZQ�C��ҟE=�,<�1�tʹ��q!W|���4��k��'KFC0����Q�5�]Bj��%#��C*�� c5G��8�Ը���ࠊ��2N�v�"�~�?��Ұ!��1,� jc�������R�����Wק��K��ͬC'��bHD������R��̲�7Ȯn���c��-��ʚ���cx�|^��l�HG�U�ï�,�2���2`�����L�Qb��%HQ���:=�Ta�f�e�O�X9'f/�Q�h�@<�@,�x����R�|�8kl�2QM��;�$o(+��"��̱�����/
�s�?-�&'#N'�&Q�	}/�I���S�u-�C;�'���Z:ա���Wa��KX�{mr$��b�2�J �jL*A����Pb��7.�������a��Fڭ4��G��j@���}��Q�[�06ⅹm�X����kc��$���a���dD�q�dD((�����c�,X�
�35� �Ơ�8��h?� ��� ���zm�I׹uS)�{�[p�t�K���n�ft�C��3_��)B��f�q=*ȱ<�"��J�� ڤ�g�R/��hS!ڭ�eAw{+)H�����n��&@a�޶�t��8.�MԖ��O�������*K�s��8�a���{��۝ߦ����b0`�Y9��`*�$�W�I��D�<֔Z�K5�N_>j��XL����3"-L�o�S�I,>�hj������1���@�=�H� �"g�VJN�k;'���Ѣ��s�o�J�E|�g�<Ԍ~ ��㳵P)�*�~US�v�E�����i��omH���maO��h�����9�/uw��c�~�<U%�b�a�m�O�"|Th|�����? �Nk"�,�b�A��Z�i�sP��QPWr,���~y��V�첊4�&-�}���s{�����>¥:�=$�8uk�"��N�dIG����
���)�����)Wf��%>O�ѯo}"���m���~a�Ĕ�n/5I͢ ԃ<-�Ӡ��6�V:I�:c��oZE&1W���s6�7L�d/���A-@O����û��D�Bk?ES�:!2��Iu;��_ [�'^��u�����s���-�o��9ݎ����6O�����!a]a�C����4�,=sH�ۭ�� �i�F������;�-�a56�><ZT ��j�1U���eb�^���_�j��=����H~���J;.� Z]̱�1����=�"::o~�}�_	������ѕ�5�_cvu#�s;�� J��k��S�� h���J��{g��gє�[(w�O<'�)�N��u耂����Y�f�\W�	. �O�gzܨ��=��?�5�TE�M�+)�2'�:gC�?-���:*��1@^�����0r^.�$��Lx��j�:7���㳛�����U��̭���ԁH��.�.)�^NP��sR�'y
��Nyw��*x�vsl!X�� �Yɶ���~
��}AE�J�O����|M�Pdh(.J�J^#�����U\�G�J O�[��s�eHݮj��ܯK�j���/����5_����'����V>��³vU�<��8)7t�CҤ�D{,8�ُ� dB�ă�)c��C��[�8�~W��A^z�Xy�X�>���e�2�2{���a�,J���QE��FF����[Zh���o�� �4��^�ւ���2"��������U�[�81����E���b���N����S�UN�YG,��� p��^K���\��X�h?�A�W� ϡ ��m���%����l���Ǥ�-^e4�,be]���2Ȍ��_�5C��W�vH]�R��{��uJlL��y�9���I�ڹ2/$���{����4S���9� i�W"�ߴpj�2Q�X��ExW�븄�y~�:+���#��� 80rN�m��e��"z=�p���5�^�&��(� ���K�܂���-�`�!8�i�����5N���(�^��u6o�gT��Lg�_%�)~Rc<IEDe}\Fx�H鞱�s�1��C�����|��g�iכ�u�xu���%�܌�ԷH��g[t����@Wz��w�
���̠)T_�1u��� ��1����|�]�����a-��9�o� �)��*h�}CDf\�ʋ��#�	��G���p�|C���k���cY�M 2Mb��V��>�Q�n�=%�nd~͆�K麳ڽ�QF���N�V�{�=O�>r��o\h�Q՛����z�����u�ʺ���r^�ea� ��Fm��,�Ʒᄱ�Ճ�$��ڽ��C��I�g�.��'�i5������]���q�l�͏��=o���p��N��LF*��xZ��m�rf� ^�P�.;�G���X�9@���� '��Y��Q��N�.�'�,�/r��^ia��r�/d`�a>�n�
:?T�g��j$�P�CF�yq�J��h�d�E�ß���g�:���	�0���+����E.W�=���ʓq����8H�`@�$���_lUH��$U����[�\j{�k��I	qeMT����X�����_):��I�r�(�� �������BO/Z�f���U�͘bNVbMr1}�)��&�?��ꛖ�X&�!f�q(Ps���ռ4�!�D;]�y6^��A�@�����'vk�oeq�خZ��ss<���Ǭ3� * �P�����a�@�&jY)���V�/Ä����b!�Y�,�[�ɖ�Sy+�U
��-<}��z!��!H����z:�\/��NW����РL������uY@*�-8y���x-;��|�&���ևCA���_�zf��J�ynA���,`��?ZR�[�f]�ن���
�V���* ��L���R2��f?�v��A�i�,�aY��T��p�������K�S(2H��;_~Ƣ�M>Ng�:)�/	��+�Nވ��3EQ�vY��z������w#���Rt�B�Q~.{O+�" ��x�ψ �5�=
��:J?���~9nS�4i�w:ڲ�-���𔻡C�)����#�7�bK!�M[�IA]pe%o��ϵq:��&gJ����sq�}+|�Y1����0�ܰ>�6r�_�4ku\�qW�W���h��pEL�2r捦dOq/��gy	���=�M��2G8]'��&�յ�";����mH.�T�ko���{QlХ�	�y?}�.ޢI�\X(nN���I�L���� ��(�"�7`����5 :�G�L%�߃���5'��)6r����� ��o�b�2�&\�[F�W�Y��,f>i?���(�n7�:t�nf/v^���t T�6Ԡ��qS�r Ҭ�l4����=�b4=�ܺz�$��u�M���m��X|�R���1��VR����tmh��1���c[+̭�k�`9�=Ĉ"�S"��j6z�gqu �T�2�#^��-~�B�<iۑ���O$Vu�VYn��zq�x�N��Ԧ���Yl;7��8�`7H��a�[�r���Of�i�<0c��d��W���N�B}$�؅.���`3��Ғ��YC4H)* ӷ������=O�y4(�k�t��d"%G������$�%=8X���̈�T��3�l�����w8*�=e{ː���v_��)�Flf�,�$�\S�N�.&m�\FKK?��u�VK�Qz�9�wqu�*��<�]`";�J�Z��j�[��7���$��^�����IJ��V�"qM����M��8��ֈ��LR�CJJ�Ff�,�@T�+�Z�
��$���D9��q��{k��KԹ���W��6�"��WIr95�t��s�5��mի�L6�+�)g.���
/���AC�p�iN�5�QW�/{v�i�R����1���w'���ƥ�k$��~��d<�tY�)|K�w���KIu�c<���{h��C�M��L�m5��b���H�A8*�t$�ºl�߫�y��	��}5��h�����RXe7[mQФ���h�E�:u2~M���a�	��b)�>D1H(���Ez<���.S�� �\�Rʽ,�s֒N�:c->r;=�4`�AV5aU�Q[O����^��K�>�7mHB�y�	R8إ���f�l�B���_��J���˫� "m��m��$�fd}�Ǒ���ʙ�q�Z�:x��	}/c�����~tO�^�FXLe�y������d��x�X4�B�����5�%�H��nP�q�x����*@]��?
O� �-Gc���������K��B��#i�0�TD��&#j���͓��m�j��2B�U�%`���R�lx�z��6R\.��6;8�
�*ء&y�#(y�[$/K�LH�׮��xJJ��5�+����UK�w��S�ْ�1E�˂�a��L{��MbW�q��>A`���6Y�9�fk
� �K�����R��0(�Q���2�o�~�Z-��)��6_<����8�8\��?s}��wK&�j찓&�L���w�Y��AW*�J��ŭ؋.^z3"��CȻ�1_r���b�}��r�|hCA�(N��v/�+ ��k�<��d��Y{=�׌��/�#��j+�ב�3öP����;&�d�&=�Z6����h�! �������vr8��R��4��Ay\
L�R����;b�|	�%�q�;���)�����I�hX�_��k�\�;B?�Р��UJ�{�U1�v�g��:C��[��q��ol?"01�d��m�=f���4#���A@�E����
:Ό���[Ф5x@����w�11�}\(��dQ7���qa���Kn�ʦɬO�a�x_�o�v��~�%2�>�� ����qT&���f9f5.��W|��ajb�e�?e����76��TO Vɢ�ylBXkt�Z�@r�����5�0��q�Qs!G�j:Tf�$�:5Yl�����a��!�.8C��9W1Av˷�ȃ��+��.P�  QƄyII���g�Q����<��-	W#���+�x��]Kc����#�)&��t���OX��qև��(�z�U�,$�x7J�-����jˍP�񸸶���8�l����~�����L��aVG]1赀�`�v�r�A}1֛�8z���= wX.VɃʮ�g����m�^��&P}nZ��O��#���H���p�����R�I,�u�gŷF�/����9���8��h376N�K���S�q�P�� T���Ե���qp��M�k.��M��$��VGY����������ga����p/(n��!3�Yg놲���WW�拽d'�r��k��/�e�u9������Q�7s���0�EV��Ck��Md���� ��%�z�[����hU|M��*�T���t�*�}��S�Z�5"�|L��~��4�ArV$�����\���'k<�7æu�%/2cH8h�%�n~����,cI����ʼ` 3kA\Y�P5"�����+,ڐW�t3>�[^q�3~�O��{U�f,l�@x{|6�`�Ӟalm S��I����kVI8HSaC$�S|=��u�`�U˜�<r5�g�����(��8���ho�"�h�@@�^���lpɍ�Q��A��d4��RW�ig��R"�N��wDcW�k��a%��z�����D&i�{�5�9H֏Q���q�Y$��1�I ����Zؔv�(6���3(d��p@tf�U�A�j�N��:x��6LQ�ҴG˷z�7�P6�5��&?p͌鞚��M[[k�i��$�����H�m��m�6V����f�?���]�Cv�����|�m<(�%�.6D�z�Pk��m
w�	���!$��:'�Sk>��u���� x���j耲�U�<�ZE�C�yV��)�f�V�F��
o�,�y��A+��_:B����s>#!Ic9�����������P�
�t5���.�f��[����'���3j�x�]������Vî�FH�"�9�Q�V;*a��{��`��/ڬ��2�do�_0� q�Y���k 2>-V�ϢږH"�+���y4��ف�R�o���B�tUjK�@Q"��Ш�cȃ	�a��k����e*�TDU=��f��f1՘~ɓ$�d���椓�O6��ɱ�=�-�fi�ou����;+��]��*xh��&\-�?t��x��RM��Ø��s���'=�Eb�|K�c�_�g<b���E��9���ZEYW�(�҈p���`E*\�=OwvS֏�n_Kڮ�+w�)F�y�nB��h�b"����3�ܶ%��)7(Ji�x|s���|�_�V��X��U�� Zi�G�6�Ջu�.���sMXY���;���6�i��x�F~�[o����������_���=��u�#}���Lj	Z<�OJ�V(�G�-�a��&g�L� ��"�|�Ƙ	
[���n�9�x�5��k����O�թL%Pf���[?���֭�R��������s���0�߰�F4����i��Q��i.��aP�}�3�\�/�^4c���zxkH?�u�5EuŶ�ԧ�,��G���ˀ��$�i�}.$�FA3_M�F`���f�Ѕ&��|Nӵ�q����L��Yh�h�`�.'�([��T�ս�C>� .����9��Y�d��7�ZkyŁ[�h��|N^>��r�I����/���ǺI�?���(����\T��L��HK�D~!�X���^��p�z�h�Y�ȴ��
>�	hЙ�/�ioU������n�_��5���3���_��WvQR�m�r�ا!�=&\�gr� %³薦|s�S|���8&�	� ^��!�i��6�oB��b���es~�U� {�.(�Ό���55�ٿ��*��#2��r�@�3�2 �+�nȑ*�֕�]�f����ܕ�n.^���g}xQ�/0�J��r�J�U���u5�|z|9.ī؁����m��ߍu��Y���&���&�/&r�Y�*��bb�Ƨ�KWՈ��?*����y+>d��ֵ4-%��#_��Ê��1f�m=�кv�/��N���D�s��u�@�=�O]jk����F�q�V�+���3�x�V7���ȇ��H��%:f���̀.�ё!�t��N�u%q��ϷT��0�ۡ^�`���K�c| '��q�B�`�ӧ���<�87���.�K-��x0���T�0Z�wŦ5��.Y�F;��nw-�p�>������//��n'zz�_s Z�-�I���L��/~b-"6��|�&���_�3��V��nG��h�+q��4�A��?7�ZU(�g����vhGO��G�!�6 �:��0�W���5?��c��pǽ��^ZM��z�o��0��l\wԬ-J��]L�gaS�l��L@�#�n)�M		L��j!�v�@I$�U� ٚ��sch	r����z2q����̌��=������<���|��8'��^�}vw��M�9�z�=_���;�`gg&
6nI��4
2�}T��	�%���o�>F�t�߭�i��Srڍ�e��i:�w�̿e_>u��:ļp�1	�6B�	Kx��k�W!���]�a_P����Ú8NW����>'�l�~<�Kİ�֏%Y��s��d�/���E5[��C�P��P�D-�������FMiZ�+*��V`��:��A����#@��&�u3��by������Nq󂄢L�7��V�+���ڌ�Ƨ|��8� L?�n��ֵ�Ů��~Gc:+5��8:�۔��6�Q����1h���_�:�ԫ�@(��H�papƗL�薱*�d�Q/��>%Ҡ��"}��
[��#�+L�΋�)�K����N1G�+�)]iL�`:���9����"b&���ԑ���P�X�Y��;0B�N��)�i��G��o�5:B���9/� `��IsX��Ё(��Ʊ~;2e�H�š�:��ݧ�<~��RRe�c�`�Sv]�aM`���N�tpL�����<"��8X�(�^܅n1��W?�U\8��@*{�Jn��QlP���_��ϐX�Y�oZA�1�G0���#� y�m���kT�hy��W��v3/�ɺ��m"S������K�u��DP�At?),��-[ ����2�4���Hb:���u�O�5�y�Ls)��-�cB�ҊKj��h�u�:���vv���޴�� $�3�xR�]�l�Y�#�&26��iE��m�%Y��z��!��D��mJ���
�[��^�!t���������ZK����l!��fhȃ���Dtw��8���<��Py�Nt��l���)C��r��_����.�E���jZ��v�3c�}!�-!xҀr��@d-h�h�fi�O�,��#�W��x?O#@��]&{GFvO��ډ�oaY0O���5� uy��H�k{�wKH�kr-�X.�op�E����&���`N����/b�!��w�i�)i'�HZ�F��-E�'���×@)��[	_��1�Dk���ď !��MK���)E�yx}��N��˻w��$�����6��̧�[	,��ƺZ[�i2.2���L_���8�eXP�?|k쿎�}s�6k2�$e\��-�Y���I��<ŷ"FÊ������Y��fZ;�p?l�����;�ƛ�=�݄񆉼�,w��J�����T����߲��g���UѽE>n�OT?��� j��AI)	u��c��"_�N��`7�1F�L�j��:�>=�p�Amdu�z���f���4W��$�ŴD�?~_���-��ut��#����T�f��X�c{����)�?�*M��}@��L�� ۯq��|&�c���>莞<1yt8[�9��6Y������)�'v>T�b��%|F�rE%X�`�P��	����-�	2$�[y=n)�������L��IAv?{�~Kq����1/i�1��D["2�Fe�,={]8UZ'J�]D� ����i�C�!�s���7�c>ŀ�^S��$-( l"��kw[�j>�C�rsW���Ɛ|fM"�b�n;��5O��ǝ6�'�W��L�$�⣻a+`��=����2}W���D,���<B�/;���f���y+gb��50#���IfVExI��1;��>���Xe����Y?�o��k!�ٺ}Pͬ���8���X��Z���	��[/� ���l3��%v�\H2i�-o�\��q
�>�	�`�a���-�B��/�PDyr��Fx��<iw(+�zG����d��+�i+�95���T�z׶o�w�d��k�Z貁f�4c����Op�&�A�-�=���s���6nG���Z���:��͂�|��JSM�<0�g	3�#f8ӌi������SC�#P�}7�K�d��>�s�6z˖�Q��%��u�;Ac���D�W�!Q�ì9��GS�l�Gߪx�װ|a�S�^@-���Q(}4t�5ʬ`"
����� 5�G�_V"�k�����ς�c���fx�d�#�~��Pj�ۯr��Ǹ��/��.���q��V6ꇤ@f�7$����^2q{q�Z��q��Sm�cI��UEΤk�f�re���T���'J�U-R���F���8_��u�7���R��ۿ�������7��jso&n�f,��M�&�Վ�F�7{�]�j�X-�l�s�Ϭj1���_��G�+/i��#�3�6���*�3��yLF��� k�^�+u,�|��N�8e��k|��z���l4��
�LH���N�cb���������R�1�zS��ӻO��c�Q�CMN/?uFϔF/���u1�K�)�ֶ]3�nm�)�\D���C(��VR��,,��$��IG��~R'�j2�륯h?� �(!^,B{�BrwRYE'����l����<��byu��:�,=�'.�v�xۯ�#ё��H��\K��)�G;�S�@��c�+j�j�j��Y��@���ʵ�uSu�P�����~�9�_�zH�&VQP�9-`H,�_@�@"&�w �\���2��K���F{,p����h8��9]0z�cs�σ"�4*A5J5�r���g���������Į-L���ď͌Ÿ�/�sv�k�d�߳�V7O5z��Z]i�;��1��Wm�z`8	��{m�������/`���P�؝�d�a�Js�8Y�0�Gu�{�#G����A̜��QH[AӴ����%c���ش:b��3��M���m74��4���Q�}���^���4���ݭ${ Q&^ц�z��=�AO���=��p���Yt/�{����5�M!5U�t]��=�����_�3n�n�J;�zQ�EH����8��6���"c�H��w	L�FZ����s�\��)N?�Oo�
���=UnS|���|�|	QM>lli� ~L���]�k��@*h5�q�g�(���3��� �$�֐D����V��@�TS�
|�4�3�t�21���#?pS�6Q�]��W�y�:ٔ����/����
`�C��9��
O�A���R�v���Pɱa΋'�"Չ�Q5�C�q4<����Ź�RSn�U�k�5����P�nU��L���C�R��r���O��8����9��{�o噙��	�5��V4ɦ,7���n'Cߌ�׆�&�uuw��y�h��<w ��h;Q�^��(]D)��ͦXm��ء����cuY.�D.
%j����x�3�ó�(�}�q���p��c_���c�,�2s�ܱ5�� �#�{�8!��q3Z�h_�W��e�\�ڸ ߹�ք� W�I^\<�\��&�|��1���Ef
��Q����h�aû���N�v�>�@��E�s� �iP9W��t�i�ɮ��IA���94�P���KG��\^�K��"�%
 ��zM�Α6�jR_� ���~��7ޜ�^; �^�e��9��ۙn���f�s��z�h1ŜeZ�fֲ�h:�l3�3��f�9-�#2&X
���G� �^�o�ֺ1�a=��^�
܇�x#.�����8��g(:���2�O�V�-���}"z>�t'"��������K�>���s`]-+J�ʘ�U��S�8��X�s��� M����~�X>��85ؿ@�Y�B�F�Rzڀ��K�����	ON�:ǹ��Z��8d�)�������D%yn��Z{�uc�N��򾻸��[>e�Y�B���!�SG������7��C�k.o�ꚼ4 ��d�u�纼9�t��W�p�Si�C�+����U�UY������K��gA���D�2�ޘho]�  ���3��(?��!�I�]gZ�R֕����/$q �=G��k�]���.���rk6�ԃ��*��hg
͂jv�`��v�:f��AINҕ���/μ�"Q�,����fQ;�L�$�r��z+b��O��ޮꈳBI.GOb>K���J��+�I:l����QnOZ�B�O�K-Q�d8�Ҵ�i��xѪV�y��*/$ˡ��?����)��y\�(R0p��X�-��BPI��z�5U	��ڍ�r( m6�C+	����F���X�X�ic2ȗ<��`��9#�ۏ&V�R����v�<ٝ ,U�~����Y&�U�F�O�ԝS\��3]�Y��7��zOĵ3�;xm6�g'>��8�WmI�ck��Efp�v>��.��.A��Pj���KV}�F.iv�炌0^[��GC?S]�-��O�e�����<��w	�C���0A�f�:�5Y8��|(?�:�2�#B�لm(��$�^?M�x{�-@��[�G(9�<4iF���-�%&G}�օ�
�S�s�e6��v˷�.ے����] �Y;�T��Xt��=A�U���`z�t�U͝ɠ�����R$��&�i7��oV��xB�L���h���7�^�XS"�t���&2��#oY�[��⡳��z�|�lG�T=E�� ���&���GV��^hԂU�7K+L��������z%3���1z�T�H�J�g��I�v�m[�9ž��;�W�i�ö]�h���� �J5��"��5��y�Q�ꖓ�V�)��\�ϼ�ݘ]I��;s�VKY���`(�$Q+��_�+�;�JaɄE�z��૧L�>r��6�c�L�ݸі�:�Tlb��IJB��2$g�v��D�&Ht	^��z�$�ӳ)T��Uyw��ŭ�5ǁ�L�Ͳw��
=���u�J^�U�)?�#5�9)-�C�{�oT���lx�Ȥ�P���&�>��r��� ����&��@�C�8�,V1�AV�p��Z�jj��v�uF0�y�5��8��d���Ĭl4\�Zy�5��'�(9�P=�ز�Qe�6�a(�1��|�GU���P��-Tk�!J�/5�7����{��X<�-�����Ը��bw/���"M�yJ�R�������pVe��	��7!D��}ާ$��($S���) \x��.�N���a��U`���p�h��S�(�ê��p�*�i����o͕�5��2�i��ڰh�ÚY��{l�s<q�揁�w(!��^݈P�@�DDԈD��3�5%��S�o�C	Պ��D��;:�e�j(�y��u�ņ����~'��{Z0��z�;H�.'J�A{�W��a��3P���a��O g��E�!�
B�]�4���$� F��W%��_`�dΕ��Xi����#[o�z�64-��*JS�|�<����x��rb��zm�R���Л��A��H��Ϳ��|�8SЈ���C�к�[�:�'x
��d49��ƧuG��ȕG��=܂�4�
�ED��t#����'�g�����V�,�Z2�����30x���d�tD�W�_`cԪ�Цᾦ7�I=%��jtG�Q�
�<^�����~�;M����ypY��u����ZU�P=�'x��gQ
尚���I�=)8��\��è�� l���Y>H��|�r
2���H�I�c[�����x`�[����g��n���a�*~,�Ps��;�-S�P,c$o
�]l3x;z���׾��O��C1�\�`k��T�8�3��:%u;�&�&��Ϫ1)�p��W�>h��hRn����Lҿ�H\o��j��1�w�����n��bE�����z�����8���5����� ���X�b>�7��I3p��"�b���|-hг�;W��.Hh%~@�~*�J�K��i���e��;�%�n~����DH��TO���U�+��rY(��<�jB_i׳�E�4�L�S��\�	�������t\��93TX�5�:犇�A�o��d��BH�sgb�Ĥr6b�+�Z!�8�w!�p����]� #�
[El��8��q���4�������[��/`̲����)j�!;���qҪ��)p����)n�ݳ��q�+��e�62��F�<��K��$��l�F%0Qs��Gb�Z	����W�7�`���n8#�N�w���w�aM��l��Fc�q,{鐛>� }���l���4�\gE"dh��z�1��Z��(H;��� �Ǎ)�%�[
�;��+�r"���n3��<CprwBc7�}c�ez�;�Դ���� \���ui���3�(�R%���b���>��������R��s	�.>˼��� S�f5q��p[c7xBK�4�曣kUs>,���]W��>��F��(mLM��#�W�ZW=x��2�:���EwTL1�!�Xې�7��|�����Z�8��W�ޭ�~��	Ai{�%Y��`l�MR���5�I�����BH���j-t<��}+I��g��<a*�`jGv��ć/�^݋r�o��D�
�z�9I��m;j{� ��u �6�]����R@3a�LC�YC'~�	]�R�3e���n��0��Ջ{5��q�U6r��u������5�=�ѫ�UKOb�������"�02�57�{��})F_WmH�5�S4��`�\4��c�������Oc\� �)m�O�n�-�+��I��8K�1lb*����������
�6vR�][H��c��Hb܁����p��9f�� f�f �Ӛ�og��1*��B8sD�4����H�t]���t�_ӵ�?R@��$�'I�!L��P �,��R
��n:!S�� ��S�A���mR�W	Sw�74*a@?�+	��e�rw������I�|H�	��b�>��?[���J�s������^�1�y
c�G:--��6HX��iۻhs�� �v�H7"�I�����?:��X*�/���ᖇ�d���"ـ�Z&}m�x�9�5��a/�"?��3��o���bn2�ٛ���E�=�T.�R��
�;NA$��1m[�����q�<�&�O��s���k�����t�R��h���oT�jJracnt^�KE�g�<"��`]���K?���&��wN�uD{�Z�7��dR �pķF �'�2�=e�w:��U"Rq^�6S��v��H��1��ߴ��5tn>YY��6���%D�1q��Y�V��U�ʹR�V*{���^�祜�������������:�ul�P���l@/��D��G�%�^b�$[��F�l���,P�����4{��Bf'7�7+����G�}S]���K�p�~�u\��'�&X^C�jD����ǂ���Š�].��l ��B��V�<��[�+Z����ȭ`ŊSo���!�'�: 0�:1�/ ���"��Nz�k,����<z��Q�=��^-�BT�G�k1(��Z��@���A����P[���˙ńr�����Ӧ&��[e�HUڍ=8@�_�7�0qT�G��/��Lz���Uu�b �d���(��`׃#[x��.�ߏA5�ɫ��A:q�&{��<y�olmE<[��A5H�w�k�,#y�]&�/b`��^��_�U��R`���AU��(b��1������F#KQ���5����P���a:�⇼"�U�wFXo���FE@.��ٗK�NC~Ph0��ф!�HA�<�T�78P�jj�X���/�m��R�n9 E���zm�}]=�;��d�Ѷ�8����\Ι�&K��C,]��ᩙ+��������9	�ެ�ֿ�(�pjoͻ02��{g-�x���>!Y(T)�v����6�nFn,��X��u�x�=&K}�F��dt�{�b+V}��
06c��\օ���&T���-R��YB�R�6����9%c�'�@E 4
,Y8���B������'"A�L��y���+�)*����?����l�Ľ5�S�SN:�d��� �S�wzS{�RH0'��kT �<���KO�-�,8�rF�L��euTi��6�/��c���3�rz^bBL�p��[u�/��D���moҹ0PX���[s��/tNM�v=-�*�x_2���_�-Է��V���N}��y����A�")��*�g�Q��I^-%�X���E"Ҫ,��3�ۣ=%i6���iH;z�G�.����!�^� �4`9�`�m�������
.YF�������_z ���a��i��l��_ ��D���F�|��唄��C�@��?8��uz��({m�l>�y������..�r:4��y��w�mnuq�J�pĚ��)x�p��SI@j���&����υ��}^8ń��7Ԟ���Q���	;=�o_R�bF]D��2Yi����?8����^Zέ��c�0��J$��Z�-��k�C�Wu5]!1B%8!����
�E8͖ -�c�c��2A� ���\��������X�^o�U^�tI�?Y*�6;c��DQ)�J�����c�Y�h|���;���J1�YKĒ����X�b��g$gq-����?��޺OJ�=�)L�[u� L�K�x���c�o��b��\8���������"
�I�^���S{l+��w��˥q�!_Ӫ���v�&���G���r�p���/��?�lԜ �P���K}�
������d����V�%&�ǭ�!誃7�<ƍ�hk���(t����3�_�\�IO<g��Wbƻ_e����K��_�0���R��DhԠm��Yv�q(B�U��=��ci�mt��?f)�M�/�YW���5���bz4�b[p{������W��,"`���uA�\eE�2�˚�34�yΛt�SF�K��#����z-e$��g�R�u���J	x5۫������ThA���ځ$E4-���1�u����w��Dю��;�d�X��+�,�QZ�"Ml�}M��m��eI���F��E�t��=��v��g��b�x/M���o�vՀ�κx�I^�A`F��I�� �;��6s9S����M�-Ƶ����xAKŲ ;
��o���E�	��_��ֱ?���{{�n��@d�����}M�1�G� ��K��)�c=cd��Yq�𬒈�2]^{){�z��q�}�AcS׌�3��->�k�D��s���`�'�Q�w���Ng~Bb�8�d#����/a"LBC��K��.����鰍>YF#��G@3�H�>����s-����?��et���Jh$.VO ��_�"�9�u����ю*��;z����[J5ȹU���}��%�������/��;=��o�	��lk����j�ی�)�̌٥��ɉ�:��!�hf�;k�$�3���>凅f�.���uL�徎cϔZ�l��� ����;J����(d׹8Z����ݮ�!&�J�}_b���}�O΁����E�f<�ᑒލ��!���=��4S�;����J,�`���h6�J�ĳ�<��_18;9�V6O�?.���~���F������bJv��q�^Er��|b �qW�zߵ$B�B��"�Z	��C�a\�=<��ͭ��X@�M�0g�wRm%r�$e����q��긺�ٞ��ӭNX�d��}t뻻���O7���A̵�؎Ԕ���Q�� ��p62�Z�J�u�"5�qI<j��Ѭ�K��)����D�>稞D"���"�`�?��f���g�գ"��m�s�Zf��˦)������Hh��،B�r�:�bn�z'��5$�:�O_{aٖ���p�企���gu�x�#���*�^�#j��:)�ty�{2�z�2I�ĝ�͉Q�%D�kr��5�65���j`g�S�	���/�p���i��UIQos-��rOm]拆�&�8����� r �2E5������`㾭�Z"������E�#78\!m�����-��0���	x7(��Q	��5%V��Ib�q�
/�-�@��P��8�i�ד����K4�l�T8=x�Jq�ɲ.s#�ee��5Z<�Q�۸5
OD΋��&~�E��YQ���K�4߿:�k�TI��٤�z�U-�up�u����m���s�s�[�nݶ;7���2���zԬ�BwQ�M��h�pW��r�ݯG¨�Q���C}P�u��g�-FK��>��3C	Z=�)aY��@�l���-�t,#>�3i�XPA'�VE�V蠥D���g�^�^�M��C��n��_�q~�Y�%j��`i��q�Q�az�`��.R��Ի6(�w�����'���nˈ1�ZV��v"	3X�-��5�0v��#WaVRP��.��#ߘ��D������2}	��F���{�D�:ܿ�����Ezi.0ݚ.E�%�>�W�`X�Nqɽ/���``Ua�0��t��&z���1{{�޹)ۖC�`��9n��Ol�b���)�OV��č+��OkO=�+k��ú�� -^A�%�TC�cBn��.8�3Ey֢��#y�nw=�Q�4�9	AgG��@�X��A��@�N2� ��ǘ�Q�lw#P{6�gg�X��h�_ob��\[���6 -�3>3�N3���R�����