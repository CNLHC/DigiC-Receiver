��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK�E2����Z*_:�����T�f���XY��G>�Ҫ�	��4V! ��9ql�5�T�=�Ħ�i�u=���ҭ��!�O�|0�}i����^<GWO+�W��]�x���%���P�#ZA�~T�H��}uF��O���Q�|���}PQ��X�p���.�C)V�,�ҝ,��ȍ����3��}�@���z ���f&����O_&:�Ë����;$*I溵Vџ_�Z��}.͝30�n (�2؏��]�C������|�i��6@,ǈ�>m�7_Fh�� `b����׿*{�,' �B�6YW�p����h��Q/H��W�|8#&B�������?��ªJl�xȦ��P��`���D�0_�]/��x'c��I���o�5�%oh�� 	���&���9�i<��~��`��])�N��-6r��U���~�Ԅ81��:V΢D]��^��`��c���[ʗ�5�Kƣ����K��a��Ǎ�99#�Ak:·�l:l�jc�L�SSyi�̌���*)o�c!yq0r]�A��;��`��FV�>���O��8��+g�J\��I��w̟K��"���:��wI��Վ�	�86X�JA��.H��
S6@$���q�뙖�FLG���m%�P1~�do�2���3A���Q�|�L���{3�u�T�F�lZ�%��|��ݏ�F�Z��ǻ�Ç/5�$�?�xSO<;;��r	�rB�}��K0��#�W��&Ϻc�a���=��0YW�9�(Z���m�Ր,g/?�����/���9�o\ߘ-jrr2�$������K� n<lk	�W8�k���a�>f�]L�B,���8v$	��<wbܵ���IJ+�|޽3���%1��_�X�����zQy]��ҩ���ќu@�M��k��c���&��I�e\,����-���+řH!]�A���F�c��Ȉv�քCx"�0���#��Ѵv
�YG�H���Fȭ�B��gʼ����	*��-c�/u!��M96"�����Ň0�*yt��0��Y<0NXڃ�7}��3���R9R�%�n;u���� �H�1�Yk���R7�k/Kȅ%��u�@��b�~��$�ZK�x,��v�7����Dg"������������?c,QS��st�O��Ek;H�0��a"�����Y��d���PG�CX��؝+4��2�����9G֍��J#�^���/�������H�Z�ga/U��l�(t,&Q��S����A'��AK�k���ߩ�x�pF��q���0#�0��,��m﮵kCk��),��* �\�� SR���C^P�ݪTy}A���.�P�C��N��'�#��{����#�6�D�>�d��xy��\R,*�@6E�C7%���8oo�GcpM̫�3��5B�e~�B����T��Cy=IH�N3�yEc�>����-�'�H��H���Y�����+V��kD:��L���'�� ��9�e�%o �K��rϳBN����G��b�)ތ�닡��d�A��v~��nH�wVQw��*���.,h�d�ۘz`��� ����5ϗ�)n���ử$����8��������G�����ޅ:Q.�u������O��#`4~=��}�Ե��z��Y��O>Y ��F��M�@���
q�����1�j�K1D��ƆYr�
AhV~�n�3�R@G���uS�Mkբ�!O2�.�tԨ���1�G�r�oo�JW�2B��ګ����߆�����1��ɤX'��}���K?E��r�����@�:��x��2��q��Hm5����G�h��������?�f�]@�Y�g7�Ę��nseSѪPw4p�j��#ȬRM�;&|�L2�%2�Q������ϥ��d�8�^�:�`��e��4s�W?8�Y���xN��y�J����l���ίꉟ�Y˅y�[�@k||�-ᾈ����3<�."�wuD�ד�#stcʛ�b���x4���خ �����\��� ����4��{�[n��%�Y�8I8�aT�E��_I���M �K�mA�g_�9�lYU�ei=S��.����m9@�3?�b�-F��q���s�A\�p��P�_�x���X6��myqF"�'�͐E�a7T�g��B�F����g��k�>B>K�NP!)_�%6����4�qu�;���� M�5��FOt�h��_������� b8+�oĈ{��/����U�CP��7,�}���Z���Ⱦ�)�L9uV�4��P�3F=�\�hT=��k>9�6�������S��_erc���'Xd��}�u�c<�.�㉴�x�<0z^/�V��F�U9��C�~�qX���2d���}�T�`���f��߄>s��9�BF����?��������H��b�#P�$l7�Qx ��U#��_V������Ծ���h3���jx�[���mY�Fdv?��"e��	S<�H�yAğ>�jW#�����at/���]1]c���4?f;�wr|�w��ȿn��&�%8Qr�+�eEؙ.[�Ӕk;�Q�z���N�:!�ʸ��(���]z��N-�Y�_��M�,�+E�^7��eѲ��XQ�C��t-޽��n�(����g�~�t&�~[����>wfԐ��C�.��T'������S�A�~踴�r� �ym������Qz�g|��R؞%���1[�V�/doZ�}��iʟ~tk.��v6��0)\p����kZ��
��,x��<{Z��F&���|���N4��|#���Y�G��<�0�dJZި�bC8�8�4wÏ��!��q���4xo��?<* Y��*�^"ܮ�m�rzF:�=���
�!�=S��W��-�$zN"��^1�r_��ߒ3џ1A�-��!�KF�ʭ�c��&�p�j��m�䢅K̾����1��#-[W�rk�P�Ľ)����#��ۨwOx��I/�8�"���/(�{�eZ��+�> rE[RI�a��U)۟Ѽ�5x|�N�6[{K�e�P�P�Y��5_���{����܌��b��ί�/�+4�cv��y�,TaW<�J������]�-��#摠n&����X�;ݠH�cc�8zq��f�?�ar� ��@���Fp�^K�[$����.��@�k��Z�tUэg��%���?"e�Q,g��mւs��{��;�%Ep��̭���X˼ӊ����l-O}�
V2��&�}�"V����/0����p���сDl� �a�t7Ns��e��>�=~X��w �*��+z(���3�o-��ɻAq}��&6!P��@�s/��Y�F���H����0��gE�}y�l��I�eY��tQ�E���e��Ĩh�^F���F�H��6oeο?E�}0EnL��[�2����J�tn{��'�� ����غ�w=��,�Ļ'�u67��Ry73v�G( �u]P�%�����z	�9�$��c��Re���m�;a���yq��c�R��z��Ld*�}�Q$��hА6�"q=7`��Ht�>v)󺿶@D�ɪp����jN,u�\؆�9{"h
��QݱO�h	t�
A�@M.��V X�����|��p�)�y�u�$l����ԉGIh��o�� ���(b��b���7��w����	��\G�8V2ZO��fU�����32|���#]1o{uY����{_W� P��2���{C��/p	<�c6Ns��Y��lSk�����v��F?�{o�ev@�4�g}=b2�[W$�Y[��l�ԝJ��5]�\�b{��G\0
�(��Ѳs1�9�!=?`� ,����c��F5��ӎ���U��vR6U����o��Xy�#`�R\`\��,�"H�;�N�%�S��*��zR.�R�AL����S��xW;�}��BgU��@��tfz/����|OY�����X�zM���zY�����m����G��L����Si�sS��"
� �}Ѿ�$L���۰�!4��htY��r���5���S #ߛ��s~�Qq->$r�� n��8�3B�|�.d�]~0}�!B�h�ݬ ��[2C>X����m:	��xvE{A�d0�0��v��T�ڲ�*�Z
m30�>���Ϣ�XQ�7�AZ��b�l~���숳���8��%��]���t�|D#�٣pN�e�oph�Pd�����4z��刴Q�Cf�נ@�pIxA:E�q�$m�|���=2���A:F����z18;P"m���y����.գ�QF�0Qoi�s
�Q��(����hq?�FG��ה�)�U��c>d�
?�Oi,�(�0���c�l#5`̨K��67����p�4kc:���3�5 S"%�hm?B���b��זm=~��%���)>DTO68�_�7�2�e�){��-�S���D�+�gq�!(f��x>�tk�\�0نj�M$����q��)V6O#z��Jē�<��}ys`�Ot����]�z�挶ik�"��3��B�K���,�s��I�F��~3E��)����ؗ�3�����/�Sz������3h+S`�.�{}��-�fG�;
$Pu�Q����Y���-�?�?�z�T^��8����̎\���@���7ܢ�B.7~���-�~��崙����:?b:��}%F�w=�[�Z+���esD ���g>x֣����YA[� cm��GXWv?���u��`�����Y`��h�Σȁ�Ny�N5m	�e���ȗƈ&�G��?OJ��U�1tE���y`L8G7�s�wo`�h�X�"Z�mo����4W�2�	4�"B·�m6��N��:[�g��W'럹���	������x�s4�~ ] }4A�',�\_��4�JtW�{Y�N�㜪��,|�|���M8���b��?G���ʽ�D=�Y��>B6��t��/�����sx��oW�8��e4��l�c�ݩ�;Q����8\�?!y���A�{=C��4��ڱF�_^�2T�� �
i�ee�_���<��#�@bWU^�Y�ّ�T5ǲ7��B�R���c)�(��ʬv�����w�释� S}"��t<����q�ʙ�ϵ{Y�,�������H��0��B0�l@��K��8�c�1���	i�B�oL��.���@dY�����<��n��Ɖk�L�<Y�F�3U{I;ӷQC(��"�o�24����kEC�/� �j�#j�o�N>�K+a_J�R�y��0�M��(����|0n0j����05N\�����]�]���_�'�_�I�w�m��:Yeen�ޕ ��ԇ�*bG�^^��@OCF�[Y~G)�:֕�D��s4�'7T0��8�s���}\��hg��w9JÊC�٠+b�6GQ��ծ:h�W�|�P�c����>��eqk����qz��l�h0�4�$u�� �� �zn���=��f�ب�M�R�Y��`B��U�y�YS<Y,�T0���*a*n�g�5�8����V�G6� ���A `��"v [b����8)�����,���m����q�	�6e^vr�d��PD9,��m�efv;���ݔ�^�����༙֓H�ߧX��I����~�H��l��&W^�AQ�9y��i/�JF쁛^p���t1[��~Tx�M4��}������1�:�'`"�K��]�=�[:��(毞�/(Ry�uBd�?�C���EpTٓXY��oGa�R5�o>r~��р��ҧE�5�O+�ZQ�T��Hڠ���f��s����9��V�lB�1NU��gh[�#����GN]3{-�<	r�ŨR��m�T�&Ϻڒ� _����t���v<|2a�|�A�],,3�B�����3�(�AT�~�~�I��u��KvI��%��!D�w�T���̵�#�/���!M$$Hr��ֲRQ<^�~�{��?���:)�qZ�woFv�:�x�z��.�{P����9�|�?��b��z�ca�9�X�	�3��'4)˝�(^����^�����"j����FO�1d'�;��.{��{�=o X֒���P�EW�Ͼ��t�g.	I��i�I>�����OC����@.�è��M>�ޚ.��Q)�Wj�9H�J��]�cB[E�v.�Ʉ���.jڴ[�5�(��-F�}�q�����C��cq��]�� J���R� ���ѫ
-R����v����k�v�htK����N1��[{'�D�
�y�F����Ho��T2�)С�S���J���/{ꏯ�c��p��Q��> Ύf
��U�M�����c�P��(�&��y��¦��B�l�u�b�lǔPe�-Ċ�)	�>�|s��R!N����,֮�:)�Q=�����%�c����ٚ	$z�J�ȗd��{�կ��D��>5D�ZS�W#l���I�g8����L���@d�œB��H�N����z,t�r�R4��;������"i�1 z�S�r�?���.8����_�3.���;0R��}3o��-��
��Г��EN��j��
��<���2�Uaa�z�pUB�/K~��6m�ɺd� ���CL������3*Fσ8ƌ$ے��O����k�K�4��\$��Z~j[U
0��@�]"m�WB�Ae�GW1�;���Pm&2bE0�%�l�@q��O	$�ݽ�,T�FnY� D��Y�%[���(�S�Ǽ:Cy	>r���j��B�<�ivǱ&?F���K�G=�6��7�Ԋ�,��v�du�M��l���@�Y���Y�f�1�(��YK��WhRB|�>l��-��c��&���nˁ)��U>��`���}�����	�~�hOPΆ�1�Q�`�l���4�V���z���P�N��8s���6�y�{(��`��Q���Z��H��Y"yN�u�r%���̢K�C^��O[=U��95j� ��ș�w|b9�k�Yt`c+Ɇ��m�MJ-�p	@�^�/�܏Ԫl�u�>s���Ѿ7�~��"xF���u�03�y�;Rm@Q$ܱDA³�w㊯9<^+,�&���$!�a�0��?�qە(x�ݷG�NJ�h�^M77v�a��M�2�GE_�	�pE���T�.�#m�����9���\Ghw-��&�=B���6t��=n�����!�a����!e7�-�2�. 8A�* ����V����m�]��0]��^m�{Ց�W�A��}�I�,���!�1�����༙a�s"���\}Ssj�����߹&oE��M����-��Ү��/k��)�W$���M	H���@z���ë��{�Ê�ڣ���G�Z7b`��pBc���t@��V/cǑ|_<����Y�=^:�)Zj��<��:�A��@7Jbs��ɂg'�|�^�Ph�A�EF?�rp���@��o|)�}�� ED_ƒ�7�"a�(e2}�;]�?=o�",����\΃��8�Sk�Ros�~gcL�9��/���?̂�{�.˞��ؔ�ٜ��=fӯ2Mo�ox�䆛;�|��'t��D9�BZЍ�����؈��?hTL:Rڐ�/|YJ����:������OdtL߮�1����4h��q5o���|w05��~��~��|���O��S�g9����t& ��a�;*�������VM�F�'�f��#jMc�h���Z'TU�=fm��H����P�+Li\���ԓ��sq,����Mh�ׄ�[9
6��Р&�+Z�_ARc|����m� �#.���z�ʨ|�wjVZ�_�{nU�_��Ďs���L`�*�=��?����UdT�����{d�fi���d�;2s�yr��ˢ:�g����2x�x&�� -����S L	w�rS���ص���r6(�>�M=���^~/���_�o����!�轟fژ93��;��W/6����6P︐l� ��[dy�q�y�*5��?戋�%[�Su����0�O��a)�s�I��S2�O�����jJ����[d�x,���4%��3�Y����Ioo���9Y�o�";N�PL$�|�ؠ �~Z`9�U��:-D�d�#`]�����\SPG���7AAK44���Y�O.Qk/б��I�*���d�]��w[1�6��D����md��W�p����"�$]r0:�5ԝQA�Dh�לȣ/K�l�&�'�q4�O��G�}nyv/�n�T��U�ۋQ\��i�X,��d{�ۮ'���5��Kڼ94�l�WT$�K8�_���� �������] �U`.s���5��J��E��)F,��_���ǫ��i$@�Q�ÿ�G��1e
Qo�%�k�&´�xT�5['>; BK4� v�_�:C��<�Q���OZ��W�j��~��P�����w���ށ�-6�Od����˭!ni,"d���WW"���yN�f��;E �~/�"V�[5B�H�b�=��R��-�=7`��<K�hO��դ\|B�w&?H�*��О_��F��YbZӮBha/�S�Jh���Δe�ӗ\�U7��;�� ����D'�Z��4P@�߉�/�~���	�����t�w��������i�otk�c��!�զ*�<��vJB�P|�~At�f�T�Cr��.�9�Cw��u����_��z~쬤��J��O;A�h�1\��M����H;���}�:���*[x+ ѽ�k+���PP�Ec��R{���d&n����%�gU=>d�Z�ƿ��Z G������и'�_��U��)sQ�ۙejJ՜�$��Ŷ<�&�fMM
��Q���^:(��=��`�e]����X)��<N��A���Q�X��.���fDa�^�X{�����*҃f6,�/.�ΰB�U�da����?J���kz� �GԾX��YYd�|1�Eu�1�b��dG ��@1I��Iފ^d(�"�ڼ��v)��y=���0܎���PвrF2��,SG"�5#'㒁Rh�'�w�hC��=�`�!IN�P��Y��̺h76���ٷ��H��i��S�7q@<���˂��<�6V����Kx���R���*�JDf��fP�Vp��m�$u	>�����9U�22��,�o�y qepH1S#K������Z�,�t��m���!B����:X�7$d̠���Pݮ���J���҇<�g��Br~��Sy��{;��;ǒL��sK��&n�_�)l�䀎;�@�R��xq/Z�JH�ئʳ��)�:�!Z�|p�r�̬ʹ�}���"�b������5g2���X��d�h.�sN`��Е<��y-Ӄxd��۱#��E�B��Ϳ=w>�	��N�c�j�U&A��JG�6�P[�ֆZ��q��u�*��J���,( f;;C�7��_�������e������5d<�g�`�J�ǀvx���J�w��9��@(p��-yc"�Ƣ]	���	����hߖ��.~%��
���fU��he���?�8�"=���N��7��{�R(v�6��zX�f���AL6���2�g�`�E��ǖ>�ZY�|Ѐ�҈0_��IOh���A�����wCM������Y���>��Y�vOnВJ.�i�3���32�}�)�E����CC"G�?��r&6�ힹ��}re��~�n�H�������uI0�fX��c���{�� ������N:�1�7�;��O��	��o_�K�&��ꦁo�G+��G�3]�NmMT��Y�ݢ@�$<͉���v]Ĩ���eS�ȧ�?�v΅̈́	��B�������x`x�W���zΛ!'w�����3�:�-o��y���?t��t�<�H,^[�|���郜1���
�9��w<Č��O4V	hUo���I�$S(�tttqP�Z��t����'�1l�J��E�p5i��E���Q��z$SM���OW=˿�w��[��u3u ��Z� �q9�L�z�o��̯����:�Z�*IM��f5H��� 	��s�:�JϏN��&�>�-�u�y���%��^"�ʻ�Q���8r����2HYc8Z�(	�{��-���T�Y���%��d��F�\��=��m��2@����{�7�vN���t�(����QI^�ވ�e����OO����<y%g�@����s5RS?�R������(��lΏ4˳�;��.G���]J��z�� _.�%m|F���`er�9�e��? r
"��^~D�qv�
�5�T��:�q,X��?�Ok�����1-��#FŞ�<G��w����W����T������Y�\�~�F�o�=�h�]	f�BR��އ��+��&�����P�gϽ��Bڸ�3�JI^Fw �[��n0u�;�JRҹ�gF�~sN�f�],Rj"͡P��ʋvM���<�2�3�c�uD��s��P(q�X�";Y���1�����A�Ԙ"b�`Qa���,�7f��uK�a��
%S����/詩㢭(� ]�N��*U�PXn��P�(g��V���.�Y�j9���wn������~ڮ��E��M9M���v��0�忺�Pܩ�Ҝݎ��z	���ʔF)��D�5�[A�G� ���� 1�T��R9�6����
���>���Ë�����nh��ǍfI&�Dg@��QdeviH��vu��JG/a�|�5�R�a�%l�/�:X��"m�QDB���q�q��ңz\�-D���h���'�� ��p��q���SqЪ��9I�CWzr�髴#����<��u�w?b�S�����!E��i�	�;�B�b<�7ȡY����m�F����'����%���?0+/4�3j�4��͊�o�˟%;Z�"�7�_�:A}����޽V�ʬG�c+G�:����?.�{���0/;l;]ou]�2�ɼ~��O��v=�A܄�vLg��r����=����/�u��$�9���83�z�Wx �D�VYֹ��X9;�\��q�%IQ��f�;�������m��	��nݰ���q�ԙQ�,��qi�O�d�D�{�M�È�����g�e��"e�#�ȪL�����ng��ƽ jF�����T�E����瀂�#J�VIr�O��?���`�6F9�^��y��\���tGM���7hTA�Eit�E u_T�WO��n���`�4u�����h��*��\�p��7u@A}'��i��%!Z6ί:�rK@�M���F��jY�!���	�k.����`�Z�@z�h�A��$ {��WybCYJE���Y�b�Y!�E'$1�����.'k�c8u��L��b�9�@o���`ًzm�S�!	��OE0��ҾA�O`�2�:��!��C�"��8y��.S����Q4z�R��dIe�l~9ͥ�؈���ahH��F��G'Jg������<jW3�I�Æ���g�*���Ǜ�ײW��� �������QS��:ώ�`�^/`��7�y�m�Wxu����I�h��Y�hy���k�_�*0����
#�����U\7�Wkяۀ%įG�4�A�ޒ2Z��OW��)����,���}����z�;+`�;���j�v`�L,Ͽ\9��\@�-���b�&� ά���(�c��V�\+'ui1o�5�Xb��%������,������3�^�ۦ��	�wS�knMK#�|G�s�$끒���sJ��V�*-{��U��5��2����E�@���w��A�Y^7��(u!n&��#��k6���d�g����g#AC�H������U� �3#��d(H�LL��6TG*���6X��\T��j#�!8����f:�	�<'�Ih�f�8�[��k��}��I���b��VU1@�a��"�^RzAn���T�iPƻ��R�WuF�nc�&�Gy���nospة�� f��?�۶��} Wȅ͹f&{4�����i㋞i�b]�+.�)�6+�����S�i�WMX����&5m[��D�])}&hbZD�i�櫸��-���f� )l�(��9>e����B�@е�w>=��.��\���?����*����})�� ���%ԁ%�5���q뱸�9�~��g'��CHT�Q{J	��Y�N�ٔ�N�G��\����J�Ϫ��VGAj��b`*&���3?�'�z�a�N��XȻ�ζ��g՚nw1Уac�0E��a�͗���Y|��
�rl��i`z�D����Uէ��V�mÕn~�s3j���Ip8A�Z��8�U;>�* �l��ʝ�C���+
M!`���=<�b��B_4`��Z�.��E-ZX��0ޛ�b0�C�XY����L�cU�m&��1��|��F��3�V���q��_H�2�i�?�<�0M�>�	c�q*|wy\���%H����F&�e̾�m�e�����0��2mx��iOe�~�&�� a@ؑW?X����)���k/*��!�u���O��K�/�t ���[�ݕ��������m���Rq�hJ���[Y��T�|�r�֎m���+hZ�o8T�0s�Rc�"�j&�,σG/�KE&�����7h���E��(Atd���ٚi`�˧�?�	��
ҵ��6�����Z�pr�;�}Y��+��.E�~v\�8+g����u�?٦O7a/�Jt�8�I����˳hT���{A�H�[�t�)r���cW	���h3�F�65�x-�L�w+�4aMs��5��̼�=��d��kg���a\���t�0���+�h���<����΁D|d�e�j���@�z�Q���R���62��k��X4Q��Yw�$��W��i�_��2IK1�ˊ(VLn�q�2E!�g��DP�$�2���P�_|$ <�6GE.�nK�%�$.�M�	�M�7/ۭ��@;�ЧYN����/4�B��D=����,�������Ku�I�"�����I�y>����aOj��	�F���N�ҹ�Ou(`?�܉��f��AVd6�A� B�+�c�(����l�/�E̷�z��[EA�N��E�Uy�HȐ��q|�;�V�Z>���\�<��D�C4�s6���Sj}=v��6/���r�|B� ��q�1/�z%|�w�ze[w@X���m���c�Ѿ~�B2��Z�jp�h���o �`��P^���<��QYGiw�N�s��p�~�P�����M2v~t:��}��C��:��[,e�3b�兩{��dJ�b�������}��J����&y'�;Y�y�xE��]u��Z��	!�6���B���Ɋb1~GH	D��ͣ��0�Qn�̴3	��5S���?�}�k��Ll\�
�`'���t����$�1`h��ѝ�88J�����)���DǬ�c��{y�@+��J�/��0������A�=�=�G�w%�
�ƙ�Y��,,�>��XfH��^���Fu�GTSP��FF��4�� ��d�����N��ɚj���8��v��>�4;�ʇF�[ y=c$C��/3*����\�th0��*y��&qo2jw�ש���d<Q={��O2p�k~����v"<P�3��H� ���.*�`x���YWP��ҳ�g���R`q������LE+ W'��	�`�νJ�q�1���s�l�a�^�n�}c^ �@�x�a(		��H�f�W�����'9I��S/��P�TJڅ"`i�~�[�7����x���ǝ��	&U-�#*�A���sկ��wY��٫M�y���ȗ�������Hx�s&�Pg���Л?/��@�R�"QW]q�����J�zC��2Xq���U���������h ���I}�-.����~���:��8���*�ѕ������	r#�}�����G�4������yd뢈.�÷I���}&�3�!ѐ�E�ִ�V	�P�$��GG������)�wy�L�Rp/(Ƭ��:u��Tj�@tRX�L$Fr��^+��ݶ�;ޟ�{]e'$���3�;��<�e���\�U�B{c��!�Z5��g,1���k�]��5�I������{�~������erPg�	�y��b��ۖ)Ȩ�[@}�a��r�䨓'K�kLo�O´u�|�K�A���ד~ϥm��gj7-�#�D���%�Jᱯ�t�K1�����F�5|u=����1��l�s��#����q��ӊf�ٮ�@+�Y)�46ҕ��x]>�(-����:Ym�Q�F	���v�է�(���\5C��A@�X��Tˆ�\v��Znn��Ar]nD�u��G��������ŀ/��kGI�T�1<�6�9:��)31�w�N����䗰ߗ�;z����p��0����gS�`���
�U�k�#*��ӜM�J|���XI���׾.c���]	+��/�Gb�@4������{�Uo�%/=�5�q:L?��2���;W���!�l�Wj1+q�R=��ռb
�[�	9��G���m:�;�`�J��&�����+��L2��.3���ؓ�T~�d���E�B��/�,׭|���H��
.�B��������=x>�XIf�+��Q��%�9��3Pb�;a�^��;����QSNL8��k���+U0m6{�����F��7a��W:���8��L�)����Ws����Mj�z|�b=,��y҂JiN������n��&X�2E�{nܹ���Ov����17��%|k���+��"����_������׫��M�f�c�jQ���Q��E"E��u/~��[���p{R�0Pr�.���7����wQ>�aQ�����:�^�HW9FR^}<0��1�6�W��28{RӟZ��I'ʯ�W��,�Nw�"q�u� 7�V��hU�	Z
Pg���"C��i�����г�Y�� ��e���-��.�h��k"j��b0��@2����������~�5�1D�����ܕ�DT�0���;6[l��; �^(�y�i �ɾ4f�������BK��XN�R�Uv��0^I V:�,�CǱ餐�7U���k���5����:E�۔S�^�f����{o�S��2oOq�ԇ�Ʀp��p�X/�k�N�rfֿ2�"O�nw�(�-�J����*8�h���O��^ -; ߷<�w�fێQn�V~����2�����mʹ;��扯�_����H�V���< �s�_��fw�Gf�>:��(�ڕ>I�1��C���&M��bל�1%�*�:�Oό����B�J�榌e�Ghcq.O�c7z�,��ż��݌��9�-��q��$�{ǭ,~D�0R4�/[����G���̜X�. �Q�^=���ɧ:5�Y���5��恮����J0[��N�����*�V�-���~~-r�*$��%�Q��G�=�m�ɳ��iw���O)���'_��z�C�4ms����Dp�ވ�h�|����bd HUw���������4��jZ�R�t�M:��'j(����giZ�X�$�;��l�+��)$�ͱu�37���h�r_a���9�(���4&����_B����Ed@�K�J�z���B�1>��>p3�`��^Nz�s��f8�)&���مuh�^)s�Z�xlG���2�Vm�U��!����ᚴx�L2������1��O�^�-���հ��%��Uu�|;�zA|X|��|������gY%@��i��]gb��C�R,��E.�
х26R��G. �FWP���f�xNա�Z���+tU�1�N�bgD�L�y���b[%��X�`y���^1��]/�-�2I,�	ӜS��,|k"E������A��<鹞��
#��4T+�t��HX�=sG�r5#�� ��h
dQ��>ң�G��]�j� $�([����hƺGؓ&C�@������:9�Փ�y�1��_����q@ՁP�쀜�T~�z�#��IH�cS��(��@�Z$�a�
�A���<Q�C+'܏�Q$�|����8����93��_�?=��
 �����aC��c��ܣ�S�]N�^��2F7+F��SI�T0�� �D͗���{s�X2�;�-j�^����
?�b⡫��{m=��gw���*W�F+��zcv�[g�n�RŖ�n.Ԗ�C�m,�l`�r�ц@�؟��D��[�5˙��HX����/�z3��?7.�/,|QU��Z�)8�*�9c���	�Y����/Z�3��g#�������\]R���bl��+���8��Y�F����"�F�o�����{�$�[0���;m@$i@�#�C$�<B�[��h�X#����N�^	��v�y��J�� ᖪ�c.��ҫ~��ߑ�pu܆:[8� ^Y0�Bs��1���ݟa�����y8�*�cQ��\�[���aǝ�D�O"mU��7��Y|�㈼�6����Q�o�7�,�<k�}�r@��ȇ���w��v�N��$F�ze��k~s���%���,��p�P �����ŉ���D���^wL�}n���c7���V����4"�&��qd�*��3tJR���3�`�P�I�,���6d�#ϓ���i#)�p�a�#��<���3��o���;�,��Ŷ��kAεG�]�a�� ���Ć�c����p�\��!f<��[�������.2�"=�Um��G�Su �b�u���(���uz��W��������7�lr3a#�8<!�/rg B�;;g�T��+&?�a�'�	��6� q��kByo�o*=��P=��������`�&��r%��M��_�i�������(���Էn5�\g��{e8a��0ۛf���o N�>ȝ�Xk���O��>ʝ�5椝} �!�<�{&z��Z&�(�[�	�>��ӭ���b���.�_	�{V��Xux�f�Qv�޼W��O�����ڴ�kzx���E	��_nq�>�ybY�_� ��>Z����e�)*����:���@R[�H��:�^k��9�5�>�D�6��k��@�ˆ`߲�y���!���s@!�6\I,/��&"|(���_�:�8��F1+�y�1��@e����v��:rƥ�K�����n��ł�X�#a��{0��,d�������f�Y񕎀������X�Zh5�ff5P���_�#��2�v�O�0��]�O���	�E������C�yow$RP�K�W~�i3���>�%\��wr�Pw��|�����`�^ۃ�쓒���s2^���!ݐ�Tn�ΐ�~����zB(�R?I"�a4��n��v��F;���䬏.i>��{�CÁ�U��L�j}�+$Ҥ�G���x������eP{�����TC�'��NX��Ihd���Vx����I��H�+�gO`u}f�����.�uifh!��1�}\6y@[}�D�d�pqN@�Ƿ���SFT�!%h��� mg�4^o����a���k�Q��7ϐD: @�)0��$Q�,W��p�	����%�$�Tv���69�-�YL�I�M�f��	?�d�ǝ��x�!,��"��������k���EXU�C��5_��7�V�\.�xc`.�:  :f[P�SEͱ�y�P�vB�\�X�bR���S<T]vhJ6�E�X��<<4��o����&+��_���y�����KO�[�Bs����s��ߛ��F�#�A�� |���������]4�BS����qo<��׍�|s��!>�Z!�Z�A�Z�l:ꁪ!��D�c3���ƞ�H��&Cs�"*�R@ �Pyv ��?��`�ۀ	nSK��>��+iu۾�z��O��M@P;�9�7(x�H�kҵ�y�t��$�تΈ������`;q
ߵŭ��@*٣��X���{*��Ӯ��l�ʈq�PW��ߙN�������@�Y.f��vu+�� ��{��-�f�:�A�X�X6�I�
��X�&;S�o�$�KO B�g�"���������	�B�+n��v-QF���{�d��k����n{�;�6���Z�imߜ]�$����I��/~��'QO]\���/.�	a����ýq;��{@^0�-�O��@�JC�
�Z���
����7���wD��ˉ�]�#Z��yS���_[�|U�������P�.��}}�8�������B!��-><1F��</�ѲB��O��0�7��f��[^:�"�;7ZrJK)oͩ�;�����[�"�\�I{,T+�o.?wu4u1�~(.O�Zl*�gu�e���.�;�I��gvV��Q���]��/X����%|�Z�6	���.�cL�����Z�2o�;X@%���w�^����d>MB�a`��3��+�;k��O9"�ɋ�g����z�ܻ[U�%"�ŭ���&C
�%ߜ�����ܱ�)`���;��:Pf�r�c�d����:^�wT�d5�X�˱��8�����K$�أ�?�z@�]�-�$�v_���2����[9�c.���r�ӆSZ���!�i�3.�/G�!�o7��)���M� Kߗ��ց������i����0- 4tXH=#+��!�^Kf2����Ǹ����1B̡�@k�=@�Ey�����%ޣhA��Q��,p�T�;jϋ�%fB�m��(��q�NLx/�Q��m<@F��P���-�4UW�wklc��J��X����_��Z䔣ZN���R����&^�^��+��7A��I�)�u�1���/T��Sf�����7�>(��Q&��� �/����Z�V�vw ��F�Au�.������� {?�����5{���ϒ�qWS�#[��FL�|,"(�o,V_Tce#��k3Y��ơjh'���{,��kT� )\�;��Og����Z��5IN|4��t�D%Qeq �����W�t��C�7��U/?5�V���!t��D�G�Z�o⒫+Ɵ]A�J����犁�l[@�������D��;f2:���˟��2@y��(�U��NZ8;p���>� �q�X�tb��k>����),BS�A��܈�_	M[=�Dk(�10�fJ6��n|�
�h�z�l�Y��dq�})`睊}�q]lE��gT�f�������`1�v��] �[isr	�y1�b?�@�a��
`ڊ�����%�"��1�'Z�w�*�>�?�
�r0�%<Α����=���p
{�-���z�;['sWK5O��>�%9���Yh�W�R����٨�ĚY[�|�D_�^@���7�wsr�iROŹ>}j ?�Ǆ'v��E�t��,�]��&"à��.�5C<�\j.��4�HF*�۾�_���N��	<��ڳ]��-H��N>����J��ۻK�oM1��+6՘�/<�>�X*8M8�zf2휐G��O�l����L0�T����w�7��	Y2:T��V$�YH��v����vd�.¤#���V'>�r��=�,���&(��2� B�4�^+�΂�	��o|(o}�kܲ�C���}ƆӦ���=:�~�5�4s�NB�T�㡲�M�v*I����C�{��	�:�#VU�dƶ��W�d�L���9]I�E��c��<�{���l^� �5�\<������c?�8{��EaP k���W�1Z[�0^�^,ւ�x�l�ǘ��I�C ���c�r����s��Д�i��4FJ�=k���������$i�aZd��=�������t�摒�m�խw���[�B׷\KG��>�8��7s��=`�s"��B����Z�=������R6����r$8��	�_z_�n:�(u�C{��S�5aҋ�S,��^�g��	���J��� P,_͓�iT[k�>PO�A����K+����	�y�E!gF#�A��m���*N�9�}�ࠟWU�X�v(�5��%x��v���td����~��4�)� �خb��Y�G�eLdNd��RT���ۍ*�r_X�����.j�9��e�P��7�zeFl����[���t��J�q�B���fu��Sc�BCz�5�ɾb�/�.�S������ֻ	���)��	"�r�UЎ��B�y��l��|w'vPy��K��D;�0EBl�t���3�d�
�#�4o�߻����C����v�fJ��:#��e��%��g��Mr���ē͠���ip�TG�Y����Beɍ�MA�|l���w���%U&�c�3��x�HD.iZ�ʸ�Uco�^�;����,t���-�x�W+��e>�ƈsL׾���ڢ��`,~��\o��­:�e2	����k����W��
	�\�rI�0���Ԩ�����E0"9͖�@3�1�8_F������k3��S[ `����]�V��\�!��j���^��S��`����<UлML�3NeV�vv����N"����qt����xz�ιk�ߏ�&���7��0U�d�#�_�>��� ]?O
E��
u�M�^�_*37�B_Fm%��ɾ ����0���}�>
j���2�*t�n5����MA�?�K+@�+w�s|�*�l�G1����(���?���
�������h��� �+���Y�����+ԁ���ȂcPy�f��λ{}mxV��
 ���D�j�~���)�� ��%�;��D��2���V�v;�7�@vut���T�b�M �c��>BH}U��w�Z�EG��cN4���!�~--�[1h,R��>��KP5o��i%,��ѯ�u�� d�ҳX�����1
@�|N?��*�|�����\;^T������c���<�^v�U��(�K��.o�S�5��8j���힉Yw�Mt�6��֥꼚��2Rr膉?�Z�A��p��Ue�څ����+N�J�����J���$�5]V%H\7�s��nЉI'�íBOC�?1���_(��޼>���Xh��wK��E��ٳ�̮e�r�C�+�}���`,t�
Z�	�YI�<v�o$�E�	�	��=V����u_6��\�#��t������2,��>�=>�6̓��!�ڑM���Å����E�I�����Ƙǽr�a����]&�$dǃNy�h<����8<nI{k@���j���b~�su{�]nH�=�w���J�a��P�&ĵ(��b��~tWT�E��v�O ����D*���M������E(�p~���bd�V;,� �/H�`�ێ�b��͢��CD%�냒�����c��U�NF��0��PR�Y{Q�bCR�`��!�)�(�W4~Zwr�����Ħ�1�ӹ�<���o�C��1Ё2Y�v�a&Ac9\�_=��X�{�	�bo�Ì�|G"��!���oa�ܛX���j��}@&TܿU�����6{���?�
D�Y.�=�h��(�p�Xu]�yQ������$�(�Ww�<3ci�U.AK��_�W���_��(t�^0�����Ӈ�����h��'���͞glc1����,�g�|�.m 	� �p�p�_�!I#�+�AE�9��8��4�����c���T��T����.�=[N	�h�����˹ǔ+,~�KP���.�	��UO�
��G�/�v%W����}���㭊����;���\�ި���� A;udf�v��­`�[N��ҥ��D�u-�s8���#W�h�ҟ#��� �cv��:=-&rm�8r��P��X�O(��ԛ۱���)[_����(<��~�5ǖ���$���X�ש��"ueS��J�
�n��?(V�^ ��RGo ���5T[(Xʔb��0P����G�/ǲb㪗��Vy�7�+��(���j4L�f5��Cmʯ�)#�����}F�O�/��Z��j�Q6D�;ڶL Ye�,����*`�L!�i)*�T"����>������V�^X�[ّ��ޅ&$�iK$ܨ���te������ �<[Z,k48�0a@�ܷ���H~]�c�1��U�v��,A2������~�A��z�G�#�����"5I���AQ�����A�Q��ka~	IA�[�.��PbCNUl}�e5�>h�\W��0 H�x��d���n���V[����Z�@����7�oL�Yp��!�قuq��D!D�Ю��k}�2��bmJ\�b��uV�����_߳7���SO��FÓ��]��"C�4N"�d(��߾>(�w��R���uRs%��q�!��V�=��L�����ڡ9�⺈"�Vw��(����tP\Z�~���P"�U�"(5U�vG� ��
�a4=F�A�:!S"�Yb��k$�����t ��<��@�e���s&�����W���P%���n?�,�`嬅�>�Q�2���G��B��L�N{ ��V�)�PP�Klܢ�m`�_!�YnIJ�,"F�Q�YD𕫔��?O�J�+=��=Y��+���U^f�S���ENk�f#6~I;�e>*��� ,y��!��<u����PnLFonB��Zll5�H��f��~[�$�C�o�@?@H�ro���%������7��{����f1x�n�~��8���Δ�x���&���Od��ݓ����̷�w� ]Zo�cK@czt�X�X���^�{�pC�W�U�14��4��Ƃ��`��ڃ��Y�����;�v�� �f�4�e<Pq��˺@�]��yz� M��G�F����}1�wv��tz�5�V�j�Gf=V�+&���2{a36C�Mx)�l'r���/�C��p�~�,�u��A�v��h- �EU��bWB@�u��?���w#?�k��U��i�{2S�7Z_?}��;��"��.YL���x����׳�W?͙��܂�mجl��wH�<S�H��3�z1z�����<��M;�tU�`�@��Ѡ	�tL��{�t~Ǻ{�ŧ��S�:R����C�0��ch��u%��t��C �;�WA�n+�O��k�	���;&s�]�P�P�.����L��J(��p�h�S����0B;��e�z�;S��ps�[/	P=E7K��L�����i��#��W�iG��f�;�&������1�z�쬢OX�b�Ss��+_�9��]sS����ap�ң3F���,,k>�9,��{IRK�J��6!]������&(�������D��<���.�Z7ꇘ�|�)X� G����c��2 ���iڪi��ﾚ�9� D8H~feo��wC�PDٙJd�)0��T=w�Q��=�2�b��7"G��"/\6�c��|�c�u&@���9��)�%�%qa�^�ׯ��!i�q>����9�r�F��TI�?ZƕJ�������;z!\�4�ڋƘ����W������:�J�G��kAM;��9�A��R�R�)zV(b�@8&Ƴp��uo�p�l������^���&h��Q�׬C!�E��g���07��������Tۧ�{�3���kd&}sd���z��ۍ�[���YR���.�xLˤ�Φ"�t5�F9�q�r��Ux���.Ԝ��=��]����o����^����+�8�!��~�Gk*ݬ�N1�%�ǅ9�E>-�:��v��<�vA���N�����N6�n�_w�FbZU�C���T~�45��q��	��MZV���؁�Jh�T쑮Z�����w/�%��.�WF�s{���� b� �it���\��╶���|w�oL����vw�jm�K�lg�j:On�T2k�;�"d��ޗm�1�yY�i��/T���q����h��Û#a���p��l�h�d���?ѳ��K��e�q
l>��I�L7qv�N^�u�W�k��	�C9�+V�NU�6,�{�̇��,��Q�iTk���_���;��A$����N�- �M߲4#<����wgP�]�bQ)v��\q�&���������}O�U6	���)�8'_�φj� ���	m��[=m�AI��{�?��$��[����FެW^7�ļ�*��o8-� �!�,�,���x��ڕ�K�"f0��/�u�D����]���-�p��ﶤ�?�u-뒾pN���r�,=�x+�(�4\�E���M��n���L��n�)��*X�'�Csj�������o4��19�<��1��1�6������:�ªs������>>J�8�_�p��j��_We1r�䨣��%�Ъ0hX�	7��.�_Z��_<�Ix���=&MN�F�v]ئ���"�����^�Չ|�J���@#��W;O�VE}"�&��
VԖhm�(T�A�����<���֖�^w+)����@�zcڟ��?�f��eaz��C��|'������LU��=�t }��Ӆ��:p����s�'��f#[Ʌ��8�����<ee��l�m��yy�)��t�#h3��<�@��ݧ��JF!*�Ѱ�J�Wq���6y���OP��#vB;�=� �z�h�dm���}�TW�s�;�B��X��%������}A�[�8���*�~�W?c�
nVt�a�n@������2)�ǽ�T���#	�n�<��o�ӗ���Tu��O})V�F6�{������B ��Y��:����u����O�y���� �p��s�� Z�c��ٿ����Jz��@,'��4�$��3�%��¬Mq���8�@�:@���f�RJJ��?K3<�>,�����~�8nK�e^qEx��g��~G�ŀuLĩ �ӂ���Rg0���K��x~|��X'u�w}Ӝ&dX�5K�!��F����?1J��8�A�'�ѐL��O2��0����5�mA�f^*���5����G神%��E�����O8�ǆ6uN���!��#x�Ø"<� )�,����Fd�:�>�5H<��� zq�����c�@�'2�;C���樣�H�����h���� (p�3�W���т�b���A�S��#Rw �s4����D� /ߒ��{=�neY��k�)G��O�p�v6ˌ�wcM�-*(a�1�Qp�p)a�u��*���{MûA�޻����3@'a���l|��9r���g=�^l&\�1�%6"�Lg�䈚�D�\!F��MF<�Q��3��������;��q�� �~"�睮���a���9��qTq(P�5��t�y���U���~��8���E��L0�|�ʴMR�m���,����Jb�/9E�9���氾�)����ka�ƶ6�Ӡ�z��E35_���g���U/5��76��}�ر��I�Z~�$R�-���*OIQ���ҟ�� s	������d腆��[�;j٧�z�q5G�4�S�/㗠!�>JwJ�������z_���3�G�"}����nFe�%[��Re�0��)��S&�<���A���k��Sk�7yQP��9K�)G4Y��*�'R�ҁ�e���a��}�3��q��-HTt�����~=��C���(u����N�W�~Erj�xJ	�u��(���V�ٮ��}���W{���e_�<��M���^�if�o�n�%�0�3����L̊ �RZ�|�)O��#9���ն�A8.�X���,r{�?L^�������W���<��؇�y����Dz� ��?�V"���3]Z���*8��Q�އ_�Z��U2]c�\�[�m�{�z��x�ܸ�6M��|�'�t��;�P!�T��I�n�K�T��#&_�Ս.i3΀��'�����Z�w�=�hD_��S�wk3������?O���v�ܸK�)'Ʒ��Q�8�!�W/:�0���"Sp����<�T�}3�tU�^�M'(퀂}�d�qx~�ܸD��B�J����l�8^V*�_��~zo�
��=St	@��ich��X�P���+��������]2����-�1�x��U��е�A��K�_-Ó{�t\�LI�G���`��sb$�]�V�o��h��R7��U��P�VYW�Mv�B���<տ%*�z/[F��I�T�zwy�oS*T�M:F�������e,�4�O4S�
�^>�?\�p�'c���6фB
h(GM�[���z̪��,�w���f�e��������{,�B���A�H�$Ĩ�jZ���n%���uD���5=�Ez�M�&�xݤ�a�vE�X�FG��m(��g�C��e\��Y��ҳ�#n2h���]�%[<A��t��dZZxv}M��g��\J�vd��6e��%�\�9�fkU�o��f�Vf���]Ç�שx���Qr%�Gu��Z���/�@���;�p�Z��edh0A�$۔��F���9wX�<T��c%�d�m�7؉��㥳��_�xB�x
jRWB^"�z��=��9�\��r�"�0rP*���n����-Ux6R���x�pd�LR S��J#��"���!�i}$������x�
�0�oK#�)V6���9�G�ӝ�T�f��uHi����+��q��{,��퇬W2��-Q\���S�?�SK��F�3�aLv�Bv�z�,�uN���t���l"�����x�K^�)�0_�8>ܰv��5�5�bj�YF����|{���j�����u�U�~�Lu���O?X�W'�gP�Ϋ�]�_�����U ����)�)4-M��Q�����1�OC6��Gj�R�$��IDk�H��-�_$ 
��ًB��h���Ȃ�=K
�����3*J9H��n\u�W� � m,��kY�0��V�Д*���m��dQl�Y��l�%ڥmvؾ��˴]���t��5�wf9���z�^T��!�Pګ�芚ӆ�pXGxm�jHx�t]�ϋ��Ќ/����RWO)�l��>�w�7�ϲXkI[�A��l|���D�Q�CX�D0�� ��Y�HI-6��XW����ˢ����`$���.��mo������uqPd���ZZ���"�X2@��7  � Aj���c�/�Nؤ�#���Rm���A�v��΀gi��.����q���oY꭬���<u����#C����=(��Y|�-6L�F7�`�����v��x��z�����M��#H���x)�-z��4�ʯ�+ƝO5Ulo���R�~�Qf�8�h����Ԩ�2	|�	�����n"�w��b���s\ܛ+��3#�� �^g<<�5��
P�լ�TVgL�j�F8�ĳ�`��։n�<�7\e��G��U����3N��EE6c���j�����ݏ(�P��O������~�*�4���j3Q� ����W�/v$��|�N���_`�g�=��WZYh?+���t��\O�a�:S���;,�$Q�	��:l���#;;u��l&n����$�m�"��������g��\|&щ��<1C�%�2]n��3|��.��O���p`�/��~f�`��o>M�B�a`���n����B���8o�q_S��)�r2�i|^�Kd�\E�̱;u�,������:�y�kȓ|�ʕ�m����5�X��{GX8�x-6PX'�n3�@sed�� �mW�����o&6�"�����_��|>�vVj�\��y;d1�u�J�.18~<x��F	Q�����:Ъ���~�(XŖ7`�mM�U\#*�7n���cD@,����0�_�@���>�_���R3�,��>J�&�����`�xSOS�	����I�;5)g�^�Y5˙�J7<�	�.��2�x�"�Wt�Q��Ao�cђ��&ZON��Ӕ��hhҟo5(��ǟ�������+v^�瓥�b�H�����]eJSA�"�L�֨1��\���J�վ��l�����|���A2�Ԏ2ح0��7�-, Mvj"9:����m���6�AΊ4��t0ݼ����+�����Ҽ�ܧYL�B]:8"V��/�]�{��ܭ���'K�q����Il������?O�~����T��W�a��j��դ�����ε#bW���Y����E1U��XG�00�(/��QV.~��f��'��yq�}�#�yn��e�NQ�+��R�#)Q�.�C���iz<m�A�nQP���8����]/���"+�)�2k�
�D�l����^� a6�:s�.�p�A��_g��&!��R�O�����x��ݬ�.,Q7�y�0iI���A��Л��T���'`��! �=+�ccG�Z��7�����ks-��8.,JFWxC��	+5�m���R�$C�oܪ$�5���{,*�eiޑ�(��~u���l�&
h���jZF�G�� y	�4��:��j�:�1tPЌ�ߣn���"&^��ϥk�}��/Y�IAY��}܁I�3�&�����A=NV#5�\t��G��!�s#RV	U�zM� ⺛N�Uc2������[ft��Zp��`���!�C��}<�|j�� 2�UΑ�$z���$��N��x?��9o�%��1���Y�17;�O �v�����	w��`�D����3��L�wJ_ؠyCik��'
&�֢=d���h^$�1o�
�&�M��Hwj	�'�K_),5�u���ɢ+6� Ya����D���Xw8���=�x$����uF�P��=9m-�9�N��E�ȥ���+��!m�����f8��>���W�r�Q��QZ��)�B�����Z+U6�6����>�w��I���:�n�^Z��n��-�d�N�^Nz�w�׽�&,B��