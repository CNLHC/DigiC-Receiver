��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk���c���k;���5:,k3b�K� j���U��r�(��3΃��%,.ʫGHh��`¦f�U4�Z��Ǝ,�"�B�G!�&!)/����[܌�ń�=�ά�,1�}H/��PiY�RvJ0���T���^�E%�0|���D�i^i	�Z ´g3�ա#� �X���h���B~�3��&�C�I��s���h����rԜ��?0x�l���'��L_�:�g7�w�\n�U����rO�Z�j7�i��ٚMھ���
h��Ro���Z��;JF�� Æ�׮��LN��A3���T���i*#ȏK�@.%ܠf%E�����Y��/#:�{��m+Ԧ�7ܫ��8:f@����}��dB�p/��Q
�ڱ��.H+�%ede(�Fw��sUHxa�����陻�ƫ��y�
�Q�1��k��^ʴ�̕���l2x� �GQ�!���ך<$X��X�����V�����kkA�@(]�ƭ��S�+4G�IB����i���O���+�Y��-��qdV��}ޅ������j��LԜ�-���N�4�3sf�j�'�st�]�h��G1������#�s�y[e�F��ܼ-�䓣�Z%� M��������,I�;g�����_� z��x��s}nAVw����j����?A�jE�k�)��mm �s�r���\?���y�л��(E�M*��| �$+���+Ye�	q*��p��!��}on=��6�:w�t��r:b*R^h�MH~�;:����D1�S�Ah�#���e\AnH��18���Mֶ���[��z�,���dC-�X�$2��F�k
g_��|�mવ>,%;��/	r�=G��r0�f��w����kRr�h���v�~&n"�>�:{�m���ٹWRKQB���e���v�k��g=F�bO���m˶��Q�H��;���z��2e!��Am�P��1�*��=A�!s�U�N����A.�{u��+Z�������q~'�	��[��Lu��}�p	���^.�0�B�����^�\R��< �.Z}�P�	s,5��&�t˓���Rʇ.��4����h���}����e�,�@��
+��2��*.��5D?b� [0J@a�����d8�S��z� }��Q\��8wN\��^�1����pүx0
���y������j�X��Q��amqӝ�f�kR�ۢ�����}��M���IúM9GNd�WߜH�oM�))�0��@j̜/�{t�����op2k�L���U@�
r�;s{��S ��-�
h�
�r�.i�?�X��_7����tiH����A"CD��P��	j�)K͸�5��Nr�p�"�^*b��T���ҊJꌅ^��̝5b5�h`����ӹ���p��{li+@�uX{ㆋ�M/ং��0��:�㟣�%
�#���M��)��(��oӚ�ow��~v���],�=�{�����7j�7�ʼ���|�����rt\,�c��3�+8�|zcMZ�H(��s�Z7T�� hK7ϡ�v�g�1��B%��'iE�r��t��V8��ߗ�T��NOB%�M_�(��X���g_��ր �JE�=��C�԰oby95/Ӊ+W�p����}x1��H��Ĝ~@B�D;�3��2�O�UX~KPڬ�����U<��aD��9�����$�y�Y-�S�ꄞL����6ZL��c�PGj#9�/M�"�씌�mRG0@	l?����D:��$u^��"��%�!7�t���Ϧ�8w6���b����O�����|_�ہ��R�~�2mgYr���ʒQ�lܜ��! \Y�,QV�j��G
�?��=�n�d�/�}R�%X3ߎѵ��[}&{��ŃB0���%�,�Q�.���|4%�=;���l#g��|����'�/�h�-<��;X�K`
X��'���I�Z�Z�I��h,�İ����&n�j��7?9
�a6���gg�l!a"�n��������d/�u�&Cq�o��u��́�7��PԀ�>����&0eGK��U��b��B�^��=������_o+�uWۮ)�*�]��7!5̦gW���1ooE�p�SB��s7G�)Ukj	ϔ��Y�0 ���E�;�t[�q��i1�}��ת�&<���0��!��g4����RzH�:�b|1��9jƱ���Lka��ko:��9��n9:W�sԐ��ڐ���
�"�v�~X7�t{l&����[h3'���?>P��&+�H����N#�����|��`4��f)��YT^F�a��(���QD*����΄��{����q�8�b�i���|}G�[��_,	�S�1*�IM%���sEΥ�,!����L5e�)2�B���=I���+z�P�5���$`֘�M��&$S�)��)�1�޹��uF�ZT��B���y�G�Т�M�#�þ�� 8�8��m���d�c�����=j2c������� �J�.ۀ�WԽ+��xR�����L`���ݭ,p?x�S�E��Yc�%�T�z�䔾fc���Wn�y�zg�.{MW�s�v�[�?�6�y��w�{�p��Ќ�����~�M���ko,mT� h��S9��s��6�T���`��d��V{�~�Cz��܂9����l������J݇���\9��V26���s����2J���*�9d����0s�?^\�ίK��9#����R�@?��Q��HbFw�S��X�ۇz:v��`.�<D�� ��~�У�����g�Yxڧ�O���ax�U�J��zLV~��E`�%|V$�ԭ�.a��9L�ZI�,�����ved`����oe& ]�S��
�*���uҷc�����[��U�K���;͔��3Q#)�q(�ЊK���;8ZY�f����|@����~3 ,#�Y���� �#7BA@-�d����)F�`OT�D�n3/�>��.m2�K���S����w�KT�$D
��~9�\/8����%hRxU��^�;���������,���̀�=�������!T��k�ʀH��G����e��u7j$��8ii�!����K5>�M/��Ʌ��i;�ȍ�j�%��8,��4�͈�/�,
-��F�q�Xv�����&���%���)�/�`/r6����V�x�#��))ެ3<��c#������Z�&o�.3�`}�	�nPp��M��B~�����Fb˗��>.)r�7��qB�*=>!@����w9@�8Dze�Bw/�[ �~[w'@X�tZu12Fw�u��Z[��5�ը(zq��$�`}��`�a��O76t-�
��Sp)��m�eG�����r�F����x��]G-�u��n+v��Y�sP\'��POM!_�vo���$�[�R�N�/2����w�v�=����v����X�����j���F3��O>?�Fc�l����g������VOt8h?P���l�{QR��vccT8L����k&�w���)׺��ޒD���YD0m+6�[�T]n��6uFXH�>®ݏ�r���Aژ�
#�Y���K!q?��o�9�8��N����"��x����d�>��$�TP�����y��̾�K��E�� ��dvwn��~�'P�T�t"���8_^2��&��8�"lp�!�aH��*"�h�7�F.aq��w��'���H���˱ٚEYӯ�!L�VK!�Э�WU �t�[i��#J�����S���.�E,{�[4X2�tO#�9��p�r�q�`�Qm�}M1���,����_O��8|/wU,0K���	W����u@�����gF���;w��K�v�1v�t�#Ϫm��¾NX��fg�W�_j�Te� �4`�u	�D��@�}W�_�9�v�d����o��I���E�� )j���_�tF�� C/�1��V���aM����m�n��6S�Am]uGc��G�lP�>w	�������='�N�ݙ���Y�XT}TKaJ��m��Q2P�Eb~�x����6�ڷZ��2JZ�E��V��XJ>��W�m����ߡ'm]�Pt ɃAgFg��@	\hH8S������6A���r\�N�XI�V�������0C�tM��Y��@�i�)���Mz.v���N�5%�?�W�˫|+:����Jm>�M�(��
0�ʅc��zyq
��	�0�����|��9��٩/Ƀ�p��w�a��=zi�ޫօ���*j�X/�n)�|I#��8}�0ݟ�/(d2-�uS�2�U�X�_�.j"��p�1Ō�nҬ�vҽ=�T��cumRB�䍫�R����.�,��}c���͔5��4�g�*햮;�<��k��#8W3������D���j��4<H����	7=���>�9�>�J��L�1J ��έ�y͊M5��"vmr�jO'A�}>����M���i��Pe�6��1��&)�5��猶dns��Y  Q�HJ�����s�"@���������H�ߺ��a�رP��_�v	�j���1@@Db�6Ls�:�_�l��5���$�E1��H6�v��H�&�V�w�I�l҇N���be��+�V��w�.@I�A'Z���	���Ŋ��`��N��:�����k>�z�DW���/�XO\�&ً{���8H�K96�H��e��aرx���6}*�R�C�h��~�R��:�^gbw���N1��˩Ԁ#�0��-n�-�'�>��qA=ǿ\aYGGU�i霋�.�h��:
:�~vъ�3��B2B#R��w��=�L�eH|���@��ƈ�!��;/tU�V#�Ë3��H5��h��P��Ĭ��Ͻn��9��l6�U�"� �i����b�ņ�	��փ�^2��G�[��g�{>gb�ع�x /���	+tm��|%�h[�� �����x�E�Dk-�d�C�+I{l��A��C6���ɒ]��(�hl�"Y�Y~썋�6F8#����b��(V`�����g��س޽�4RD����7rh0�񛁍�Hm�F�����pp,f����(��%�L6��i9)���T9�����*V~�	,�}� T�+�ۏB��I�|P�2i��bHb��C�!�ĵ-iR ~���\�,�'Ӟ�wZ���޲A� �Cx�G�i�FVH\%�!�h\)�nWq�+�@5��jQ����̳��3��[5-:{)�%����l�
���FX�h���Pv~�G���7G�bU"�bō�| �{�98%�h�-L~�b��	�Cu���ot%�>�k����+MS�f}�'��+�#<{Oz�@����t?wo��/�t�rcD�4Aک��vŏî�\�X��L�w%�*P7�B�o���_�Q�&i�t�G'ˬ�n]����\����5�+��:�`]e��_>��]k��yc{��
������4WI��,�#8����8�T���y�jY�[ ���U��]��w&�)'�����#��(�a��Z�E��<y�)�{A�2H�����<a���nOjp�
dh���4a�5[�Kh����X���ލbm�)j�&xϋ峉�/�F���f<gl�g~+(������/��y����=,���#�3�v�䜪8�Y�G�b:��H-:��_o����3�$9�9�,�A&E�	YgX_�\�r��q���T=�����tk���P�ɛ�"����JR����|�45�XD�ͮ#!c��"P�������Ò@��� �K@=�,Z\?�����z��	�%?�kD�m�EYg�^��Q<)8�JB�r՟����j�������q�d�V����Y;��(A�q�R�msREѓ���,""��"�T�":��#0��=b�R-E��΂s
N(r�lJ��K��R7����i�o����'o���Ъ���㼙(�])_3��9���)�܆qgj�Z#�c/:�3�� \���-�h�1�A"���)��Rt"�<�G�Pdvy��,Fe���T��L��N��'��c&�ܯ��M��]���>�Ƽ���n$�-���D�_�<�Ҷ�y����hćzF�[��7����2i�k�^�����Ǖ|E����:lv���Z�d�A��t:�J�r5>�{я�Fsa�2�z ۚ)>$=_�����/�;'p����]~����qՉ^Q�aE=o�������B��C.-�
��s��T�Т����/~��o�r�Bǫm��*`�nNJ�
�^U�	� ���%��c�N�yJ	��6�+v�A���6�F��!-p*5�3t������k��تy�.�n�Ģ���Eel-�����lU�|����4li�/s։-	�[`�]��>�(�e��&�Y|:���{ш6=g@�}n�����#�t�	p�`��[�֕�_���({F�:xA���@�P��5Ȼ[[a	���M�+M�	|����i�k�U|.2X�1�S�	��d���!��O�qohy����h_���ߠ��b(��e<�R�
+e
s�|�����#
�O�	��q����n�Ǘ\�j�<L<��N^���� &�h��N�D��4H��$�n��Z���2�5(��fj6��dW�j�'~���K��O��;���w.���C�(àPǓV���籋=�>蓀#�Z�c+�A�쮈�@w	=�c`�d�5�_f4�	�2�p�د��W�Y����&�L�*�1fҙ����P2�D�3gVw���M�H��<��쟇+����1EAP%]�F�kb9T�9��[y7�fP��!��ͨ✤,���5n�ք��T~�Sz��,C�"�)4i�w���Kf�llI�����E�������x�P3~Gӫ���w��?�?Ɓ�0*I�y�_wi��K6��7mb
j��tL��b�ثJ�����G��c\SL��|g���s��s�+!I�4��T��+<o��}[�������dv� �N�H2 ���O��iIg�J��U��)���� 7JrS��R�^��x�=-��=\Ƀ������v4A�$�$8P{R�4�j]�Rk��z�":�%Pu�ȓϰ^=L�L��r�J�Z��<lL�a��z�uR�,&���D��꧝�h�Ż~ s�7[�k�\I�T�㘢��?/B"�:~������5V�bO���@Z��ui82��1��7,��teCZ�;�U� ��Ã�J�L�lإ��K���6�T吠�\#mW�l Q*5�����ëq��9�C&������_�U��
�Z'�u^,�ܢ��yN�����h�A֍+G9ӕ����Q�	Y
�}Q?��
��47>�ը���i����~�x����	T�[�F\�S����3sTԁ�jv��E�9-n�W��
I�5���l��L��z�F���\����y���O���g0n?7�[l�%jٌa��4�h��\K�NH1���2��Nq��z
As�}�F�,�aB�x�
7;�����l�@��P�ڿwhi�xZ��mUz�L�p(�6��"�C�x��(��2W�1c�ʄ��>*��'�w�� ]>�0{��G�a�w�D��������V���Q�)!���I׊����Z�b2/�tެ�e½��EK����*�ƅ-�&0ِ�)(�"����Hn.1Đ�d�z#?_���p�[�\z�7�5䖍���i{^�io;#䲚%U>%���R�ѥ�h����8�i1E��,ǃ�Rol�n6 �ZS��Y����܃�w9�:�6�
6�K��I_�҂w��hr��.|���%t]YQ�X�*�:0X48����RT���#�3̉w�<�opU�8�������{N�:s2V%N�d
�W�W�b;�%P��M�O�7�*_ڻ��+�v�ŉ�_4,��Vu���`������B��Ur�"ЖF��@{ô�lX��=�p�\�O�6oNO�nc|�+��iPvɹ�T�UCx�஭�B#�
 &��q�6Ë
�Lfl[.v�f�*��eQC'^'3Ku��V��Z�j��=��k@BU�����׈�Dt��Ni�Q�/�]+1�PV�i)q�s��Ѯ��#"���𺃀��P�q��΁ xEۓ�/�BR��ʲ`~}D�:���tӘT��I����n�ÓS�@��\v��69Uö<Y�,��'w�U?��t�@�����*���)L��ۻ���+�!�a��D4\��-&vTj?�T�]T;b~#�����#��<��X�^�
n��S��ϸס��@gOBìc���r�Φs:��'�5
���?b���'��_���-��k򬫴7_��hQd�l� a2Q)��^e<�	u�ZB�լ$��bJ?�A���a8B��*��x�IxV[��e(9Z]����&�i�+a<g����b��"�f���@f������3���%��s���N����K�*��.^�c��Ih�%Ͷ_eG��Q�|�O�0�Z�I�0�#�#{21�m&f\��e�H��(i�v-|�5�i^ f�CZ���od�r�qu�����$K��y��� 5�����^�VÞ��� p�mB����	Z��ns&;<~�^��o�� ���	:�ƩW�^S����4SJE=[�R�����`<�_��t!�� %{y��4��
��_nw�tI.�&��� zn���X�q��C�K�y����P��'ƴ�|]3��{����޵�7UW�U����#_�)�:�ڟ�� u9����=�f�`H7�rt�m3S��Mc\��X�q(J_K��L�q>��%�Yl{,�����4�|�~3��Jgi
x�D��sB��?� �c��V�6�Y�����N}x�G�M;#��4�R�9����"�&I�N�Z��漇q�MS<i1��9~6Q¶�%�>m��̫ `�q:�+�ZK�b��f\��>�`������� K-89��k�Y`Nֆ��t��D>�~����cgH/��x�i���Xy���,W��%��WN��a~{͓C�b���b	A�Ї�E(���]3���ޕ��x.� �%S�����7����~A�Q=����{�Dx"�r b촬��`Bb'���C�8�J��(��9Yvk8˯�~]�|N�XlT���`��h��\�~b����̻�)�??����|�'��`>�+���y|��$��!ycU����F_��Z�z|�`8��I��oq��z�y>Ͼ�Ѭ�'`�U�e����UaYL���0'�kī}Vǳ��)[��$�ȑF�)uf���О?���~:��V8��kr�7�o[��mh�~#�GhZ�a���aoU[�?N37Cn���?Fa �$�!$EP�0���Q��(����|E�a������Y��oz<�k���!�7 qF �{�ê#��I��I0�9�cv���H,��5	$:F[��˫Jd'%=�ZJ\�2����4������}���A�$>1����*��bn�	#>���A8L�o]^�{?�� �"}�zL.ҽ&g��C���Ưy��*ڝQ��_uo��AJ�P\���V���/N|�ע`ٱ��U����/RNt�{��?��F��L<]}���@�2��.'�X���J����z�f9��	DIL�����vJ�;�+>�)��j����j��{�=�kΡ����;�NhN|� ��J	>]��ҡ�T4�*z���b�2���PG�|�=�iͧŏc8k������D�?��v1�3i������6�w�¥��/
a�8�D#���0��	_���}�D�ukq��O�R���{��������L�r�9~��y{"��yd8�J���,�0{�y+�a�0�)���`�%vZK:pУ������F��g�v�����8�ό��r�4h�S���7�
7e�bp ����.xn�)�gPG�N�Fk"nO������n�r�p����� J)h��^�^�R�ψj={�?b��=5I,ի�]��f)%�
A��]mP:�;�òs�'��!Q���p������*�6���4|��+�f�pA�1#���o,�V��b�A�B��Q��V.�9@5����_�?�.I$���mGK�e|3��ૼ���f���u��!�~u��-nB�RLl:�%īH���M{�j�)vpwʑ��-��b�o$�
�����+C�S���F  O��k�<�NVm�������Ύ��Ӳ�^Ŭ���%������6���o�c��s��Ԩ-���x�]+��~�Tf\-�&��0)u4�ir��;���0�xr��=Ho��U� D�����@��ѧ����Wf���]U?�)b��'���"`��;�U$.}��0W9S�#L����@gĿ�7���qZ�~��P3�Do���j��^������v�f�p��a'�4�^�a���)[x�"-��Ql�����ѷ�o�x����p��|���jw�E�f��q��`.Ql�H��r�2M�a�͑�������	օC��&�C���]�bm��M���,h{_X��ৰg�y��#|P<�+V�}>Z_g�B�+v8x���15��p�lq�Y����(�J�9:�v���?�z�н�2�[Xcn�!���u�����=�p7y]�q�_\Z��,Ұ�,2�.U=a4��T��3���� ��j�bQD���p�.[彺  ��Ƭ&��NO���o�����Crj�f>"_}���@Wt(E�x��ft'�!�[(�Ǆ��.�>P��nx��-����J�Uߕ�4D�T�b�Ų�_�vI�+�]J�ݣ��G1�/z�n�T_PR�+���A����ks�6 �����Z.,��j���e�
�D�j#!���Ȋw{<&	��C-�C�pT���։Ԙ� �$�p�����e�x�d��ۑ�M���L|v�M�n ��ǻnp��.W�_���t�+V=�,5��XO�`��jUSL�t�[Bդ� qa�����/5����b�*8We�,���.�oy�`�,�Y���_��7˿��g@�*I���fd}�d��z�-����S��	[t4g�~0��/�)[�n�,v�* �_;�#��"�b��&��sd.�@jS��kn�!�l�5ϥ&TS#��B�����C��#Cmg*O>��b�#�Kz~�����>��ø��L  ��o�O���Fy�|�	��
5���.�t��C�%���� ��/9귱�����T�}t�՛:�2Ut~R��'��S��c���q����VЏ?C����Ԍ�G�)X��UFe�"�E��$��֦S�M��B� ��z9��b�����9܊H����m��iS��$��P�<�  )���/q3N��X��ߙ��7��Y�:���8N�9��<�Pl���Y��p�hPp����V5��:��C_7�h����R�&��ԥ�|u-����F�׃\Ө���KJH�w@�����vի
$��!�#Y��%r:|zV��/?�C�K?_��˦]�G�R�;��Ss��u���1��S�w.�C�_r+Z4{|9� �Y!&e���,�����ɶ)Κ��"_�z�f��X��4���ϢqH��_.-����z(�֌7�g�&�s�6@�}�^��w��(��u"?�B��κ��dq#�H��D��h]�׻�V��0���
 �۶B�˖/`���:Z� ���
�e�zR�9>b��qX�Z��j��fH��1�eew6;�G��Ik�{ႌo���Xĥ�_�&��C;c([dR���Q�8�ݵ}���ܸ� �!ċ衖{Qu%y���a�I�b���(ѩ|�_���[b�s�SFW`�$�e�jW�X�!���h����^2�����݆6��-��Q�z�1xhnN8�N��k�.��.���Nў^�:�q�k �޴�]�4��x�s�2�x�g��̂&�d-���Q����ah��F�dq��m+�2�}�B��ޭ�x�0X4"T��k�<	�����������W��@�A᳷�V�|�cB���MnҞ1Aҹ�L���gE�.�)���ż��WG���iz�,$��xH֥?0�����ڮ(�[d�R�ԡZ��:\�N�ۙ�m�Ֆv���.� �W�,Pz���|�x�Q�C"&->!Y�R[�J�ӽ��\e�Wq�5�ꀀ^�{^���[L��!�7�uv�Ĺ6��o0J�!���u:N�T`N+䄾ڒ�u>G~�,/�ϹM�<&h�����̕�cp���͋��[�',يɂxF%UEO�ǁ�a��E�H������S�b�6�C��ī+`	��{��R+�%m�M����e����RT�
����E�+����ZC�w4�AE���� �1��������2cb�0ag���6v{+㵩�2�!H��.�	�Kf�ֈ�K+2�u8oD]ܯ0~���#"L�M\C�G���G���X�h�� �?��"g�$S���3���qs������\�$()������lx�@��q���>�
���k��L�$��%��9�������V�uf�S3���4�"���Y���ONK� !�����+�[�+X�,��/#�É���lz���_�m"ݔ���G�=��ͻv��9�0�7��F о3�= ����f˟/�C��`���=�'�:蔒��1�U�����)��\��Cx���'Xy��i���<}�Cm�J�V���YzyѦnc��n�Jtt�'�G�oW�۽�'2VC]���I����Џmr�A��<�mv�k���� ����S���3����VYN��ŋfIKSgx��;e<���h=�d�[�g�m�"�����+& �Xl(���Y���^��D�^ԃ���x& ���G�M��J9�}2b��=�v�v"Ef�@V�W�f*���)~�|���C�b:���j���t�ax�\h4Bs�%%����0����2��/�c]3�چ��j(%Vy��6��Q U[W��~�s�:Bq`9�����*��U0�<�/��/:�
�w3丢�{W4q�H*���3C}҉��cҽe�D��>��^��u��/i�����dd�@��vC��(�L��ht�ۜj4��;�_�=]���u��"�ᆚ�iY�Z�S+�M:h�{;�!0c#�IX:\��۞ %�]��B��7�@���.�<i�(&ŭ��yJ����E* ������%��Jj��ş���h�2��O��	<Z:�!œ��G�����m:�� 	�s=�J01 ל8��G��kT6�&��S�Ȝ��>5R�5"H��JFt�v{���p�G�S\�'(�.�̃p��MV������Sc��wQ�a�{GC��`�5�el��
��Q�
�L�N��x�T���k���.8y4%�����Xy�� M=3/�Z���h��<����-��V q����G��Mm@5�%��R4�O��imNB5��}rX�Y����ͽ���ԃM�œQ,�9�K�,�ȱÍ��L��UW7e$��&��#K���tD(��lo�a���k��� ���;�ID0���͝fh�Q�2�!����6�����{���������Z,6E�Y��~�f[ �t���s����� *��F�YI��]�@ڗt��y鍁^�=^C��**���`-3��5��5�6�%o��mP0]�`�A���%�7�Ϋ���	ȡ�v��_�z^j	`~�j�q���F��#�+�ņ�`9�̒��Y�|�]8��-DA�(V[X%�s��h�)�l�^�����{�qo����YqJ����'�u�B�� �U�.�h�����蛂��ۡ��:��?v�nmA\vۭ�K~X��j~���*�d��?8�� S�Q��
�v�'��N|A������w� L�@����g����
�a�GfSp��}#��Je��$.b�T�	5����������\B�Ly%T;�v���e.r�"� fi70z�?Ÿ� 	9u\�Ms-��=��lF��j���m�p��e6Fƅ�z�vТ`K��_h�����8��$K�Ͻ��J�a��j��O�������F64��e?��|� ��w^4i&�r6�{�%��n��dHc�q�}�沶���q��H`�1|��-=���`#GK�"Z����� r�� yi�<0���eya8*;^�>����p���9�k�]��d�l��'^�R6�hsg��c�,�$ʒN����kn�S:��O��=����'	�7���Sd_��� 9�!��4RK- ����H��+����5�=rj�I?�u!a
�Pi42<RӶi�O�ꬑ�,�� ��[m�]N^���ţ3�)�^��B���"п^(r�Y�*�w�]���Ѐ%,��ȫ��ꠌo�uc��=5�Kנp~�Ư���yR���ao�T���1+J����<{��tJ�C;,�_�Rv��5i�l��8��PGi;��RьM�@�5�7a >�&{��+0��& i�׈��œ7����ÚHz{����>�a�wC���(�ޕ�E=%c��G�D��{+�����ӡ����^�>t��o�ǩ����U�J8����7�h/e�vLo��J��j��H��U	&��EL~�M�U9�͊�i�����[)A�\:Xkq��2�5W���,+��<�km�SY|�Z��8bҷ���5�h����'O�d�Ơ�a���X�-���>�W����dv�i*B��tTkA�K��,\�1�O���! ����'���D�CC��`�	Z�hF���ի������ T�Rk���^�\뼐������>Z<<q�f�G}�X�M���_�AG��(:�̸	- AV�Ui鲘Y�L��ͦ���Z*x!��H�$(�"\���hez�����]~���g��R�6 T��D��Jě_���W�/�VB˓�~@o��K�a�L	�1���p�&�*��B$��K��-l��l�%�	��3�8�bJf��s�����1RCjE�g�.y�o�XUx�A�>�9�T"J@Y@Z"a�Z����s&�/�Y�B��[�L^ݸ0z	~���6���Ɓ�@���!��i�<~�Y�
���!Gl��󶟲2R�+ t������������^,��/�G�Ҭ�&����Vb;�Ы�I~�Ơ�#p4E�mmF�F�r���Et"{�ݲ&@Dd�)L�V���$��T���Z�4d2�a4�y�
��@!q[��jЃd$m��9�QjBW���)��8����R�\�H�W	h9ъFl<���z��ѧ����岗�.��;��g�N�F�ىJז�j���z���2��_*�]�G�o6Y�:�����Q7�x�$q�� {k ٗ�{���oj�����ջ��P�iðA�^�J�3V(�z1�,�+{A __�m^��a/b
ҁncޓ�H���p�G��0�s6<ɫ��D���=�xn6�"a{��w���rna���\�
�!}=s�G�%�)��#U���u�Y�S�c(���q��)!��O�|_�xaϣ4���*e��H��hR����q8��;���jq�k.�~l6��΀�Ғ�����]�����x��T���<��"��X��R��c�^�f�Շ{�ԑ��%�ه���?��|2�Ԁ��<���^�#>��`�;��;ݯL�ɑT(�S��0���B�mX�у'|
3W�h(bwb�f&�RH ���`�����~!����Yc�����*SYP��5��5�aͭ:Iՠ%˩W��@F�\�����Y[�7u�����ۚ��=���êu��-P���u��\�
�]�f&t���O^+_��qX4>�Z��z:u�= �ܭ��T��ؽe�?(�ȲK�.�J�"�E��WSes�+y�&�Iϛ���hKW�O�u1]�F!;��ʪV�4 �8��_�^���0�c`s����ӻ����`Y���&���a! �7�â��W��6�-A�\s����f��S
B��8^wd�߸0.D*�xӇ����u��Q�]�o�����%�ы�+��ъ���>�#�v��������0�Y�Y[�q��	g;��#h�z���;��D��nʈ<10� ���4��h������tB6���{*H ��Ҙ�c����ė�������� �[ތ�`7v6*�&��*udU�
��x��qi|�c�Ôe�@���>�F'3���'�ǹ?e��so��A�E>����2!s�������ٶ�@��vn���Q�9�j�O=)�7������(�����Ub7�w�/��h�B;��Nd��s�o��a�}G��l���������"i�Bx�.nm�4��`ّ��ZǙ�{[@̋��@ͮH���
�P�j@��0��Ԩ�F5�D����xX-�$�}'�NrI^v0�W����)���X�A��s|�-�J�G�% FJ��4�ճ���q�67&]�<��AmmF�!!r�;�54���R�,��{�qu���+���B�,5�(�te���pE�����7�xo|S�K�% �Pw���<X�ȏ�A�w#`]K��b m75��-���:Υ�݆�FN�A(KE�a���I��K%!��_�&l�몱���b��o�s�6a���5K��P��Y�CB�"e�j�U�x����d$<9����0���P1�q%a�1(�)�r�jD�1J���<�p��,�@
��+^y>`�
�� D�ߔ;F���g�H�j�2�M)�J%�Q�	c.�1Tٕ磞o㚲1SGJ�LՅ���ch r�rݞ�!��W�%����{��-R���>Ŷ����.(p>Z��������$��95�SKŚun~-����7%�6��{=xo�i��o�����h�Jx�L,�:��+�ˑ+洢����О�ߝjL1Ũ�Ev2I����[��٤��G������'1��m��P���d�����"���VTe�<ʤ]��r�g��2����=�mJ �EE
����je糏\|��L�h�,/|g�5xOS�V,z6:Ԭ� Wj_.��x ��+��j��\��MiV��D�Z����^�����K��x��Ug1��0��ӯ+"��E��訌���1��u�I;�}.q�i�oٶ�U^�Ųչ7Ϲ��Z��\�bF���3Q�����XJ���n�M�ϏI�����Yٰ�fiH�Z�[���^��f�����u��䶑�]wi3����QЮ]�"�M���8�G]�s��Փx/9�1�y't���x䷘D����o���B,�q�D���\:�2����G�[�H�6Y��\�q}'b�;���q���-�k� �a,ʝ"����d��_t���J]��t�W
l�>�[೉"q�˙O]j����x�Il_"=��h;������e�O�Vk,�N?|U>�[�@�ћ��{�����j.�vw^�$�V܋=+�MoU|i�Gxٍ?��V�B��]#�M� E@��9P��@��4�s��K$�N&���B^�+���?����y�4�ĥ�i�ٖ����Al�:k�mI��ϝ�v3x�+]����I���㩕�χH������+����`�hU�-&0��U�#P2��PI��<(�"�<�,���7 �S�`�6R�6�t��dR �������?Ћw7�7�_���ేU{(�]�@��p���'>������*�����%�pO�{�^x�wj ӹ���DV�gꀯ,��jEG�B��޲Y���b��e�՛W\��Yz�f�_h@���_���gk[������z���[�pc�~s�����>�3�z}	�:?���L'��_=�
�k���]���z��֘BN��s�g��u�>���EݛQ�K);p���3�?d�����0���G��j�������\�z�e����t�����*��)�������f4:�~>L�-��F.�w�~3ʐDN�Xh�:�IE�
 ��B�̶x2R.$߳�83����ԃU#�ۂ4���;��k���/+}8{�q��|J���on�a��'g���>hA�AN2�^�r����TvL'�����kː˲�j�f�=����TK��b���Opg�b�W�`��k)�P��b�J�$4e�(��+����8f���w��V:���!�;��mV���l(6�u o�c��b���*(�i+��'�YyZ7��~PA�Ǌ>'8Rdy�ި�-܌�>S�a�8��h)�����umu���#Qa�� M��R��l&aˌ�)�~��E!3�V�9�316���j7��uV�b��Z�z�z�W�XG7��x��3W�+�9ρc�{'��=�����%�c-�g}גv/�M=�e��i.t��Q��Ws�f��ߖ��fi,�5M��O���k��鐰�E{��L�s��h��i�	�a&K$��{#ȋ������ytC�=7�7@��z�?:�E�`�/�mC���Dp*�݂p����ߊb���`>]�*W�UPǮ?b.2��!+�{��>�ܧ(g��}ƃ�kY��,$KX��� ����Ei[h���Y�(����8����3�0˘�%I+7�^������F[�B�#~�W&Y�*v�a�����b����/<c/B��`��|�ܔ�<2���-��O�PL��Y�I!,����e�$I�@aj�"��N�,e_ %��
���׸ت+���fI���|3_��K=y'������
�^v��c����A��$�g�Fn�{��������[�e��K����n�Լ�P��mQ?g{�]3�!�A�u_ܝ�$�<����{�Gx�� ��~={�����}x�<�b�|P$	�,ゼ��J�\�ETx^�xI=~z"f��"�D��Rq�$PL����!aV��ge">j�ML&��i��$y�Y��<�P�����y3�z�8��fi�Jj��
tk�QPR��F�Y�����Sc�3\�_?SZ5}�	�Qc��澍I /���h�e�E/�l�C(EާYH@�Sƙo���u�H0���	b�c��f���j�K�d07��{철���h�D�P|"�zq.�Cݾ6}��Q'��'�+b �U�3 <���������
��{��(Ϟ�����=�4��/�thtG����D��ְ�+H���2o�T������=	�DC�f���ZM���� ���'%�L<Tb�,�[h���R�a�_�a�ׯh�k[�"�<P7NG�W��=��BX�T=� *���ެ�4��*��Y���`��x��cf��E���ȶ)��y��e��nle�C�u�Y-��y_o��
�о<$�%���	��$T��ˈ����QH�x�X�h���'�����elN�lWJ�`��q�	d~}��攣7�y���׏��k�$�k����(�n����~����π[�#���w���?�Mp��2oZD!�6Y\N�v��r3��n3��f��r3E�!^����"��P�b�q�Tަb���f�B�^�
W#�Ջ�E��"�1ڃ�M�eke�VJk���k��ۥA���ӧ�M`�LM˼�,U�6�Nv����!/�A���=��)0�;J��d��;w�����^�š�\�V�� �2�V�?����Al��>4W�\m��y݉�ߕ��2�n�\� b����Ed�U���! x�y��:�t�h
��i]��Y�Պԑ�^�Q~)sl�n7�������q�
K�<*(&_> �˄<��㒉�)�0�F+Ҿ=y'h�S7J-LN�&�$�R��0�����鄹���0���������T�7��Ξ|2
.>u�|�#���<��h��tȲ
�~�Lb:)|�ޭ
��yVɃ�	��s�8�(�B���#���-Ìڮ���H�^�����w��6֙�`��~��:�v�c�$�����[�y�<Hr�a'	��#�ᎇ���R��oЛ��U�����Hhp*���B6PM/�Q�9�J��c�� ��5#��E�����Y�J�k�0&�.�2c|�!�9�,���]T��D�h��_WQv>'p&�Ui���`�-OP^��[H�_��{`�eZ�d���V*3v�-���4B��f ��S�.Q!�Sg: �,�\Ŕ��L��s�/$!��]��"��s;��G+�:5Hk�W���d�l9b&L�� !�[1�Z=���`4@>}Q��%7<����>�l����4Z�¨�n��wF/��7��:�lV�R��Tȃ���?�v�w1����T'x��J
-�E�D@��@��h�#�J]��fFG�5`��XL����o��a��/�V!良��X��G��jS���Ue s�#�����2.�5�aT��q$Z���{���ո�Q�C��a�^�#�!���"��<�`�En9+��&���p�KO6l�;vQ�I"��$�W'.h\�<��[��tG���%ۦ�i��	��2o @f�*�n	0"}T7+��]�#�-b�7z�Q�牼rIm���;
{��}���B��B��N w�dpx$fy>},�h�y����7��$a���@�!6~+	�ՙ�v���|��jE8�OH׷l����h�+_v@궍�����
�p�5�L[fp�i7Uĳg�I�#�x/0X�@�������r&�;������@�*'�z�6���g�&N�[��f����b
���ܑX��!A?-(�y�NO��}����Io*qa(/&������P�;�k����a6&�_gԺD�T������DP�_�Kn��3Y� s��6���ĪaI�ސַ�o>(U�7^sqh%T�R���5�	�*�)��[�>=�z���)��|�)~47�S��nLf4WJ"m%�3�AG*^)�g�nwo{F��i�U�	�<Yf���-O)ﲁ�Zy^�HВ��U�-�	������s2��gi�і�������V!&�jH3[k2���
vѷ ��S1�>��~Ȉ�\^�cGu{�
��X��i�y��=�SHe�S�Z����J6ښƣ�x�uv�LȥuU� GV�/�onq�#��^�ʷE�t��9�ي��Hx�A�C#:#�C���,���g�@���.�A+�DB�m�0#�v����0u�K��s�����R��fhGe�T:u7���!kx3���g�����]�+Ŵδ��㎺�_SHg|!a7[Y�.|~��-=q���"Pm��K���2J}�'��Zs�>�F�@��`�-󗳸X�[�䮸��'��/�	�v!��#H���>'e��Z�:��NF̵�|dK�g6�����'��^�}�L@�+����#.����	>^w;�h`��a�zh��൱kk`v�1���_�|�f��k�A��7�D'A �/�ox`��)��������/<Fr�A�>��Q�v�<�7��
��� ^z�J��8i
�w�K���E�v��e�YHZ$F!j�\ۦ�
����J�5�V^X��a_��+�����v��쨨 ±֋�y�B������-_�i�Z���u�G܁`�zŽ��X��!yY��HXI�>W��;ߓ�ɚ�.�V܆P��ݱzpE�]��O��g�Ո� Q��g ��������۬M]̤�Q�R�����Q�	e��U��g�tQO�4h������xw8}J�A�߇�r�T2@-�©��;v��Љ����ͭrF�{=���Q�գ�����=���D`�'���ƺ%g����{O���h���롵�̓�StlL��JQ�>�u�N=8�V<~
�|HvkC��3�(�L�E����'�/��YP��45m����v3Yɦ��n�,Hdm�U1��t��}�S�~��Wf��Ι�EEg]����(G�9�J�\:j�B=+�=j�o}�����䳵�.B����~�VB]L�2RA^�>���%i��7��u0N�����m��!+6=}�UY[R�R3�M�� �y�
ŅI��KZ��lD2��W�K#"ߧ�Wc�P�'[|���~�M�*%D��pzc��L�:7떦r�r:l>�|�G��FHR_�8:~I�l�dN)>��b�NO����BTK(>V�Q�������H���*��/����K�0T��Ax/�H��bF��f)�ó�lh�ٝ�@Hn�qv�M�9���3:�rU[^��+�uF�^H��-��Bn)x#�1�E��+��S-�D%��z)O����C🗑�=���ϻ�*����P�ӕ��V,�c�hv���}#�7E�)�)Nˣo��r���W�	+�Z��/������ɽ��<�`�W �-���e�]��r�Sl� �#�ȇM[�ʜ�̡�+���Ek����`\�O	a;��ɷ �[�F��&ty�{[r,!|b��FY�Q�Y�ӵVӕ��X�]� ���ߨ�H��~��Z6�I��`5�Po�xNYf�(�c��=�A��'��j�Ȍ�#IϗÍ\�֌H�+��ܢ�~<��7Qos�b3h�̩�(��8DJTu���4A]����a�x�0'XE�^��.�����*��_p�w7��.􍂍E�^�;h��^<�.��ꏐ���	Qdf����=x��+h&wR0t���J{��v�_�3�5�qs�D��tL���f���b��A9'db��vc�"&Q %Z�5��Lv�����v�e_�	U��
!��M��/2g*r���v��?�X��n	�wɥ�������ث)�2>I��:�������Y-���O�����*ɬ���Y�3"�]R�)+���=]���rO]QF*���Kd�w�P�"�C�7+Ȉ�s�2i����}c1>�+�'nȚ��H<~X�{����Zv�j���.�d]`^�b�u<���Ys��0��]J��+a�ae�Fs*D��浾����.7E�pf�̶@k�2wv�d&���M^4��"w��33���vʝ�up��!(��t��I�7�k#ue�	��򾯄`��.3�� ��G��V�g^Q*1�N4p�#��|�RR|���gL�	*��3g�x�;w��,�3��<�v�UK4[���+�(�v��nc9����D5����L����&�$3�� �[����j����~G�2_?9�y�z�l��@Q����2��}����5p��䲦�]1�Ը���~
DF�Z�1���*��C�L~i,3�3l�}��ï͟�)s� Ǫ|��-ZEשMB;�>G�Z�!E~�!�o�.�S���R�B�P�I{����f:&�-�c)�y��Ե�,R�k|K�辵}U����2N����Ũ�
e�g�H[��� :F��3�*�j4 +eO��E/ɱ�B�3%� @8
����5�D��K�����jO&U���Eb�L����[Y�T������L�FE�7	���^Q�u�����AG:4i���ȓ;L'���f��t���fcbk=4��4͂-?��	�8m���]�9�E-��AyH�7���:�p�Gt��َ͊Ss �ӶE��)��˘B�V�7��5z��m;�j[n��T��7�4��#�QZ	���\ȓ��5dS�Z"@��y���2u@��G�D���Hv����B���&�S>ɂVӬ��1�I��<����-+�P=|N��L��bwX^���ޗA^;�� C�J�R���9�){)1�6�_{\�Z<���x�ʔ��1�&��
��ݾ�u�T��D2#�=p�%M��-�,[�Řr����^3 ���������c=�����1y-��&)�gt>��a�|һ��'���3�W�fC1��Y��ҍ�s��e:ٞ��J��Zb�����Z�n������C\5��PT� ָ��yy��G����A-ǩPCد��52�W�׶���\�0��g%����<��$�ځ�3�
q�p
*;�o�d��`9#N�����Q�d���� V��>���e�4���'����Cs������C�1��M�m���[�ܫ1���_��'�w�xh� ��\�Υ&Ġs�!�nj�	!��B�%�5��ߍ,�2��F��4�̋��=�����@�߸�Ѹ����d0�v�+Hf(]m�ȷn�߮\�A�/����2G��g�s�G3��Oͼ;ؒ��o�n�O��ͳԠ��*]j�hj�Fij�l�x�*~��[��.��m碚�s*@w�,��jKi���g�)k��G{�j���W��b��WD:� ~4�!��9`��|�N�h��j_ǖ����3 �eA�Z�X���3���na��m���(�J�D���"���A��'ǴՐٻ��E�n���G�D��r)��%�0ڭ���=�6~A��W{Po��v���)�ۋ�'$0K��/RZ�U�F	�B�b�jӪe�0�{5�_~����rh1kÄ\+��f%lisC+K+h�@�^���;]k�KϠQ~,Ǫ!"(0h&��oT��1�,�����i���>���@Hn~�=�d�"��b=�X4�&�.�m"���:��ŀ zb�tL�����:��h���W��=e�+_��U��m���|�#~��A&�3\�����ffh�<RI���k�I��8S�V��f�e3� 
��^���^���ۻ�t)��l)6:dz#)L������_T�0�&>����YY��6W5d�3��hYX���c�C�/	�W�.����B�t�ѡ�h���t�:��P�Q �͓3�j	"u�uXk���mp�+�Y�!��l^�U4i*�>e��d�~ҳ%"v~gρz�1���`��AD��I$���`F5��{�Ҍ��k�����"��sk����$k�)�_�)|S�wD��Y_T�B�c&�xc^�U����PG��M/�%�����+�o.K�"��73�hݤ�ZWQoK
�J!�X�N����h��S��WOdh��h�=�r�8�o��*f���G)�sPv\L����I�3��7��$o�mbE겅�JʵF*EY��S{�cj>��A��e#�3f�YS��z�D�R||��D�^ɥ��2�)��D��[N�n���?�xK�F�h�x�%�c���ӗL�;�,+앛�VpC���qށ��s���0Yso��D*I^6��T�͢�ܾ}-��KZ�oۥ��M�C=�h�_R�;ap�s(�D��uru� �5C%���#�as�L�f�XK��ҡvqڼ"�+���q>�b.^AsC��*��Ą^�u��ZL;���d�vAkA�Ÿ�6G����o�.J�_�P'����D��c)Z	��.��S=�s����zٟ�`W��B��m�C��+,Zq����ȃP;�r7�N�L+���Nm[��v�c�Q�ϴ��>�\z��R��	��h\�K��b�����+$Y���]i�oQ� �@�컵�y�h��@����q/�����i�tѧ�������j
��K�
.�X����&�+�{��U`R[�7o�Y���r/ѭ�V�fA���ϫ�=#Dv�r���aty5�Ȇx6�]�t�XY������h��5�����7�ک�JG�oEl�>�܎��������Uk�t��P�Zno^H �J/�uɠ㑂�Zɴa"���֞�+���}�Re0D� ���Y���0{b��mɍxg�3,����W��z���q��@��y��mC��	�$`Ҫ>�@L��!�s�\�����^b" %Xx�g�����] �`#���ŻT��N���B^����f��>x���P�	��7=y��L2�]�G�D��k���eA�bx�F f�$��Ј`�N-NW�����p@z_ɣ�VXW���V[�
g�.�.W)I�+��yAiP��| ;1��ʌ\��+��<��#}hp��A>�N,���Պ�q�N�LM��#��?s�ǟ0De�"�E��
$�&G�+��jQ���Z������eթ��ϯ]�Y�,L�4���!��\�旂"�͖�C�v�����@�X7�f�r��Bжm�:V�w{��SyeIF�==c)�#A�Ef沣��^Ѝ_�q)��J��r�7,�w�[�$�D�!��8r�-����h�L=*��g�H���W?P{��{�nV�+��>�@݂"A�6�&>��ZC�;�Ab@�H��="����G���<��N���&�1��oYY��u�~HO����&������&�H�"�s{�&�$.�r�[��Xѐm���S�5u�&��+#���L�DG۪]�7Rkc��+h@�s��y��(�\3�տܼ�d8�v�4�Ţ�8��e�$�p��܈����XO�Wd�vo(�&���������CB\����"N�(�á�<��|�֢B{5}/�a��|5�ҬL����9�#��h�Q0��Z�z����Us�0�h�ɭT�t!��A�z^Y�}U!cqtx2)Co����w�P�/q\&�!��{��)�%��g�%���QE��)��M��kG�-[��pK��+ ��%oRǂ�뭆r.�R�(�5|��Qje)�v���E��*=��q�j�W�`���e��y1O����`�����@ ��m#������̪��֊��.b�wL�6�$�����x�>1 �1���� ۺ�^��6���C�Y���_��+�����ė"~�޸��h����������d�rD��;���
�=�rLa�je�&�Ku����g�0�����"����ۂ>2�V�����MYUǏ�>��'bj޾��lHe�c����m���ro3��ßv��/���7)��� h�V���&4�{4�)a��=����i��MlD;��(��r�<�ۻL����*���̊�l�ë�E�I�
���a���'%�UC.:�E�^�1>䦨���GJ�0ST��;(X��Л9f@�*2���Pug�,u�Bd.�����C����]k���*��lWv�h�z���Pf���s̚a!n�E�˵�%�������o��+.n��*�Xΐ)�Ԇ�s�u)f)�٘ծ�d]��r�.�N�f����Y�S�B6����%q�xۆ��47�v㉜M*�������z�(.p �*^�T?����g̮�5�N�0�;B+B�� ��i�J�N��>��]�� n��u;D%V|���7P��~y�e_���)o�Z��]:��bn	Vƻ���]���+�ä�<%7��n�Fg�U�	J{�H�����D�rOe�F���at��3�J$��X��t�N7�Q��Ib-�賉��������2��@��; �޷dm��Q< s����c���1�D7@�Z�>Κ��b�*�f_PG�8'nc��љ6�9 <��ǈ����&��s<,�ŴS�Ce/���*�4�1��=�ɐA����CPR���V��f�������١��+u�`�hĀe�9��9f2-��?�@Ui���c��Mh�l3C�^� VA�W��_Ǿn�!��8�|����F�x�����R�=�4;���@ܶO�����_��9J]�\����(B%i�W	.�Gf+bI�z�=�1��|>M��Ľ+ހ�O�L�=[v�ֽ7�h�K��fj0�[)2.l��}jBL�)2�˥ѣL�m���x*Q$�_�ֹ�4��Q&/�+(>D\�Y����d�d�ϟ��)�nD�ZluTڎz���:XǪw���Q<�y~��+e����z?�w=����4��N;_ꐍ_)���b�t09/.d�GK4��1��oڸ�9�G�@��1Z5R>9�:痌F;���v���y�c�[�!EB�1:so��c���;�R��j(�Q#$��K�m�L36��:����,Rh�7�b�*'TP��T��i2@H�����x��_紂Oy��Ɓй��׋��X	��J���d��b��e(u���gu(>�{���j�Dے'�_K
 ���H."�7�AL����U�(�T�@�&����VV`�jc�K*7x2�=p1趸a��aL�9~�$3uI)3�?���½fa��)�a�2�c�G���{�� �� �K�2�=U�Nz���-����`%m �n����wr��0+���}d�O !>!Q!a�� r��>3��E�D�z8π���"��5��B���O��8/�q�(�nOv���r�x�n���LQ��V�Yk���nj����u�[A�:�L���~]�q���Ǳ&K�K^̣���b��L���~��������&X�~���,m�ҡ�O���.vlܳ+	�ƽ�M~�h,Ehn�P9�$i;���jC4����|9��jyk������Ah�_p*"d4����A�Fd�"5v|�3��Q\��ǾV `�8R_�,H�%z��oC����`Z�쯢R�z�������oNw����Y�n�7>�T���Ԩ"��X$��B��GNG���^��˛2o�<7������ke���?�yub�Z������'c�G�d���>4��G���ܿ�] �В����0��>�������)��(bdX��ѩ�B0ܞ.��2��u���H���\_�M�8�zlr�H�_d���`#QI�D�����S�KC	�r�M�6��C΃F��_r!�޻�X�1�{i)���������\>D�#�3�e��rq�&�h������E�r�]8�>CS���+^04ú�aڡ���(u},RI�������C� [E-�u��b�j~����D�SΩ�~/����NKb&�к�� �ʡ�'�G��zѡ�)�����A@�����v�NR1}�q�m�r�0�����p�@�`������M�s����kG �I�=�8c������?;\#�0�W� o�fm��}�`kŒE
�q�I���i�s+����GAt�!��S�D?ŗ�*܊�$�����r�@\�3���"@�.%	;Gq�EF}�0����B���־'���>g���g��}��@������iٖ���.WÞ��w�={���umSc!���s�e�@{�Q�����gn
�ڳ�e���08�늺��fJ!�
����
[9ZM �e�^0�ރR�e꫘����_O�A6s�������\�ܳ���c�'z(���ٝ���lot��H�q�gE�Z�MzV�f��M9�G�����"ܩ˞,�.L���1�Op)���Z�DMG��v�R���=_�?��ݛ��p��daR�6^�\d*{ٔ����ȃ�Y^:��;��̑���� �Cn�����IШ���x�]�$�2�y=�ĦΰXE�d����ty����H�1M���KflGo�n�C:�LS���`��+�
7�P���C!O	4)���)���,
f;!�(AL�}-)}t:)��ZJm%/i-�RM4�ߢ�'��u�3����1`�V*���8��2�F^��
1x4;�7��x���R:�;S{���EF�9�l��N�lx~�¾4Hdb�t������e�<F�Bvl[�ʺD����w{*T�#�cj5Q�p�PfA��ɱ�����z�uq���Hl����R+�u@T��j�G|��a#^9�
h9�ِ7p,ѫx�h����`��A��z�������G�-My��Df�:���m�<�{��|d�>8�.p�� ��'o�H�[�;��ӯY�����MP�}Qk��P�{2�Z�w�)g1� Ô �P���˝�!���_aro'L�P ˧�9����T�;W|��@��-�+�s�Q�F5;���hà�)�<���=����5��c�uK�0&��n�u[6�X����	�j�5�F$c��`A:�u'�%�Љ���=�:OE�����r��J	̏���ph���n[M����5W�C����@���5��I������0�|c��9���Z���x�rXD���v�ƌ�����Hw�&�,p�P�r�]�{��N�;P�<��&m����]��x]�TҡL�Y�k�Wbn<��,\ft��nZ��6�?�5|��ӟ6H<��䶞�z6t/
������JSI���(*F.�i�cd��j aD�
͕*Ӷ�T���a/��tF6vr�\�H�#N��c��+y��s4\'b�˷~��l���yЀxՓإ���p�lU�G
�*H�#qK>A��w�����ʌ�Y]�����^��S���� �����E"�m��8��PZK�bV�D���{,j {�SO��M����B�	sM���-���'c ~�K�x��%�h�>��+�� �;b��"$��&�����{K�P�!}}�uX*�=˺`�6c�C������O2�PSu&�g����
�7��!'�e37r�
������s=�Ԗ��1��Ɗԛ}D�v��:��kB*���eDnA�s�O�Sr�ksY��]�Z���#���v�.K�a_�[dXz�c�0p�_[Z��̖�Q���YX-Jd��1��\���|�l�w���M�B;�#6s��6�9O5`l&�����NO�rg[ܡ�#���U�Iщf�ݭ�
�b�(\s�M�$v�.�%v��He�[������߼k���֍t��8��Y��Z��f����}AW�A���Ö����|�(�j[��]�\(���o�V
��O �tl���<_y�F�=-�7�2P+��$VT���{h*�ݝH�7�v{���!f�Z���>FN�/l�����s��è�7@m�v8ja��?�}*���0H��|�2��9�s�D%3���<�ݧ�|Y���x݃�q�|	�l��q�`��q�&d�h��A�ʘ{�y�Їy�������M�:mR�+d~�+�p=x��@P�p��)��$�2���1b5���R���/kD� '�i*q�C͒���QR���vm���HG[��cÕ��v�ٺ�R��ð��t��<!��,Du}�A�Z�R)��
[��}�������2G%r�wI�����Ə�ؓ��]o�Ī��)�4�� �\*����zE�'�1$|�zao���&oN��4h�b?���e���!�Ϣ^&j`�?��
��0�D���(}�*����8�C����"�{�b���C����򘵥���v�cT�ʗM��^���d�̭�k�#}.J�U�����ـ�ݠ���,��������b7.��bS�Rǩn-0�^_x�{���j@�TT�5=Q�!��C�U��
���$a:}?	6~��ڷmTJPiv�{�Dc����Q���k#��^����!!��Y����3�'2��܏$�_�ڴx���d/\t��:0k�jb�l`�����l-%�˝&�\J��S�md$d��.Fi��RK�h���<s���c�1H��|��g�{u{~��.����f�ủP0p6+J�<X!;Up�lj���]�Bڂr��|��3`nx�gTT�]���E(W�OFYA_�!szyʑw])aѢF�tA�qHk�����?5/�&9��c��Cr8���x�K��No�H�Lkg\��-�~�cx��pl�B"��0��>�������w�:�1��a}��OM�����
�Ҕ���� �pg+�e�	27�O@�9�!]+#��n��qy�7)�tOe�'ݴ#jdz�/*nH�|�_�7~���VJ�����s.+�?�E+���ϋ���3X{���b�][�P�k�%5
�$r��� �ņ�r/�45g��}�$쾚��P�t�櫼uu�ɏ�s��Ԝ|��P���_Xr.Y¤�c��?�X�EL3<ؓ琺�Hן��e������� ���HY'#����F�=�AJ��uq��uӁ�슭�H��d-�樤��a�eP�ɯGlY����@�|}�N��)�i�q]ʜW�6���<!3�$h�ӘC�WB(i'��˦��J�!d�9Oر��ͨ�j}�)�N�m�Ғ}?���~�x����Uc�\�n��/����q:�VIV`�x�CVS��1�B�,m�f;1�9Bc���+��?G.Qu��T]�ʧ���]Z,/r��itx�;'�s�Q2��8-���92��w5[E��1.�!�}�/e	ϛj~2�:�l}�e��y21��[��Wy�*�|w�f���rJ���-�f�HL�&K/��0�|p
���"�DM�Mq��]�N�'�� ge����5��Y���?�5�fS3��ѱ
���O��5�%������\��o�Բ���8szF��&ܙ���\�[{&v~٣d��H���y!ؚN�����ED�.��Ҽ�.n�VlN̲г��4�2:P���v|��){(?� |5j��fA�|K]�?�]��!A���d�v��y$�1���@�v5���K��.{g�0���I�#��p��aޡ_o�6�8�s��Bu�Nm������~��菸��&t�r��0�B�.��M�9���1g�f��g��P�Ai#���4M�z/�wN~{��,�/`�a�9�/Mz>�Z����@l[Ir����v*j ńP�7��qeaͿ9��	a�i�5~�o�h��1J2I/����)&�v�e�b e�>�y�[W��.�TS�����9K���{�{%`;�W�I���R:;��[�*�L�n�
�y�<S E1�UX/������r��݉L:4ud����V���x�z�̀��hG��yy���|Ab���7U;d�𦬆��#�0�iU�T�	F��˴�����҃���2\��x��p�9��n�,��վ{�;�͏���X��ad�����c�Y�WdO���=��m/