��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ�����cY�r���B��HA<�����N�#8is<M�NVYwׇ� 09�)�V}�	�NӃ+C�_��H9eo�#X�)��m�SM4l�k�������xD��$�ҭR�1���A��Y"���7��!�V>�
#���R��g����&�a��ԉ;�+�C�E|7�}��(G0Fw�#"n~�B�4�����b�F���m�C�����Jwѕ��*���>�،̉����t�,����������z�}��N�3�A�guC���P
al�IT���~� ��ӊ�D:S���U�zp������$"�i!aqݻ�c�yz��/�i��D�%8+H�T�B63Rۚ��h?!�� ��Q��Ip-�AF��
a�J�#^+��6ȼ�s: ^����'�\c�h�ע7J�o�8.��`0�M7�'�@:��q|]��]�*������G`Q�!~��Z`O�x���|9ҳ�G��:�����(�{Y�ya;��H}��Hm��s�j߉%��m�����y�텿�]�ל�z!�.G���z�uB���<�Kםv/����ʮ�ש���J�#.�H��p�R�m&Z
��p��&լ�z�(��C�.����/w5�Nŕ��=�p��c��<my=Ys9�a�v����"���~�ȳ4�X���G�� �i��)^s��k��C��e&=9OR&�0���Q�_
��ػZ̆�PH���U�n>wQ�t���M�V����$r��,\2��'"��ො$�J��L����\��V�"�����a�������{_pJ?�#%[*��0|wbv�N�ނ��[�����Y����j1�����S?�X�|�*09�T�1���8�C �hЄգ#\������������F[S:�%֙�_a}k-E�X�H������e~iU]�𡁆����de+����(��-�q+�NE��O��_p�  �}HSь	G]E�i#�_��Q3\}J���'������|'�M���8B�WP��$�{冽@�[�(�!��o�_�?��vA��e�H&W��MB+��mV~픻��aE���넀���V�t�&;�7�B�� �^V��鰢}������#`Ɇ�O��
Z6��A���>/[ϓ/Xku��X�DAA	��W	��*5�V$�H�M	�w�[�Ň�+S��;��8�~��K���n;.S��|.��%�f�r"R��dD������}�sr�b�:Y��vX�U��~�ķĎ�ڵL@�f?A�t��V7y���o#�UL�:4R]|�A,��9���-� 9��(�i��g��&�%M؈د����jf/��,��c&���Y>���o�� ��z=���������cf$���IR��ⵗ�ҟwbU�4�>驫����ʒl�y�U��l��9�M2��j<=ΜuE�w�lCt����}��W��`����W��Mqo3_�����K�@�5�n	B��#6�2$g�'밎�l�33$e�����*H\)�N��?OQ�ϯ =S�|�$kr�\��?���2�6���Y���to�u��z��m����'���ZF��O��`r���w�0']���8͸���铼�Y�'a6��6R�<�G������E��r|��R�҃��& �T'=�{�A���WO����=7�����3����|�N�M�~��앙�n���(3)���X����.
J�6\_ afY�r����;�GWc�C�Xt ��N5���oI'ֽ���R�%�S'a��p�B�=�	�nHH1��H��jJ��d�(�����絾�~>���&#$X���mS/�&8�|[�c�������>Ԃ�#��O�a��$�?m�Q��1��T �J��_�ć��]�rD��j�lN
��h��"�Tj�_RZ>zoѶ�&9t�u�<M�ܗ�?MX��	��x���[uK���6�P��i!J�G�?4p��n΅�\���ѿ�8l��:cj�(��VZ "'��ٵ}��3��W]�!�Z�����z�f^�}��U�7��5��(�c��;�jGC>q?r��2_������G/}�!����3�0Ѐ�Sk����l0�vFKĂY��{�A��Iʚ8�f������\��Q>���-�2D�n$�A
��l0�cV�2�h���\O>�~ݾ}�-&��7�N��*3>�KksP�i��ϣ���C[�����O�ƌ	�[1\��x])��<A�MT(�W.C��=c&ΪQ��A��7�W�r+���Wْ����B�"���\�흯��VG�!n[ҵq��"��d�ezz�{��fĚ���!����7qA��N5-]X=�!2aqA/��d0ʛa������<�CPo�V�Xq�R���q�C��v�#�kc$S&;�įm����q��\ &�z�ՋVsᚉ)�\��*���eV�oj�2�j�?�X3"�gSq�<Z�l|E��zT\��'k�C�#����c�i��׹W���|�m��8H�@��KY��kxC�Ϙ��6Q�ώ�8�O�gi��u]υ�v)mh�e���|Š���Y*o0B��x�Ϋ7�'��1u�N�˽�Ȑ[���M�:֋*ö��K]��?�Z��A�vw���P��SHa��t9�ΐ'0�w���T�뮝�B���;��D+f�ԠA�0�O��F�Œ�\��0�D�E�l�����q.���Ua8"���boR�@$a\��c^�N���Y��7��O�_���h
�AO=n�_떝�zU�;�\���M�?o�X�F{��М����Pa��S?�������5���F"yp��M�s�,� )�Z��9jp�N�M��7��R��0�d��x$zf����|�i�=K�S��}D�P��o����k�.�D�^��o�ZO��U��#��젠���d"��ԢZ�$�{��&��x�+�z+Ү���k��XK�&Ey��nfj�ƒ��?e:�Z���Lm�L)xI@��	����qR=ܱl���X�L�{:�,�K;�d��MY�I��Y�T@���o�c�Ǵ:|Q��6W�s�G��2�KP���4�5����È��[�P��vgr�� 2Y�U5�JW�Q<���|�ޅ��� j��?�d�7�Ɲ
h`9�4���g���0I���䏻�3���"|�E	|<���o���3� Gg.�<
�o��a��	{�X��bt�*AOtͻ�)"�Di�)}�O|=��p�v�C^�=��&S�+�S�������o����i�|��� ÐR:W�ϟ�Į�r%�f��p���:� n���C�רM�ɸsS9p6����[�'�Kgxz�;j����� �.���t5h^��<,��U��J��P��b&>.���ץ��}}
�ƪz�\2v�����'?�h[q,i&"��K��D�1��u*Z�� ���&!*�����l�?���	�3�mnQ���H�}�%(�X{Z;
$��l�LRZ�$�De��!|ƃq��`Gs��#ʆߜ ~�$JN�\���>��~��\�^�T�R���fY�����b�x���Z�~��6p�`
�S��aRU#��;� �8Â�n��O!�X�kr榜6:���XF9u��&��{.�:��-��x*�~����4	����ƙ|�#;sp
�q0�b��р��a��9�H|k]D�� o���"�c)B��8�*����&ң�v���[0J����)��18W�7�PK�Ӹ�j�`�GSEW{�d��QL�2T���M�T���1NG�6{��n@�ߜ�?]f����:p������U��<C����UP�s���SK���eCs_���ٚ�t\���m3c=��5_
&����o1:&#�k�c`$A�ֽ՛��H7�d��f��.�z�xyp]�JM�>ë��
%��W�9�|>�X�c�I0�<R>l+��N?�(xfhBy5L&)��)k�ctE7w8N�H����Oj5ލ��Q�J���g��D�&ұI��%X�m`�B��8=�U�Ů��X߆*�[���Y`���v�>X�"��<��v:d��*�Y|:`���2��SoA%9W�ӎd�M=��f�� E�d�G[�@�~: ���]�ފOq�դA㒑j��~rى	�^NL�7�1���f����NXX��f�8��^D=)i�lIv�?_y�*����'qFEYn����͚�X�����/��y�I���S�u�۪|�
����蒢7�Ee|T��rc��S�v�d�,�:*�)����r�O�.k8�q��j�"e*_n�	�`�jI��6hbR;�V�,���>ǈӦ��T�=5A��$<�b��콰�^^9�￭xgu��M˕
���-m�3��������M���|Hq�Knp���Y�[�@PT���2q�5�+Y�#JB���,���.X�P�6���`�-]���D�����!�1㚀�k^��}7>�,w�iߕ��\�Y$/���p��
Ou��}!l��m���0�V���=ސ��P_n~�C��m���p�m�a����������74h$r���!��qH��ɡ������e'H��}��8oЪSb��.,0���`-�݀�v:���a��I^�ִ��u@�!f�A��P���D�>�s�wI�/�
�ڎqW�6��:r<K������~�<w��-�Z����t��T�S�xj(�4V�M|hAm�&���L]��4��L'
I�l�6f��D�蚣�.zxwv;����8Q#��v�`���ǛOi�OH���~��q�.Վ��-���Nr98;������v�l��uA'�>�G�n!HW��nS��ѢMآ�5��y���ΓMJ3�?��7��h�iE��+����P�s�lt�Ɏo���rRџ��Ђ�����E����H���'�`��Z���~{OĆ{/s�\��t���	F�~d�Y�%z
�8%I�f���kzܫ�h��%��㶽6M7�S�2�n��I�=,LdŘA5�#.���0���r�͈t�=��ŹK����h.���>Ԟ�>po����בi]^aU�d�[�,��Hf�d��!Lr>�Y�w-+;6��c��mw�%��I̫�������?8�������������$F�
��H�o��s�<�̿c�φ`��wD܋ �௄v7f���5a�,�>N�{򙞎�C�8fO�t�_ \Z��%W*#�"���&�z���q.��1�ތ�R�M����1(�ޏ!+��hǡO� ѥ�����UG�e&a����S{���) �ێ9F�i݃ѻ��q���H1�f걳L���T1ؗ����ܪ
��w�+�#̮�/����>��^X����'LX6س�ȳ������ �TȔ�AL���a����!6ƜJr�K9�:�ܶiҌ���@N�(x�%����U/�ۓw@�n�b�B,C��EĥEx��,�N9G�����S�3����/arZ����(�t"�a
v�Ɋn�.k+lhU�T5x�G��?�=�0�vC���D�N�/t��jW��T���k��V 3��y�%���L�ѡ3u�%,}jfN�<r�@I�c�
�	Њ������X�k��1	�ׄ".��$��Y0��tk�	!�eH��0��E�f�orI6A��xn�.�c���L������&��y^u�h�c�5A�U�t>&8i��s��/�B��
m{��R�G[�#��h(��w��ym��*`�����Ǌv�r�87t"�%���D��VŦ&�&�y���U�+����/Ÿ�U� .���G��ڈ�|���qì+=�����E����ڇ�S���I7tJ��,/��qn��O��a;s?�I����I�G_�#=|9JΌ!�Q��2��%�A��	n�c�0l��&�^�:\"\#c?<��̫�#��7�,a��}�ؼ�Щ�&�:��1 B-�Wb֖�j�zr�=���W%2�Ө�GnzBv�Tz�������A���,�)�,	�D���r< 4���j�8,E&�[��������1�] ��d��W�!l,(Ҁ��S\'Bx������>aa[i\�	j�F��y�,��i��jr�0A�>��#��	[��wu���*��d�[^A?�l�5�x#ѕ;���0:Nx�}���*e1��{��=aCq��{�B�+���y����$Z������Gm�&@�x@�~Kܘa'�����/p�9���g�5���@�����J�O�+���זI�"�w�8픅�PW^��Td&�cЂ�M��d�4������U�r��,�@�/�
r�^��j���hd�h��I�^J��?C�,�Qf�z-�W�l����-�7����c��o�#�/�Z�c�s�2!�����{�a	��.X�'
��Z�O����a#�b�����nJ� �g�E.98h*Z�a�������Gk��2t�+[�Ủ�H��);h(�yM��:&��$��\ �[��I�;�Uog;J@	X����n�eW8s��q��,~��v�'d��%��6�1����H��@-�l&�L�2M��o)����G�v�l�?9��F��=�6��ϰH�jwĭA��b^�j~�q:��=HM�.*'�Q��X�	�B�)�"x�Цuu�0�ޙ��,q��4t��.���L���^L$ss��/ޮ?�XEu1�d�M\O�D~��V����O��֏�^���aUn���5ڠ�([ASP�>�1T���C��B�m8�E�����+�F]��G����-��G'�(c t1E�+p��^��ט��x�<W&�.��.��oa}$.t�O��m�7ad/�1��ݺh H���0�h��][Է�k�L�Yu����{�Q�4�

�8sF~هٍ����4�6.��3���q`[kw ,n�A�� w�: ;߂���PR̾b��p֥ۀ�B�H"�e.���,�f��S�d��E�&Ѣm�� �B%�|�FD�i�>��T
��ov�Ͷ����*Ur��?���$�"��A�S�*:I��y�9��7G��dR��I���`H)���+�|���A����t��w}y�F���K��bH���Bjfഎe��HX�� �l�٣�����B�F�.�ΎW���ik<�bsb��>��GD����3���;�����*{D~)��L�e~�ےs�(����ɑ�a���4a�2	�cc9j���4ʆ~2Sn��S[I9��X�d�!������c�n�ߌ�����a6��Sg���<(��`�����崻��pA����c�;�\������5�؈��W�n����|������1`�2g���WV� �t��@||��)%�@;Rwı�����Q��3�G���ɝ��l�yzl���֒Ȁjq�Fƨ��l�l$�'5C��27F��ˉń.b>H��lnڌ�rV�;ፆ���=H3&���4�hKL�F�j<
��d�8]�	H�gg�*X�#�p�~U�|�05�~�Ƴ<ԁ�w-N�:hW���}Ch8'�l���p%���J�4�H�g�eg�g���`�£'Iz��I�u�T�$O�a�B|��R��a�}Ì�ur"vTk�p��ow��^������<5D�#�v�mh���PO�dG4��[,|G�+��L̷�BG�]�P�����(rT���l~�tz��p]��Z�֮�[v�7V�͋@�,��R>5{�:�Ш��(�	3:r�b1��WZH��4�{Ҿ�`E7���sK1_} 4
Y?�OV�݅)i������������;���4��+�m����=���*-qw=6��(���Vy�_6}x�Fi�g�N�)ݦ )�8J�"������Y&�ز`?�~��7P�5���ͅ��K��%J��Z�����Pa��|�x���wk����e����Kc��P�4)"��R��c쵇�#߸ϋ����� 7V�*#�A�VZ�8��7��H�f����	�_S���cU��C��pQP���xu����pc+y�]MI/�p��X@��� ԎBC�+�_T�����juIO蹬��0�����m'E�F�v�>�HYL˾B�X�7�'$��E�M���^�;��Zirs�Ү��s�Yvi/�ª�hP�B��#���Yyz�k�s���'��Q��Sg�3�}!h�:<<x���E�@g.ZL�ۺ@��J��I��xz��Q��d�H����2t�H"tYo�rh[2�E{M��X
x^����Z7q��oxKp�W^�BsW�RC�FR��ī��g�$��a�Z���װ��'d%M�+Μ?c�J�vU;�1�D�:��3�ײ�,0�CO"&m%UĻݣ��yt4.��Qg��ϼ�����ȡ�ɔ���j7[~��C�=%}�
=��Yi\C�����O�ܓi�"\.OU��?D��%nMcHF%�v�C���7:m�5X�OZ��H��.`����>}-h��;p�����XF��i|/�-Q>AJG�
DӞσB�4�sޅ�%&�.������i�S�#��2*����"|��M��kS�w�O*d<(C�����0��\�LaRȺ���N�uʞ���#�OC�)(�����2�����~ƹ����UTv�j�w�l�>!!ә@sklq�1��"�*(k3/
N�#���0~��
��nӑ!��K�Z��ny����q�î��遇0��x�:��ͬZN�6�����l��)��cZ
6��MSa��B���6�6xGd�8db�������j�Ju��6�9���~&���A3R���q�R(,��K;���q��*~��U�������ܷ�����v{?ҕ��[=7�J��W�_,۠2� qa��+�� ��PU�.�L�EY!�ym������D����9ۿ