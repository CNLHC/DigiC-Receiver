��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������FuZa����cֿ���
R��U�����S3C�G�*{���c0�R�IG�b�`x��<H(�a��.��pVIJ���$NL]c��>/�lN��+փ���^�>W�7y�/�]���Dh��>�;�Zۇ��7��A��0�����4�!ub�0�ɑ� Y�
YY�����k=T��S���?��IZ�c �;��?`=��u�|�D��ul()>�,�ѥ�p�[)��;�cn�a_�ouNf��Z矟����ר/�\��`��+�̾���{��k"�%T�K����M�w#�C[��L�jA�����S�qM����S���j����N�E���}u㛯P�i�0�SvҨ����ĳ�`��G���`�L'T�'�'	%�|A#>y�h�������e���*o��C����/��|uK�0ޔ��"�(����Z�2��	�����2ZW �xiO�C����xc��5�f�
����[,�͵�$v��d�p8�yM1W5���"�s[��m��B2�����@�j��T����IӸ��p��1����g޹I2�,ر��w�W��߁׍������V;+<�YGF��]=:S`�K!�%}@c��sn��<Y�Y�f���2l�����~|�V������*.�N���/|��|\̯��gD&�|���enJr�Yhc��l"�[U��B:��D�J�z�P��QH��R�'p/Β�0�I�[��@�{ܦ�$@)������gZ�J�)�a��iIb~m�4�u"Զd�G��C����in>hOK�9��z>W����_R��M��`����{�ae�b��:����a<@l��`����r�n�~���L�1���#n��H�³��E�� `K�t;4\%����&��̕S�L2	c� f]�t1�#p�|�1�d�����)���, ���V_�4��~)c����0�GmWIW��̈h�{� ��������A+�A��H���%��F�Y���Oe)��.�����'�@[���P�k���p�.��a���?�G��/���ڛR|�nI�j J�#��;�H���9�W`1��:��Jlz�2��7Vh�U�ѥC�㛎��EB%��^�d1��[��NJAΡ�4��K0��^\�?Y���Rmp,d��	z�2������I'a��}92�`;2p&��Fs��-C�$���i�dي*K#ߜ�F�U蒹�؆����RB�eƣ|��>=~�&�e�Ӂ���f��IJ#�Ĭ���]��c�x��,����	����Q+|��;基�O�=6���]�l"| �~1�f�]���7� �>�V�Z�-4e�~�\�|���G���R_����p]�J�C��`�t�'�Ξ:A��߸�s�c�7YM]���X�r�"��f����`vt����J+A������M�D����[��>V�W���I��}	�æ'��}���(D�D-�p�w�OͿuƖ���}��9pFՂ���H�&�
�\���h���_�F7�E�ό��H��W+�\N�7��8(�HsFвy���WM�s���0�Û�ni�\2v"a?6~�\���1g�0le��M����R�+������ ���'dW�QI|C�ŷ�{��ゑ
b�PL����+�h��,����U8c��1*��ֹY�%��0���8=cTV�C��#z\B"U����A��A�7.�^6l`���@����D]�[)����\Ը`VSR^��6��N9��g�Z0��m�EP�]�y䕻��Y�9A#�Z��g �dX��*Q��[�h|����5��H`�oѢ�����񀜜J0;��LV�T_���(� W�T8K�'��ލn!�'B�n��L>�$��3qکv���j"+sܒ���aW������Q�vl{G{i�L�F��>ŬJ�g�e�3g���gå�PC���SV��ɖ�;~��k\�~&���d�+|}�:�o�4|��n�BI4��.
bH�l����	 1�� @�M�����0]!��g��������kɿ�8�����gӁ�|��<�T���D��$(N�V��Ŝ8|��)���66�$9_T���̇��F�L+�L�2'����Ȏ���U4�}���
�l�n�r����ˀdԿL�=�G���ݘo������Fw�{`���	���E�(�l���Q��
�d�90����M"�(�=�Y�6��j�φ$�m��<�j���k�^cyTK�M�£�Y?^�� &umk����p۸���R��J×��\TC�Pݴ?�q����t�w��@��	�!�]"X E��3v�j��9�v�^(�T,Y��^p��)i�C�B�|�fS����{�>g��;<}W8�i�"��׈��&�B!����l)i9!V�۬O�>f�6�:��/�M�Zc�X#ڬ����7��R���5�bo�����H����`���vT'�B���*_�r��Tt�S~��~���~�A0��#V�bh��d$���ϲXll����J���Y���&C�?�(��_�{��Ӂ�49�����^�_�4�D�")P�!���M�Ѽ� lU�[j����O���x�ep��FI~:@��ZY?�b��h�AlqEj���1~`�|a�YڦH�"���j�L܃.:��`a�h<'ԛ�|Ri�������I��W��Nq�� -��ߔ�w+�jÈ;�/<�7���V�%ߟ�bJ^~ꙸ��-��Io�����ﻓ��C��e��|_�$��0
�0n�<C��-Ξ)j'[avN��2����_]Q�9��GPչ����ݎ��vF_m���m��%��3 �lQeױ��R�+�t�<�u�|w��lF�;;��:��˞Ot�\
�*��]�~rQ�b�pbj�4ɣ��	CEn:���i�=Rp�)h�l�nkx�\Hx<�������7j�
�X�|�A�U� ˲�5�)~����~w~��c�1�����;8�n�KR܏�-n@&�;��l&]��&!VT��j�O	���#���.����A�? ϓ|�6k��c���y����E�~�QS��a�f�e��������y��9k 	AHs4_�DN_�Tn�Մ*y,T̕*܏���JrY �ҞR�S�O�j~����)$#�}�{<}�C�B������G��p�A����i��b)e=��	���P�������q���Qcfv�g�6uHyKR6a��Ù���-!��b����Jm���%�(JM�Bb�J������k�6:��M� G�s��f�-i��M�;�S�6%��"|w6���a�<~��&<4��L�^�f�N��Q�95��U`@OSK�e�s8'�yC����]��:SEٱ�{Gc����.ݣr��,]i���fZ&���=˟���� �V� �&����5�,0/�}��ܱV@��J�Ѯ�,�i{�����A��@�
{���|�C�_Nʬ�&��pf�i9ެ�9j��,+$6�/�G���t��ǵ�2�����6Ƙ^��7rN�A'�uOn;��K���tƗUr��	�	�;SI]�
��57�!������P�f$|*�aR4Ԁ���m�Cɴ�1d�ʅ'���u��j�O���_����΂g�0�"���z%�Фx3����w��\~�4�wJ�fK��� �i ��_aR.�2�ÊG;�{���q����>)l2��7C�q��,
���B����T0���kTE<+:�\�.I�R㽍cx��>��|�Z����|��{7��i���ڇFW��cXL�9��?Y��G�_L�$Q��[;d�Fi�P�$3P"P�_�i����Ŝ�B !�S�
�X��:�m��H씞�8b�E�$`�f�H$OE.�F�ɵ�z���X��4q��9��@�;��rd8�P���#?�z�`�mBZ]>l�/��#����-ꛩ�� ��k�=j�]�$�@V��h�^w��c0Uoea�Z�;kS�,�e#8VV��^tHJW�8��C�Q9��3@Zֈi�P3q�%��^�RQ8,���,&���:�s?��^3�?�KZ˂{@W��<�Ykv�����B�5���+�9�8�<"Ctd��^�ؾ@&�L#�f{�oJ(j�,D\�|���Y�q��P�$&Ҭ�v@���