��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �'�(�٦����6M^� y�N&�hM��\�[ʘS���Z���)/r݇�?*x˯F4<2>����NM��o��E�/Y�tBR�S��j՝�ڕ�!</
]ٷ⟯%��%Dq484)�gL�A�)L��@!h�xr�m����y��4�QM�DG�!S$?oH��;f Vl^7LK��rC�W���r�-d\�!��Ռ딂��?��m�-5�I����'sȘ��q�Gs`����c��� :dk#V9K
�D#�n���s!�W�V�#�>��Z2�c˃�{��d�XS_2��z1�x7�ζh��S������I0���<���o�
��Q��)���aZ&�A����x��Qn��ଔ��*N/-1�<""'��J��n�%��g��8�Z��п~�>nGy�mY�؛1������/�n0p����G�A/ܯ}��k=u�KS��o�hXSu�}���"��{ms�s%<�C	��FU�~kY��3KIX˱��-�ײ�9loG~��8���Wj������[�'���\��T]�+ʕ��/%�ų��!�ͩ��J��w?@��Fl�r� O��l������9�3Х��O����ʆo�����
<��أ�F�V�Q-�sv;L���ɟ�f�����oX�4�	�r�Y��+m���.T�j�i�8S:H������{�g�1Y��=��:³��9;[U�$����{��#dI��q#�U��ǿ���c���c��`�w�rE���U��r�J1�}qo���-��~��6��ȅ6��< �<�Bق�zYe�N����B�U�҃b��aN7"����3�'�@�s:��Ծ���̿��Z)N��(�i�"-[R>�DQ[��\ NB�Hi�	�1gi���L/��=����G4�%�٦�&	�'Zl��Z����,��څ���X�x�,��p�Aɢf�o�_w�A���?3-H����/�|H�Z����3�(ʋ	�`B��u���TA��E�vHڱ�#��j~��-�ˀ�*�Ҏ^�ɛz-^&�P��Uꡢ�� �Zu���vyg�.뒅�Cw�=�<�m�
��<K8���褎9;�[g���2u�L�R��s$E�8����J�c��D��r%0�Kh��]۸Fӡ+�K���$���n��HAVJ���N�V&�rLj�]BBF��Ae�g���aϞT�I��t�H�pҧE|_}/0�x����wq�g&�+��<®v����%]֡�ghK6f��)[�adb't�B���/�?�ibbF�����\P0����������C%���x	%��@��q�`��r'#���@F��1�1��o�G�S-R;�W�k6ZR� a���mx�],}*�h�r�d)�j\}O��A�ʀ�\s�>��$��ϥ��:�6��N��vI�nZ�C�CXP�c���sF���a����~u�	z*��-���� ��%얕���O7�cG�ڮ��	�S���վ���''��n͓�^M�$"�٬ �aSL�����d�8Ij��H���Vu2ے�rQz��ŷE|�>#}R��W<��Bc���PG�6�5dX��Z ��郌4��K��U'cR.�6�,�.�S�N��[�VT�;��/��e�h�-�����>�_.��@��ֆ`0,� �����R�-8��|bŕ܊����/�6��nS��� V$���>L1��t
>>�\����U���<�2�s|ř�,3��u��}a�J3�
��kD���="Jw�e��qnp���Ә�$]���vJ�@��ȡ��Me,^==@�&�e��vT�/ߡ�5�(��ŝߟ��b\�#��x_`�O�eb���tŮ�~��ʹwK�
�T��3uR:�f��];Ɵ'�3���d!9q��&!d����r�^��h2<��L�h�ͳ4���t��y޺�ܸ����`-d���祦bڇF����D^lϧ�BF �C�yYvlԞ'���L㫥����:6�X���Ό�ы���� ̟ex	��-����4�FI�4�����t����9�}@gj�[�U�d,�Ȧ��b8�SZ�:�nYhU�#�T�S��@���N $ͪm�$j�q����7eߎ��Uўuz��rml�.�86��߉��vx0K���ǰ�S�����1=v��I����J�z�ׯ��d�t�����X�E�R�u�d��q����^��_���Һ�-�MQ��S�'�?:���S2���;��J��m7�4J����aƲ8(��/	v�/�޾rFV���.�+�d6i��Ꮲ׌����[�<�:�p�9~>B�6���m�);¹Y�P���:µA��p�2���ݘ����u�X@]gB�6S]��m�Nt�SGE�%
�[�G]�]s:v������X���#��AH��(�	�B`%lE]�-���q;�)1+��}������fh�&�1��MS�l���󢎃Y������Ke�
���N?� .f�A��wp�x\&��9��-�'���q�s��	�{^��_\�c�y��7��ǹ֗�X.g�A���n_�=#{�?��Uv���/��X��N��>b#Z3g�@6��������r��	��NA����%s��I��b(p�hE=��<�'�p9�����x�*�yJ��3����6��"��K3}7�N������̂kת��ǌ���n��/Q���x�*���7B�q���Ze�SG����+0u�g	���㋵�i�> q$8춼�������͹�o�Ǚ��$f�p��W��'%�PC/��_��_��� ���xs�c3)��dϐA�ў�z�peu:�
��������R��>-h7��o�փv�&��i;k���
���>]�,�U�9i�JpX����z��w�w?����e�Ӵ/';WP�z�x4ݵ|G�O����əP��3lq���	���߁ut�(������aIFчX�S�}�9��~�ĔAl�n�x�z��a5�XL��+�*�l������1T��|��� �����_���J������H�z�Z��?\0��BkF�E�=�Sa�/^?����N��d>T0�|:++��*/�f���z+0#�E���x�2�~뗽{�h{��,O�q�"�s���/hݢ�ږ�!���S�hWܗ�#8��vt���rC���Ἑ�Q�?�X�؛Rۣ�i�v���}��	���&��:����s�m_�*�ؕ���v���L�ﮏ���&�^�����Ɍ!]#x�zQ�U����V d���8�&Nli�����o9���+�f�?��2E`�9X��W1�z���/.oI�[[v`J.���ė��nIe��Y�ђb �Y���c�y����;ͮb�L"�����t5�\�~;e�RDo��6���Μ�~&\��m�p��'%d�R�.r�3p^���Z":��������X���d>��KVXi�0��@c�6p��z�A50��pKn�;��]��T���l�=H��`�������Q��ȸ�
0���Y�5�m�1�?���s��8��|H�L<b��{�Gp����lqE�Z]_NX��]��DD:��	�'�s�tæ;��H%\�_w��q�)�}cF�;� ,n��Jޖ��)Ȑ��sg9��kR�r�0��l�3��@i�)��"L��/ K�@읯����|L$������&%�D��x�tK�layi ��tUdW��@�U7��rJ/��]�����} �=��k}� K�d��u�od��s;�<(%����F��@�N-�~���l��}�I4��C��m1HA}ʴn,'���ɝ�y�٫^� t C��]�i��_����*e�x�*�o�)��He���>}����}dgŖ�zu5��n��z��`�=��@vq��fɫ;iW>?4���z���D�֕v��hI�H昫�'�KD.W`��{^�����g���.�:�,ŚQȖ) ���F@q�l]rx �W�?4�ע�σt��� 崧�y�R�*,KdR��<�ҭ�a�R/�X񮟊��9A�'���֡s�1��A	[��+�X�g7�/3�'42����3	J�T;�h���jJ!�u-S�oCFRp��lO�f��8����	_��������B6� *�jU�9$�l"�6�lx&`Ƚ����2i%�\� ��}����`H\�w#��<�}uMB�����Cd�!�j�R��9Pu"�2��s��gK�1I���PT��f(��f���0�)�k�=�9��;��a�+kzǼ�|{��ĒʽBW	�+b�
b?BL�٠��S!㪸��Ʈ���d�K�D�S�ձm��;H\��x �RFK�>��=w�:��� /��{��H������hL;y�',�<ŎfU=��6׀Gװ�g[ �g��x��]�`��z;�+�-&l����Qǻ�)[Ɲ�SQcX\�����Ȅ"|�@�?��-!�/NvE��:�傺�<�X�Tv�B���m\��mC���6����8�_Zu� �
� ^\2����r�ud� `c���q����X�����qk�p�}D���1�	+��۱Ǵ�y9�| �:W��9O�fg*7��%�h7�[���N!y)z菸�>���E�\�SN�����◒�L�k@�M��Mnc���t < ��s�\��_�^�yr:3!g7� ��C�ã�|c1/Vó V�i����M1hJ�vz�B�/F�N��w�#8��c�5qh���������~Ūj�xr]�%1�ʹ�7�"2aj��sǡ,��9=�XW�)�d8��O������I��[��&��\��R�e��@�j	�>K[��a��G<^�$M�� �F��`c����"�0	Ȅ��l�_�JsO�����bV"��V���R^+�rR��8���1�����L����q�ؔ1Bnv�ӛ⿒e3%ɲ���7��5����vF�ˎ�}�צ����q�Sl��>p�7�_�,��q��G�L�����a����Qܜ!T��ySΨ3O3�L�/���ӎ�t��g�/��$����9�g$^�+��A��̮�^�ے(<�K��ⅽ���H�F)S"�l!��]H=�* _U�*�o }1�쁲�8���	�1+*�pꃐBJe�ku>0���3��efm���bd��1!��&�Z~�������kW�$�OX�h�,���z��/�S���^$�/�<���PEH��1�9m ��w/�C&�F�v����lx�OF����,�)@t���9������X�-�7/�gR�`(��8O<��eI��:���X���
K�C��>Rj7a^�bMNƍ��C�:Q�R�aţVyy0]�\����6��z�aH;��W���s��:{�	��/�ӫlM��ً�q��6ˡ%�Eo)����ͨ����<��Jʻj#
�l9`:}��>���V��_�g�Jt�/I5c�6�J� �#����j��ہxO,�\Lo2�dT2��2F,��T�qF|�鱽��sQ�^�C��"W-�Z�B!�w�f�h��2?a>t{l�K�k�ׇ*����崝NK�"Ʉ
jM����53e٦/���\���,&/�T7�O�iy����L$ga�-�M.m�w�e����Y,ѱ���p��48���vu?z �Ue�� 	���95��ꄞp��n���Xx�&��2�ѽ���S��٭�m�E>�;�Z�s�@��2m踊m՜]�l�����F�Knۇ���g��*Bak$�jX1;�A�~� �Qk/.�����f�x��O���Z��r�_U�Q�Fvڹe��� D�u;L]�!�+�X��6/E)�gZsʧ.�W�S�T���>��/.���)?8�O�kd�B���ڼGw�`�Xb��Py)NDz� ��f7y��0湸Й<���l��Tn|y��y�g/�E-nޯ�-(�y�N"6��mj��o��P�M��7���i��bS4�s���e�cq"k{3�e�'��DU5���a��d~�5�Ļ3�%q$�e7(�<t�~T�Ӝ�8��55~X ���1��y�O���$F\r����ŀq�,�m����&����`�:[�K]�q܄h�n��GVgc�oD�T!T-��mGb^�s��D[���2�}����j�%��ݞ*trZ�Q�I���_45��|�#}���L���:���=��q�L{WQ��Z$�Ö�#�؈{�w��37��1�{���2h�^�q�B���oO�Gdx����P��RD�0�nG��M��/@�i�T ���'<[{o y�5U��� �%q��1QuH�~F�a��j��
@q��B)�X\:q�b����7������~@:� �?C�#��5(�C�LB�xv����{�c!0`a_�rbt+.f����q�㭾ַ�
�	�b���OG՚):f(��e�+��z$��aVA�@K�z���W�����u{&� Kmk�������N,$b�}�me��o�A c����O��Q�-�X�d���Z�阨�����4�Hr[#<˒븰g'��.z�	66gU�!��UK�a�Q�?^&''��ju�����t1(�p�'��H9�ɬ,�6�9����S�bi�U��h�$K�)A]{��D\�����7�V]�!!����_�c{NAP(&N����b-���n,y9�ű$9���H&m�ot���֜��2)��B�`�����Q*[}�%��O�0 ������3���cJ�����G[�a5,r|��#zXydCb;�餧K���6�n����4��L#��P�G��H���g
�z�Ư���������ҵ2��.I�ԄvvF���e% Z��c9�AT�͠H���>�C�ǃ��3�LQ�J��-҇��R�}�ib������é
^�E�c���m{�̈���p\�_�5 bv1̣wBY���s��P�q{p����U�=��� Q���v��^1쏇�曡��cp���6.u�*3E�#�]��@_|�>����a�a������>�N:o�;0�fqCx�d�ȈfV��� ��;�TYԚF����C4����f/tMW��Ruݴ����𩠬So.�Ԣ�M�g�Ӌ�?�)jC��:i�|p 7 )�0A#�j�CG{���	�nq�qW{� �-\��׺�]f|� 4ʜ3�J^���JcJ�~~lȸ+�F��ħ>��q��{��ӪO~���K��wXx�&���#R:���8��h�o�g������P�0j��!ǫ�
�/:x5��dX��x�&��镟�{9��#UR^LDb�=���S�A4Z1 ��	�R8��Pe�<C]ǨSlX�'�e(���_
���e3܌s�ts0��%w^��L}���
y��Ɣ�ӧG
o�>�� �;|�C���
��ŵ�8pQ�B��"�vT����<��M��)ͱ9`f�Fy3T��	/���;��,�Y3��@|y�)YION��'#BD��P�%�9_�^�#�T8�L�#������"�P:��=l�Bd�C��B����J��S���I.�<�f	��M�Ok�@uv.�J�
�wPـk%پ�~���9xZ��·��ʜh�GM���/u���>�:�շZ!��rƜJ��٪�@�џR���8�ҙPT8,��/�-�V�"�&��ϼd$���P-u*����|	s*�Xd�J����Ȗl��~C�6�l�*��C
�p㞩}����)�V���ܩ?�nI
r�*����(�Ї�a���"Y��E�D�����ٿQ�U�m;V���Պ9\W��_��@�H��Y1�T���K+�'���=���U�!�j|G.`Xϼ�ab�jĊ֣'x�;���o	�&)��������!0�?�<�&
�����ݮ�w��O��c'�f�����s��B�$�\_����$6�n���"n/��p�Y6��l��/�4�6X%he��/�	֏� eN�C� �ůU�V�>��%Yw�ʛZ>Aǚ?�,���;�2N���E���� .��E���Kw'i>��fK�)�@=6��`m�A%C��Sx;�����niO���?���#k[���"G&4�nc��i�f�D���_���� ��"5��	j�#�:VA�$Zc�Y�W��(\���,!ǋ]��tm��+4rh�P%[���@d��:N��r����D��G�͹@	j���D�a�TdH�p�=Xm�����7� ��"r��ZAd�I���o�,���8W���:s��+Z����Zq�� �p�_r�9�흢�Ja�d{��ztX����P�#�M�>B����W�>*�m'߂�WY���\�A��8�e+�jG��D����7!�E�i�����cS�J$�Ǣ�@��f�(˿���I��̹<)�F7{\��d�()�����b�v#�!ɅR��u ²^�|\�}g�ѵ҃?2k0/����}����{�@�K
�;<^^@ݰCW�&�NG33\ ��͒]��A1kw�s�_[T��G9�����^/93�]��$$yc���:����`]}��)�ͺ*����pa�!w����.�� z�}y�%e�'T�0�*A���SjQK'j����m������fn���N����g%�*��o��g*��&=Mng��D:� d]�����΂L�A�ȟK(o�]�N��U��5|�� �z��ٹ�ߩ����PT�Z2�I]�Y(m�BX.��[3baj�6$M�vk��K������F4˙�;�vެ�'�`����Y�lK��<�?��<~}�	�-J�Q�/�'߸���H'�z�/�ސ�<f}�5�#ɸ�Ѣu`��`;�E@��e7m���ۅ��� 5�7�y�l�(�����6�84I���¨�@[;�d�sZS�YΌ�%�L��������B0���x˵C6���w�ʹ��	��"��L3#3�P��j��\�J1�'~z�˻Q��3Qk]��Т D����L�=�	��$���>��ﲫrH�(��8$ًw�=�˰�/��Ze�WA��C��u|�Wҿ����5[.�1	��_�\�]rE��t�~����{����K������:]:�fQ�ʒ[ߎ☩/ 8��v��&�옐��i@5 ta�Ĵ}��i;~|tʫ*2���%ir
`
�9#�pTh��AM��u���E�!�)R.8�����$���Fߞ[T_!Mj0���@�}�4�� ��%�0F����nB��C����R�N����i��U:&�Ѽ]���C���z>�	�T�	��Z�7��v��s��a�ﳜe��l�t�\���*�HL���'8|.�Z,41��g�׺���жq'�+/���|64��\��?J=iS�kE)�!��n��b�		����?�"�n��7O��wo�mw�lry�!�^v= X��HM@oɫeOcf�d7��#%j��ڎ1Vǧ�=�ث���ZOOa����X��q���IGW_¾�i<[���d�ǧu|�f ��g��Jۂ�������j�����@e�R����
]��5��Y6�2��51�r��5�S�F�]V �*�	���{S���Nć�T�5k��h�ˬ�����N�i���cxb���n��{���w�Sx7�t�����k�)���G�8 ,�����RS���n�7vJ���/N�4))�|�'��@$��J	�FB�MV!���#z�)%@�"xwF��*��tqm/�Ī
R�0G.����k�t�^C��%�v-������%L�1�Ӓ!��k��M  V�M������f�X}�z؞��pҮ4�Vo�\�r"⁹��q�' �	o��(D=�6��Na2�ߢ�_��9���*��P�����R#�C��E���ί��R�s9mXC���n�e�E������̝��a��[w�%�i�T&����%��:��;�m��c=�����ucsD���\��(�^;&=sLI�na7Y+x�3dR�.��b[����nDb�<�V�çZ�-�0�Q�PI{�11��ݰ��U0:�!aVXMpianz�%;hw����ʀ�q�&{Л�ͮ
=�Y��.xG�燄frʿ��Im�\��]�}�����5��=s�]��Coy�������-�Q���pJ3�"gF�ˏʽ��c�z���L3h˭t3_6�S�f]�=1,�;�	q 
!!�V�c���pɼ(c�zg������r�v�}~�Ĺ�k ��PaS�$0N=�P�M�s
,o��-Rq��S��zw���:ǖȹ����D��D}c��x��B23V�Q�5S
8���U�y�=^�.��H��a��fx�xy���q|�y���ap�9ڟQ1�y�N�;�w��L���4�M 7g5-Hj�'���AV�Q�ZO�ĥ:c`��,@��E��y�����~7u�^;���;@�Vg
P��l���KP(%,�pj�F�3��;Fd<h����-���.w��OD�-�d�،v_�|�V�����;Y��)7sM�_�li�s�?�` Ek����Ѭ���]�x�q���o[�>K(����*�T?}e�X�M@�æ��{��]S�jt?�=#��ֳ�@�����>�Ð{X�y�6s���:G���4�7���T�e!�f�a�3�∥�g?d;S�����up٥S��w��W;����}C�#��0\e�b��6[0���4{~J �/�|�ѹ�s�QF]��V��(����.�i�1J_:d�ۺaJ�!m�����,%��b ��Y�]|�ơ�f���i�@eO����<��C�@Ε���8p�t)�.��>��C7Q �sE3W<.Ȝ6G�K���z����:$o-��E� �f@���t��Z(աU��L�ʛ�WDh@��(2����������J�����ؑ�P�?Q��[���#�������[��6Bm���79��W�J-�[��uZk�>�1LX�h����_,M>�[RB/���*�a�/�X�*�K
��G{�`���Q	� �a��/b�ci�2�v᫚����#1�QSӨT�B}���/�m����N8rP)"h�<�u�^��[6�|N|D������]w���'��b��ؤ�
�	�ZAXN���۔D<}���G�S"Ջ	%w/�@��ZxQ!����^}#Y����,-7D_�X$���g��~z7I���<�d.:�/`v-�<h�;���i�/b���s`��SK�Lh@{��"�r��ˎJU��@0����ͻ�j��%�l�i���}?�w�N��K�>j�3���'��x�Kϧi[��wE�]����=�����9������͢c��ۑI��ٽcܼ���A-�&��1�?��v��\�9�V�\�޿i����הMefs�	J�ܵ�9}�`A�W��k{"�����ōV���m#����C8���O��i~��s�2lɈk>���d��,��-Q1�Q���7�t��
���W��0��J��IĦ�J7������p�>.T{�"ؿ�F[*.�Z�5VQ�W/���<��44�:��C,��&�h����6�E�N���˩�z]���%��+z��>��f>�	Rb��+C�b�>"��iͮ%Y�@�7�\��O��*a��� )���� �/X����:]y���G�"�-<����|\$�/�.��BlKM@��'��4�4߹g����D��(8Ur]��B���ĳ)�f��/�ѥ���kR]8�m�w0Y⩐���ң��O�3�G�� ����գM��{�#Y���+�m��0'��f�7�t�\��^؟�ʷȚ���XRV��{��q�O�4(_�����XF�*%�������~�Ō|X߆*�(;���<�P�aHm\���!��Ě	�`V��L�?W�b(?��U��[�4�{�,��j��bV*�H�*@SB�T���
Y�$��W��G�˯�'��bÈ*^7�STm$�؁q�BZ��]G?�lӺ\G��3Y�� �V[0}�U��{�w�@>Q�XѤa�����w�v-boV���$�]ɍ�����K��}��R�"��;Ow��.~��4�*�BIKϨ"j6Δj����|(��/��#�2��q�ܽ�R�Z�O"s+J��J4�gp��ӯvO+��M%i���A�>�[�Lʖ�D��0����ts���r��03�͑�ɦ�m�-�Y�8�f����1��Xz�n��ʑ}�S�;�l觋�G\t!VAu�w8�[��=&m�֑�k&n�9�f)P�j0U��Jzo�`d��r>���=��GblIi��i����M~�6e&�苯�W@�0zN`ŗ,2�~-�bnX�x-3X�=����ʜ��������&�$*T�w��fߵ~��O˝��D�C1�\�'w���#���~� ��`/o}�d_e;����� ҹ羣!�TK���,��)���I��+��Qr�U����'�&���w�3�ݿ�2Z4�CI����밖�N(�IХmRƃf��`x�}��-� ��t���e�;�Jiɰ	�1�M�\�ղt&�~;��t�e�@\"��ښ� Q�3\6�"���I�'��
.�I�0�#�"��_�|[`[�J�}13����ff�ճQ[K��_l(H�L��PW��r�:�#Ԥ(/X�Fu�����EPx2��4��p�I�(�U̞��*}N9R�h��M��Fǲ!:,9��c��.�!�Hn�ѽ?L4 ��d�y��sjy��*FѰ�e ^�k=¨����o�{�����a�[T5�_����>߯
�8��@nT$x���U�tM��7+s��y�_Ѷٶ٦f�(�g>���!�e��;��e��Z�j��:��]�V�$Z��a�jn��Ql������O"*ms���hlc�=����Yl?���1 '�*;��_t"P��X#���h�8ȴ�Q^��DK�zs�!巊�o4F_�Ծ�wH�~/t��Wt���<��bD���YfKc}�{����-5&
1��Rg�[���dc�#L��AQx�H&㝍4�Y�k��y���G���tyY�f�}���`��m��(Q�6\�A.��w��eN�&�<7�����`&*#!�-����ۧ�3����ޅ=�WԱ��C�),�o��Y.׈��+���)q�y�����^�n@��9�VI�T�ܿ��#�O*
DB2��UO���5%& ӂbg9
A\M�.+�_�y�T�Sca_���oh��r������y�"4i�,�b��f
���p����@�Z��<����=�ֽ`��+�\�1;�0/E����H��(q��h�`C�6&@7mn�x?�q��&1�A�s��Y����ӛ?~��?ث�q�����/�QY0�aɻG�� ��Ш©;�[.������D��S���q_�������G��V3;����{ۡ�-E�S��zN�~�*:g���K��s�_]���S43��K�R�H��zA�Ђ%�6��m켽i�:m�^ n���SanJ�;:��SYOc,����S��W�V�j|���Jʵ����V�O�5�S��v��)�D@	��(�kB��&���w��&&v��-�wF/w�Cvf`��o��<���B����n�/⺜}�8��&��g�s���s
��@D��£�e���9:�ҙ������|���S]�`��U�E�E!o�cx�Cz��ݜ�v�4�M4S;f�(+؅���W`��Q��FDr������u;���W�I��E��J6gHV��Ty�;~:+����e�I	�|��?Y���㘰e�,�9F�K��Տ?  �ERx�OUV�pRcqc�*�˦��Ԯ���ū?�c�����@j���������2��������WƎ����!�V������L�9���m��#`�d��dp,�@"��l�9�d���O�(��T��	KٗM��ǐ8�A+!���<8V=�t[	�r�E +�Z�\���n�GI�1��,S
�>e�d���T�i��Ea~��z�~���=���.�wbbh\2�ۼ|��.쉛����E�p��=�vkl�՚>�ڴ��G�<���*��� �G����-���q����D}��.�UG�"�9~i�I��TIb�
��IyH��xi"JPۿ�z�Nr���ܭ���(���e�R��|���A��}���_B��b�IͰ��kl%���[�8	#����rF0�"�9��������ii;��DF�m��D��]_�t�M����B/�IB���=�0�;�=�#��{���|��-�4�u	�˨�[�w%��8C�@� �t&��5B�
Ⱥ����m]!ɝ�V��3���QZ�r5'3^��t�R��zd�|��O>��1���������n����p~62	H�̼D�Ua��}��|,w�`��9	�a�E4�4��7V�{u��C����ac�M8I6�J�?"d�2�7��9��W$�k���#5��8�@f�.�_Cj]��:Z�J{�D$>2��,)������@BoR�\;��O� �a:��_�W%͘p�'ֺ
4r��Te�.y��<�@�% tL^y�v܉�
�?$��x���W����gfpϯP.V�Ђ57}6��z�Z���u(����>9G��>��eF�6���T�I���DkhL����~\ia?_0���P��&�T����_���>c��c��J��I�\5#p�j?6���$ʌ�H��L����'�Z�ft��)��o��i�%�"_6���?��o9�$�r�x�b8Ŗ�}A�p���\��-�Rh�	T���
ayY ,�I�U�/�L"8�����6�
� ��lH|�5	�*l!-+�qH��[�+N'h0b=���G��r��9G�+�wX<	�6%@Me�s����{b�ʷ�oU7�6��r4�gRgk��7��������u�a�e
ҿ�����>%�%�%�qܟ��ɕ��h ^ ����fWʗ�z�]�|ϬY���J�G�)U\�����۲��Eg ��t�|�dW�nA�f�Q%]���I�Ϸ�4��T�(qL��_��{�����F��5�f��~RX�e��F�?�Sò%k�i�/�$��u��D�*��$Ҙ_�bh�T�@�([/�f�<(�fjG��驷6 �'��5����ă�²��vD?@K���bj	j��(U3� C̪����|��(�e�.o/ķ۬�v�� �Au��/lA���>/��|�v�T�?s=���][�=%k�Qq N��9���kJy7� ��� 5��� Z�Xp~�r����_�
��u�i(_�=�Ch�c���%H��ڸ�$7J�k�`�c��|�ڹ�&pѭq4����@�Cf�@��2�K7�jd���ǈP�a�MUS��N��&]M]F��/B��x<�ٯo��rc�3����9ኈ߁w{����Qz]�����Fh�k6�}p�lV�~�w8^*"��#��.�]`���H��I�g\�[����_V�3�X�va�0�bwO?m��K�[/��]4���^K��UL/0S��v�\
Ł$�B�D,�6���W���F\�P��c��j>�31���H�ś�]�BP���o#O>iF�-�k��RG��&~7��G���$y
��;�8�x�3���ΐ̘ѺHg�26xc����|�9��&s��
��/�O�l'"ͭ�����`��t���f�F�4�tX��=����&N�<W8�`Y��l���#�i���e|-�5��H��j|��Z�kf����욋ru�����qƖ�z���}�s;�Q�(VC:���e� ь=$���I���dڭ�ݼ��$iW�Y���:��n%t���)���F��;_*����Ji^�Uq�i�}� ��	ߐj�棏�YVj� ��=�Q1�f*����'&�k��zxy�G��	&��\���w$�1s|Z�����A��S��`��V[�\��ےN	�� ��4$��\+~��G�/\��L�n���؟�ؠ��9�V
�j"�ל����*
�+%Kp��]�2/pg��23!u��]L�&�<��#��r�����2o�������;ػ� xv��ƌ�a�X}��#T�i��^#V������r\�C�y�{���מ8��lM<�V��KyK�P|�w�w;؍����?��c�O�-ݱJъ���]`*���
2��&��)7�H������d�腁%�~��� ��IY2vk$�����Z6�xCbH�Ó���,�r��{M/9�Q�0� ���{1� ����L�-�_o��b��\$��5�m�b������QX���U�x����~�]'U1{�sE��iE4_nh�C��WW�u� |r��y`Om�6m���>t>�H�\��/|���>��i�x�>�A���՞��Nn�=Ź���]�&�7<)����{LNPy�"�3�
��S��_�E@b0��rw�a����~�%����O��x�(��N͢r��b%�.�߾m��q0׈�ך���p�YP'�[c��,ܥ���\q��XZ���M\�������:C�s�9]���nW����X�r�|�*�<fl*.$*��`���`�:�4�o�|��y�\�ۯV,x��A!����<����ճހ�&Sv@�1�I���ڌ��E����cWϯ��V��(ح��h�@�
(�*D
��I��Q\`�B�2�����B�#�����A���]ij7� �{���<a�9�g8<B��3)w�^�~Ӗ��'�.'���P�+��2�4:fI17ZC�/����M��4���`�(��ē�<��N�#:�����!��9�S�<�o� 2���U�Uh�3��OrW�@?:�l���������&eq#��
v������W����ZP�l��Z��2������l������y����<�Ň����Z����fS��4������r��Fj<����D��'�&#�=��+��y�ܒ�� ԉ�:��1���n?�B��f�p1\D�^|���d~D��������9��9ޜI]���VT��}���wZ�� �G@����m����P<����˝��-8�T��S?7�K|&o�����1b��'��uF&.�W���ژ��C�)���SIb���K��T��p����R_[�\fn�\�c�V���/����K�M���\h���:O����� �.��Ѳ
g�%��SU����&��PcSC{�3� Ӌ+���'��r��Jp�@�,�6L���:$}��#D���V��=c�U�3ݑk��2�w��J�S0��P��M�ý&����:s�j�s����ϋ	�Q=�����5!��_WS�s��xһn�>v�x�%���+mm�k'���?�l~;W�ݑ-���}�����#KӝB�9��ᛊ��iO�c�24l�!L*�[j E�h�a)�f_ӫPm����'�{�8��H�ʘ�ZT�����X������?)�C�!�2��$S��Q�u����$��*�mȜ*q�5�K�$�"Mp9I��u��)���܇���|vT� �Q�>�ڂ	s �\s��_	1f�;E�a����a"j��_�E��=d�����@ws�f��	�Ι'�����M�][�n��L�Ͱ줈��T�L��E�5O��=47�y;cE@k���[m���F�Mw�-�������Բ����R�����s���}K� ���[��Ng���e�����u��E�yP1g�Sm��A&���fڽ�L�e ���*�����W� ��h�?�{�LW4�[b�r$E��=y*�a+D,�,���aR����Cb�j������K�\i��Y�~���FLIeQ�>O��a�� f����5��x&�*�n ����P9U�ܙ��ho4�[�7��;dKd|�`��QH/��r��<0vT��J-Є�D�oc�V������1D����b�kk��� �ф|?��.�`�=�+$���
� �L�x?��P+�2���n+~��=�B��Ol�����?!��N�
\$��W_�5#EC:^���� ��g�� �{���x�l�O�Q�5ʐG�u����BW��J�T���]D.�$�\�9#�B�L��W�bµƲɘ�凸u�)K����3�5_�/�Z%�w^��4P{�v��
�I�_�xk_j[�)HZ�B�4?cx@��u��퉗���$��
4���G�\g�@��-_�� �)OƍO���tQ!���;�������(Y� ²2b��_��g �2�%���f�*��6Y�Q����ӽ���no������a��mj	��S���>�?��GB&��P�i�YD�OU� ?h�|N��X�㌪�m�^������X$���D2V�߫S�����BvX�w�R��i����r�@^=����\�a���w�̀��l�r���4�{�ڭI�Y���@�� )��>1V2��=�N��@g� ��}`cd�+��������6_{�����J��O�C�����]q�Z,�<6Ll��@J����+Zz[�TB�~�.ZL�7��r��6�g~�b���q�Ͼ�5��ݴP�����JP<%L���9� =�
���Z�r%�EԄ@�k�D7�zlz�{u�	�� bxS�Bh�����+���- �x:"�a�！���m�'mQ���_�6�`�����/�� �7!��&"�h�o�(�/�����t9��ڝ�X�A&��>OWƏr���Iz��YCV����.K�󦎴أ����C��7fn^.rW�^���r�@��Z�^!!X�� b���"}Ak�=��K�[V�7L�����	�&���eo�i��-d�`�=W���2�Y�\q�j���r�[��O�Eb�̬ �:��qnA�b�zX�
ʂ@��n�R�v�_�V�<b�,j�认�.,W%;��)z���9�U��[}0JV�vLi�V���8�����c��k'�J}��/��CS�X��3e�nY���c.#mZ�m	g4lb�Y��)e�9#�}K�F�R�sՐt/c�;���;�۞�4?m�h��1ܣ�*��}�S>A|6����-=u�蔂�AVvk�x��J�K�Հ�i����۟�:�m��X���[p'HȞ�h��3�=��5�Cri��UC���{���z�^��A��/�p�#�fWC��@���5xFK���S;���B�[Ș���P=�D��-�ir���>"�t�֙�I{iyn��`RM$]�a��Anl��7��[S�ץq��+�Q��: ��L�ps���%���;v��8�
���ɠ:�v�!c*7��9�S=�##ޅɝ��x�Z��R�����0��QL�5�!�)B��
f��ς5R����4p�I6i�I��{�޴[K�F����X*���x�9��_��6[-���_�9�M�c6|��:��n�	��8�Y؄���OQ���[
�M����>ӽ�%t���I�}#@:��-��C"-�� �VE$����>�TqS�@�4�@hۏN+�#��i���c�;�L�Cw{�:chS�7a��8�~؍{C"��6�=��
�W�r^�O�\����N�1�q*��Ig<�}�i�>���V�� �tg/�5��Ѭ~s��2�c��k��b�����t3Vbݡ!�ip�w۲���$�\6����' ��S"�@���Y������p��v�c9'�� ?��9�c�����h[;�v��Sl3�9S\�\����3�{�����wv�J�|�ʡ�2�@�!���h�!("�:E�C�2�㮇�sS�Of=YV��`�&:T�MG���0;�~���VEc�?� 	Er���T��+�n�m1$�Lƥ6����|�6��"|�TG��~�d~ڷ$���łm���!V���#�2�ّQlg��6`$q-�C<6��,�oދ���шZo�4�	��$��ſ�U������)r�Iԋ�ĸ�m����F�VU��?��ܬ~)��2ҿ����}�����ӭt׶|�gI�i{g��,Ta�;�b��=�7?����	�Bc���k՗DAc��]k@t@��S\��a��֬ht�\9�����I�%Q}�`�C���T4
l}���d��Ȗ��^� ģ�m�I�$`[Φ�I;gW;<,Z�fk����K�Oy`k,��h2����'���Y@J\Jj}B��u`�x�F�sʖ`������͖�$�n�z��ͧܐ�LFR-�>XĽ�gNSŠ��זnAW��aU�-�(:%x�E�Y�����Dn�ʭN�;8!͆����1���د3��K{L_��Q��K ������z��7|z�<OSkU��b+�ǔW�n��2�j����|	�N�/�I�BJ�ߒ��ĥ�(-�d�=�Qs����|��/����a��U��ê`���nΤ�e%}�s\����L���W��O�f��D$6����?n]����x�?����d�}���i?#�:F�̮�n������Mm�W��k�[[�{�ZU��UP�OZ�ʑ��a&[h:%]���n�����F�A�<K��d����@�i|�Y
/��46'LC��+� ?� }rg����Hw7�e� �+'�1�P�5�#ͲxI���gy�3�����T�Jl����=,-|Ơ����Ȉ|w�٬�Lߙ�	$�@���4,��5}��'{�[��"-	W0�?{��U�9L���&�@��j�b�w�tS�Q�q%]��0��.�C���3������: ��:����T��v�ͥ�a̬����b'ԧ\�U�,+�Q�ݩ�؈D��\�Q��ɻ+0 ��7�B��L�E������Qz��g���[���WVn�*	�j��x�E��87����bbP���=h��&מ��T�c�ɱ':T�ѹ�����DV(^��rko�`�}S9:�qp��u�H��������X扨T�7�Y�w�N�	���/����PW�Ɨ+�e�^{�$㎖�kX
���?8p,uMG�)�.,|_C9~����l�F����?˭6�_��1�/��'l�^�y��;����<����_��G2�ag%1���O�:�1M�k|����&�1m�c�~jr�+����V��9G�M�ʲ������f���Zf1с���pc��8H��w�Ӫ�`�zޅW�a�H�d��D��pR�1!M$�;Yrk�O@-����W�J��1�<�.	���;<��U��o�'&[v�Y�8ʌ��F���]L��z?bKy:��k���]ס��8e��-S�H���B��/�k'4���]B6�R������6����_t��*�ed���D^�/��S�`�D�������)�w�[�A�^��F�tVL�8�e��Ôd����L�?�;rP�����I����x|�4R4�h�G&�H\��5�E-b�8���\�xlQ��Ğ����oP͚Wu�>�q����H�v
ӝ�oN}���^{�F`Y�6���q�~���ڻl�=�k��A¡f��Q�믆Ǔ��3v tY��� x�Z(Č����Y$~غ@��tJˆ����HO'������	B+�`Umr���9��Z/����^	T{����B�&�d3.��Y�NH E���NX]y��)?�!��=��zTC�� ���	���mS,��P���(�o��)�^��YL5Q������%ָK�u�:����S�G�rc�:>^�;%�,�������5�!�़-��=��/K�?቞L2WG����I-u��M�>�����"OF�9�r��"����������ڦtJ��wnj$�@"I>�>eg��p��B�ffa�&DC���;�Y�aD��Zá.1Q���s�?U�sZ�PL%�s�|lANR���\�s� ��3ґ�m�>���L���c{iI��j�g�g�F^�e�m�1V�[�7�/���M��E�+���P�\k�엄�YK�:4��N�}��1Łk���=���
N���!m,�r�s,s�v�T�z�Ԕ��^i�z�͌�wuk>L�|��d.��t��,����c��7GJ0t�jof<�,Y�2��g6k�ai��y�`[�I��:3�9������b�}�<%{&
X"2���sX��
&�^ ��Dh�yi5=!q8��^�5���o�rܽ�wd��^�Sh�Φ�Um��U�L�R��M��==x#D
 yF�;��c��T��m�r��R�F�좕��$i�u]��O�
�Y����%�'���mХK�eGH�E�=�)C��"򤢕�n<��Y���:��g�g�Ń���6"����!'�r�� �~��we����G��2�`���'���,�3�p�l{4� ���Iٓ\������Or��*�Ɗ���t�+"-j�����[��?i"��I'���k��@�� *��r��U����A*v"�.��!��t+.��-�	��}�+�d�e"C��0nR�ʒ&-+@J�;��
�7J=���ۏψSG~�d��tE����{B3��Ǔjs0���c+�u�Ϻ��U��ۿG<�N�����ea�֕�=�G/���lI\�m4�^�|R<sIqH�5
@�w`�U�����vU��\���}��%m9Xwp���"�CM���j�>W�e�����
��j��2Q��%i�tV��X
1�?'K�Q�`.�۔ҏ�a��yx�M�R�^�\�c�t$�B�`V��Y����?���l8ç���MF,���������r#?7�~�IWd'g/o�	�RFۂFXU^03�����!�
���9����\�^ C�Bc�a�j�՗Aӱt��%��OK�s�1��8g��/ qa�v��;��>ai���m�Kg��f����<�Ki���1��u�:�\�;�}�:|�P�j^�D&�e��{�1��j���i_�V�gm>P��̨���~�M{Qc/���L�)2�h$Q9���4�'�=)ON*RB-�����	P�MN������djo�ҵ�>}jm�n������vNH��#�_�Kq$��F�wx#�v^N��C ��,�6NaGM���X�|m'{�s���f
�ь��)�0���(�+��uq7LM�&É�BV{��Բ�����g�YJ6��f���Yf���.>Ta��P����B��gb����T�4MRF�3U�́�D��l��U�^�[��P�J�>���^�p,��"�٠Ϊ�:�]fg�F ����ދ�?�Ѧl�?�y���]�ې���D��tR�T��O�?$t����=�n�z�E������U���9��j������v��밚�ky�d�J��Q��=�y�Ǚ�\�/5�dot��(�-O�T)���%y�����
���P ��;OKc G���Vd����Y��仸,, �=�}y5�2�G�@�盁f�~�v���߲��@.`�?m.D]�PF��N��K�M��7�n<�1�rB��/�v�\0��,VVk=�s�\�[G9�K�%��Kw��S��a�TΓ�y�7{��*Ƀ��f] ��$��Ǹ�r�3Lb�k����6�XW����3`��������$_q�^[&x
�b�1)�րѲĠ�L�Oi2�<fǑ�c.\"��?�d�?�윻�cǇ*i돔�T�������v��/�Y:OD�� ����<-	��g�̱�j���b7H�z`�4e]c��[���?�x\������.*����ϛH�5fvMP��ytwl1��"
�z�������@���M�_=���"`p�i�WK�wK#�՝��s+((��u�<�V�B����~�їy��Q�5ϝ��8�IN"^N������u}�[则?�[7Kv��Me�<����[��a��(��{�R�`&�a N��k>�����-���/]G�w�E��g�'�֕�[�mIV�<�+Yg�!�N[l(��hE�'Jo�7�@�5e�H�j�v�c��l✡�ou�Q�<{ث��H����.(J9!��>G�Wdg�����p`s
��r#F"\d�5`h�|�cd\�l�L�ؘ�()��kv(��W��QP�g���+�{r.��!���R���e�*�e1��Ht�?��.=��X0cV�X���S�o�򑹛t�+s�������]S����˥Y|)_l8��1�^Sw���T��M&��b%^U4�\��=U&�|���ij5��:��M�M�{�;Gr�g�D �Ȯ}���vY���T�x 'f�����yz����c'��hV��Ҧ�Ɛv�c2�9q��@��ܵe=�y���M,<�7i�s�24���b�hR��At�45�Ӧ����o5z=G���ʳۊcT�	J�DJP+c��r�~BQ����3XN,¸��$~���G����d!=f�i,y��k�#Z�IȺ�0��"��A�ER]*��"Ϣ��G��Q�.�����X��^^{�fs/����0��זX"�ׯ��.ZH��D�
ykt�~����A��Q�7V���.��%W���T�AF�"T;���eM�����Z_˒��H.昀�~ݨ�8I�� �#{�N������I�a�Ad���
V�6ޘ7(@�nZ䌆PY���D�� �;t͡����4r
��<"ɞ�4��`,�􉞼��y܃�L�l��'������~��vqjѧԎN�F9���h���0Դ2�v�d�C�4Z�S+�zͷbm�f��d�9��E���L�e�a���$�%��%Yx�W�
�\���&9�f��6�J�;���YN%�a�3���ó�����G�rHz�������e��G�R���̂6,f��z���(�Yt*֊%�drwT��H2?��蹑�K�� vX?��1�@�I}�P�:Z��.�£;_����b�.0����}OR��r�*��dJ��/�,!F�FR��]'I��;��(�l�rį�m&D���4�>Ǖ�s�G��]+�����h�%�J�1QW����܃˹��Eۘj�у���݄;��8�ʎ{�����~���(�q�-?���9O�,��<}A'ZW�b�z�U����O�*�v
��z�t_�������R�r�B�As��q�B-qlPU��!�@D�(�>�����wT޵���XNj����$�d&%L��P�
L�'�yv_��$O��J�|�uNf�Cp�*��9\��ϳ��MG�8i�]�/fW+O����k����(O�pjj�hJ*��� X�GG[{�7�Ѫ�M�5p��������_Bo�仜�.��z��6b�;a{�W5#���-�ĕ��a8�{�e�?Ug��ֿ������0��b�9jJw���-�`�P~oo�����k��57�{�g2h���p.�	�!0n���(�(i����g\noޖ���|�Ś����?���ĠU�&D�`T~{z�C;&K����iAf��p�s���r�eP�^55�ôGBB���<��PPv5�yPN���Fʞ��x��ߜV�����|��o�ԓ���-xQk�� �S�f�s�!:/��E�q�������SEs*�fZ�I4",�=����#<M4g�0
m�[u�Ir@��ws�q�B��r�d�g�ˏ%�z.�\4���w(���Hp�nY���[?P)��O�H,{��9�WhS�;8)�\�n�6�|8��X��t{�~��!3E4��w�n���uV\h�a���A�L�˕"���[��A3;mխ�l�};2$Y����y]�xad��-���ke��WW��W�2�Vr|~VG�'<"̉�T`�����U5^;�m�']���&��֘�VqC����e������_�s1`��	������W��G�"jL������g�G^MY��1�LU��,g�1���*���suj��2p#e��� �7�0��9*���:A�H�~��TL�C�ŝ��W�xʜ)�rZZ�
�jݷ��CǕ^��`iȢ/��q�z�ϖ�t�`1�?ŷ����Ѷ}�\��(E.<�Ѭm���1�OI�&�e��f*����YM��0<h�{�MM���ֵsJp!����mK���D���P���PHN[���W߮��B�o3�X�Vh�'�� ��Թ���Hq����?`Α*:�r�}��LPnS�*���������\�G��sg�7��>�D��6�.�*CU��²H��v����?���+5k��q�n����U5�P��	����:q��4����#��3��I1ٙ�Fp�y�v�����Κm�6skW%c�W�����踠 ^�;��k��S<$̦��+�9X��Lm1��C�F�ǚ{�7*)ű���;��{�3&�`$��!��箣�FV��I0�;�V��mŘ�O�����⸆;���/��4�g:��)"'����
F��P_䒅7D����ڋg-�!��q�K(��Xu��Xg��/~�L)��@�,�����k��-��?����rGDE�( *����M� �3���&�n�!T�3O�Mt��u�i�u���GZ-����`֠���r�p�o���z�(�N�OJ�\�	:2�V�a�8,��ސaF<6ןl�r��~~eܦ�i]��Yhݺ��ߗ���;��c���=��vײc���w���͂*!���0lm��%���z7r�vM/�ֻ�Z�=�ǃw*2�O�7�y�0S����6�R#�cÙA�	�;*"�3�'��Hp��wY
ur�{���� ����>���q���m�Կ�(�Hy��[�z��c�3Լ�� ��c֌e^W�B�+�h �>�"���m��wǊ�&�b8^|�IY�~O��r�L�0瑪b	��b�S.�}(��u����J\R�&�/�N��_�Χ�˞?�HT��:��%p����B���@η����J����Њ�r�ry�j���n�l%)�(�Ҫ���r��qc�NO^s[���K]�檭 ��h,FQ~��p��ezPs����G��t�g�c,pN�W8kc��u>�Rlg���3�Ci�~(���K��Eh+�b�I�4�o�"\k���
W7�U(_s}�bČ�� ����ve��=ɑ5o}q�9�YÅ/���G���^=��� �n�~f�~L��'���ym>�@�_��$��F���T!�}]�cS�'C�FیyX?Z����������6����8�(�<3X�Y�	��)�,��1�j̔�e*�?�bq�qe��g�"$�(N`]ͮ'���nxr�~O@�g��d�Jrƚ��h��T�$|^6�QW���=�U�6\�GB1���� �Zlv�)\����7m/��2�9�t>7~��^�d�i|#eI	�?�Z/�Ch�#<���
�>��kS�&|&�u�Vw��k�}r���s�x����+�s�=I�O���~z4ò~�~�.�zZMT�u?���,���{&fD���;�~G;�H҇49��p�:b12N���N~l�3O<}� ��NU�5��G�։w���,i����4��$lB�8)`�T�E�2H&�b	8�SZr�Oɷ%��*�xF��8H�U�|�n�u-��y��1���U�N�ϹJE������8A�YV�~�YiF�J^d�h�0t-(�1�8m��/��0�:2j�.&ӟݴ��X����8.��dH���4��g�1��=�#ݾ��/�˰p�[G������qE�!�"�Ci����~M���<L u��ox���=���_�VW�;�����7��~L��W�g=s]F��b��#�3S��g���j�|'�@m�J�Q�i4cS���e�G]�&YH����ҏ��N�s���=*�on4X.o��aU�V��z(8<���d1�!�F�qe�y �[�(�?b�ndmC�����s�q �� �٫�(�m��{����%ȇwe/�i�$��I@�˕�K�Pz`*�Y�5rQN"A5)��7��/���:���28ڞ�C��Ry<�8���L��#�$��W	ğ�#ߵ P��Ky�3�~�V���$��-��1��q]2JK�f1�3��7�J�_��J&���a���D��S�Ӷpr��k�&b<��O����M��ԍ	��S$����j�L:>MQ"��vYS��93ԡG<A!���ZM���:M����toℒ������s}� �pX����L^�[ѷk���%�%�G��k��w�����!�~����⁅%�����I��h�כ�9��2c��A����%��ozrӺ�\t�:�qK���fO藱�yI��H��T�
��yvb��:[�����uE�ǡ��,H��C�Y{���i��ޘ�Bh;�«F�b���;��}P`
Ԕ��Y��^>&k��t��\� >�<׻��<H���.}[��3�����_�W�� -T�Cc$���[��&�9@Jm	~��q�H��m^=�D��.�Cʥ�)�gj]���K���u�0�PT.������x���H�]��ѫ�)U��W%���:hY"���G
+��[��e%g��{	$�sj��� ��u����ו*:�Z2w��>*OWΣ֏���s�uڊfR����4�/������]���� d��S��_>�6���˫��F��f�?ma���t,y{��礃�Y��3�0��xobH�[W�r�3b��e��-Wp�My��>���$�&!�I	X�E�X|���9y0�Rp4���A���MK�v?��	�D�|m��
�؅�Bq\�t�	~�g������H(��{Kͥ�Q�8��������@���ߦ�0�"��0���'����{�5!�j�a�Q��������Ž��D��h���Yo�P��MR�Ik��g�g�i��%A�0���<�|�VW�,��Yɘ1�w<�{�
قQ���68��0����S�'�Լ@8�ey�����ްb|Û���!�sW���[�T��4(X���K�ؑ?�~8p4�)�|�R�e�`�/�d�ľ�0|��nr�u�]�WnȸR��2n��iCD��3��eF˂�X#�R�2�V��ǫk��u�dh*���1���v:,�1�~ť��z��]'Š��b`��S�:^mGY����"�irZw�K���������@���u?����Zب�z˧�����y�MsuV���o�-L��}�|*B#1�EG`#N�:���y�uu�Y՞DH;Y��+�7	��c-z�3�ي� j_��;���1�=��ś`�8k��T^�Q�B�F���'+g���X��v�Z����M]����(nX���n�=�,���r ��0���
�P�����v�Y����#A���5���b�c������<T]�
�M���ԗX��Ǜ��r
���_�	�ֱq�]|M���ɐ@���JNM�C�;wp]�>�;����FM�u�p�P/�7H��6i6~�+^���|6�08�9�{-T�ZI#�"��=Ю�#R�,aƦ^�sZP[Z/��&�׺�����D�
�)'���ڮ)���>C��!�3�d��Opڈ*��Zl��jz�u+��7����iJj��H��jX�I3�+�Zmk�?�B|b8Nwq~����=Gm8�����G�̈n�#ޙ�ʃ�洶��+�襲�&eE�(/b�͕��c�	'�K��b��2��_$�}��Hlص��`)��t�t#s4U����&�8R5���g1���Z�����2oS�k��M�|�� �e�E���N�a�'���lm�L���E,�{��ӧ�[��c��N���v�^��������}���:�β��͹Y�!�M��zD��t�]�උs��IN�����^�Ü��N����f�ɵ5�%K?��������5��"p�dP��YW�%��	ȳx׮Q���r{�sG8<%���2��G=7�.���f��?b��mI�c��}�/8�f�FD�6�����ڽѵ59���Қ������G�B��ޚ��'��t]]W�;�w��M�3�S��j�&tO�^��UT���,#M$��g;���Q{w�i��Ԫx@&�{
����Qn<?q�Y�h�ܼ*� (.jq��6_�mP�8�bh|X�����!�ܕ�w��pa̬
�] �K�P1Us���V1��.��08�\PT0��;U�2��uJ���9��(ۘ��	 �B��f�5eB������(�8���͵a�Y�[@c��"}|���l&��δ�N튦gG��'۟� ūKTͽRY�u�ps�<@9B�A\��S�*�FXb���%A����˃F�D�#g:>����֞�9���X�Qg��ɸ�@9U�E'ړ�dֿ1;2�n���@S���j���s�?�����-���7E>� a<Q)cˬ	�f�w׹�x$����ǫ�2U��D@z%`#�3Ǡ'����]P~tڦnjlˉk����`ۚk�C+@�:�o�K���$�_}! � �'�^-�\�ÕW��s���39�]�p��m��z5P�Ӡ�3g�޶M��@"�o{X\@�C�8�s!�A�:��,A�e�.�����O@	��ݒ	�96�X��z����I�{�����	��V�nS?z��&��ҍd�C��╊"knN�}AkK'M`�r���綐���9�;�hν�,�ӿ�ҒP���uZ���V=3�e������){��V�XR��JF�����3d�bog����r6��M+��<���S�8|���/��q�!�S��?P�`�0��y���Q�b��4~G&m� nϷ�7���WD ��*U�e��%\�5#]�%Tx�����_����3����{���@����`���v�C�|5���#�!��~@�|-�-z���pJ�Ҭw}�o��2�ɾ�z!K��i&G��}�}�S,j�TF�KH��#0��~<�HL#��1�P���"���č�@�tN��b��蝞�����0cb�tDg�&�۾�u������p��|��
&EP�:)z�c������ER6��{G��v���0ˊ/!�)�C��%�X5�]��/��G-�3zm�1#�s��@�%��sC'�x��V���.�����C��5�5<f�J{���CLn�D��4ٱ��NU,�a����p.��j��%%�Me9���
O���7P�h�QE�׀�RV��
�ۀ4z�xg����xI?2{JK�B*-ry��:y���@qBא�S�%�*#�������^����k�Z1|�%\����?FJ�nД����C1"�C��)ٟ.��8q��ClqF���c�f�����1�3��	�FIB'ѹ�{=PT�]	(�S�GV[Y��Ԫ�d)<�긽�b��H���նA�7K�p1*����R��t�Ͳ����뇫������RKㆼ�����J#��_��o�o뺗���B�������=];���LI,Sqݓ���c�q�ҥ�}z��!\%߉�w7�ϕط�	��]x_�wih]�77r�SwD�	 ����鷗�	r�T�[I_3I}�GS�_��H���l	H	�cZT�t)�K�-"܇���Q.�(�DP8ߋ � �WA���G�e�Ơ�j���H�ݯ��3Eɥ]+u`K�=��p�����}��e:�\P<�<^�N�)%����q[��!7��>@��Cx5�Ź7��*�D0st,�ew���t*��7�ö�P�#��x01=�N�����4|�H+&R�	k.&"ȨrLK����F�����Â���o\��sͶ;��'����̒�ĸܘְ���}�-�4JL6آH�lV�	�#�����J[Xv
u.Hg�\H~�{R�ב�%@�Y���~�����w�`Vru�'"�x��- �J���?ı:ƛ��G�=&���m�С������s42Y*�C�N��5�!w�����Q=��:Z�צ�٤O��?�����.YS�yD�b<4�T,�gC�cz?�i�����_)�_���)�1�bqI*���c����<�~|�T~��Xd^Il�������+m�S���h���'���n�E�U/��i�Z���J|����g��	�m��=��M�ِ�Zh���V>�7H��g�l��� IQmÅ�Q��n�Gq�9�L���<x^���?a3RcY��t�Z&H�A�G>�H �2��e�#�gpٗ�F��йhE�s� �:K���D��:�B\�o5�Z_p�"9�d_��É,�C�L��L���"{�xx���!-�k�A|<O�ХE� [��]�� T.塚��.��7�5ѱ���Ro�s�'���d�>�B
JɘO؅�)A���΄�g��g}���T8.�F��\*����ӱ���*:n�=�pm&����n�.%��Z2��{�B o���,�)ۯF� �U�P���RE�n�(���߾k���G�KtS7"���BT_sHTn�¶_%���+�䀈�S�q�q�����<M	j�c/��`81T(�G�Ce1�C	���"��� �S�_e�s۶�] �r8¼Q�Cr&|�|,<�<>�b��'����}�V3��st?�`���(V��9���]��<�fS�k����ĊU:�H�&�o���cCjLV�R��R�p�f#�]:`bcZ� �^�:�r�/BUӾ���k������Y����i� 6<�q��7��xnc����;o��UD/H �g&G�{��&�u��mY������ɪ6vU�P?0���r�/%٤��,9�(h�e�'S�|��t�MZ�G:E<�x�t�Y��{Xi�� �H�n���(��a�LV(=���� ��t�u�r�(��$T����(�ہ��$���6��yJXZR#Q��9*qa5JZ@�[�ϣ��KSs J�\xa�8�[z�x��h���y�"?�\D�Kzm������"���r�-O�B,\z���7!Q��_Vv�^FތV�]���$�a!�?xVL�����`���Vх�B��t(u�a�~{<+�h�-O����t��4g��uk�O0��#WY���p���h �5_�(t������w	�Oߗ�5���W��+�����Hv݁�SZ_�;H��k%��Ui��v�����7`x7aͤE�Ο~�	_.<��`�a#���3b��)�x읽j����2��<)n�xq'���9�DóU�m����7�O����"���so�^ڼ��c����X"|:�HN�B���#|�N�9?ƀ��j=�5D��$�����"H�]��Wֺ���]桂h<�R)Z�VWMT�q��� �{����V톥��
�<����&�)�n��������s ������9�W�E�g�D���O-Ḵ6uxՋ ���t���#op���>2�n��^[��xHD���s eE�p���1�]��Fj,Nl�a�����,����ze
�ˠ4��1��!�4�@�	��A͕)z w�e�7I��Q�3f��C>��ɢ{�?��x7�%�i%D�]�9�Gc#`����n��������3�v��h�o5F�l~����~��F \C��>W���e��u�^��lYq�2��Hh�󩿙��Y�H$�B�u�s0��}��
�-�l�碯�n�l��y�9lI��	�&�+\߾��P3�X��0�6P��g��x���bZ��yB�<�*�f� �m�k�:߭p�Ы}���T��Dj�0rQw]j�_@�].�'������3�P4;��ä�n]xeB�8���u��s��@����;x��?HC�#-����!iV52�{��<x 1i���G��qM6�+Tg-+
��@?DƲk���{���(��u.v�**��l�8�ݻ|�N �r~;���|uϱ6�����S�چ91&��2DUҼ_p�&D�mH�(f�Sg��v�9~��|�˙ꄨ107'�o+��,��2��fTS���tfS���/��9�txQ�J�/2:���_��h8��O����k�l��-��ԑڝ����9(Msy�!!ˠ��j9��7�����%�T�+x�zco&��i��/Vo��0�JM�U5a"fx+`���B���)Z~I�,��籦��KY}�ភ����~�&�r3�=b���(�~��V�v��K)�μ� ^\OT��?V�07��u|@�"S�o^����
�������t��n�qS���4�l����'���K���/J��W���״��	�� 6��Ki�*O�n����
0LRv��iu����>�`zZV�����g׍��ʴ1��P�8���hyK���{�ҦP!�x�or���'eHؐs��J~З�7#�v�_�o�(�9��	��4<��e} ����u�����k��ɛ�����$�BS��?E�	�7-��e�,��ӻ"M�珐��9����ɜ⪍��A;|�$Op�VB2 6�8)� �5c�8�ne�o�v�5��ԂqU=z�}яU���tm$*��?Q)�Y]fO%
<�0y��`(���ms�"��_�$��n�F�Ns-z��X���YTW%w��+�H����G�l�yڨ��[�e,y�f)��h���Ε����Qaڶ2%Ƙ2tT�ɜ� ���\)�^p�Wp��~vd����ZΩ,�'����ܮ��xfޙ]�j����.6��_��e
ظM����	SX�G��F�sF����n}��ߗ.MH�Yq]�p����Q^:�X�)̘
ۜ�;I%r�G���9z?@�:��T�a"��TZ�?�!lI]��;��X�Fǟ��/����d�(�n�侈 ;��ZgO����1.��������P��$�{�r��P�q6��7T'�y�4" ��pmO�q��z2+J���LуTP�U��$���B�+-d�y��~B
�o8�,A �65��þ��%0��T��)��! >��q�ZC1�k�i�|����uv�|��������0i�CjR��ԗN��a���ը�ă���KՈ�'�^�Jx�j���'��/ZX�����4!�SZ�^GQ6��}�ؘ��eZRP�4���dh�5
L!�(�P���`�ivd�VF����R[6��B�J:F��L�6�5�l�
D��v�(�{��a�O	$�4���7M�h��q [��P�y|8
��>_�\�FB[�ձ"ǻ���!�s��,��EU�T�`��)��doJ^Ӆ�r�p�����8��m;T��>��N�+�T���,�0���:���]PW0�pM{��mmu>���*Z���1n�4�粿���)��5���@u3���T����qw���S�lZzqkq`H`�U�7	��0�Te��x?� a�w��(�ɩe~32@��t*�}��˘w.�-Oè����'��Zl�?nt���@���Uf���̭op�l��A)�:�$�zr���7�sv�r0�C��y�}%$�1{X�o�8ѯ.BJC���N�xߎ�7���,�8D��u��E��>C����u���X�cT����b7{6ksk�L��ƺQ�QOrL���������p=g��Tp�
G�v'�Q���$��h.zM�%F�n|�1���_	&xz�p�z��8y�_ŵ}e咚o�a|Z2��ԑ��mm����ki��`�u6#^��M��4K#u��@����l�G��l{��<���I/h v�������(����f�S�nWs�z���)���>���)�'�� D����ȗX��:v=���I%!r.�D/tm��a6��&��u�ѻ;t�i����M�nۺg�%� L࢚�yz*af
0�2�g:��
;�=c�0���4r�%Z�J��MN痦Ny�<^�R���k��<&���6�^;D���=Q�j�2�I0�N��f!��ye��c�sx��P!2�]x������4 3�W�h�c�
��B�1In(4j}�������K����+�x3����,k��ۉ�.Mhx���t�� ����_wL]�~}��6$���d�8m���&�Ѹji�ީ~�r�z��B�V�7ϛp�V�u&W�i
NH�P��j��&�1AW(�l��}���5@����u�,�U�P��A{u3`��jyI��1�����:��ָ�o }~ H���~X&���h"-4�>Cު�a*H�;�G'��P�J8�1�c����zp���&T���4\�������穄lPEY��$�ph����r�W�.�ֽ��3h��qH�:�?]D �0#�s"sY3�?A5�h�\e�!�.A��Tq!�Ta�eXґC�*����A���(3"��Q�d�xZx�e��̔�Q�������T���:��rb���m�����R
'ȃ5�� KA�����/	�,��4o�i��h�۹|,��&�T�LB\�d ���d:C!���bȩ��h�j��Z\�$�!�Y�dAɆ6����m,
�&�7�#?���VԳf1c��$�����Q�nS��1砫��;�# f�`X,�8_�~��[��ş��g".���;0��+�2��E�v�4n ��'ݗ�j��^ {꿛�h<�p�[�ʠ>�:��e���A��� ���Z<30M�k���]%�\Q��}�����7�� T�]�Р}�������q�!�y��}��1��/0�����i-:�ծ]�#���l�ԎqQ�mj�~��������L��G5aT%�;��r��~JԶ\���9xt����@*�D�w[�4{|eT���O⫢5wu�U�z=9|#4����]n��m��C��3l�f%�f�, �^�9Ҥ����؉�e �.�8�HG};�Κ����&O�EW�}	?j��q+A��q��ڵ��"F��ū}��\��~T�1Qi:��������zībW��O�g�ٕ�=��%�qD o��rG9Ɗ�C��x�m!�kB��ğA��Fm��fAP;�I�v́��~7��ۗ�-�6Q�E9?�b�%e��|�"���Ъ���
oA��mn4Lc.y(�0�V)|wqC��;E�N���;�7�[� `�!�������쪘Q�ʡ�d|L���9�΂)�J���h�bj��!0X�\�������xa��GBJ��bFǇ��K��,:|�a��߿��,Fn�I�7�G�~��HmZ����uW�m�A�x��"M��B��|��1��5���Qx1�Q3�=��ݛB˃���M�^-3-ۋy#�����v������E,�d Y��"R
��+��JBt���(�C�9V[)z�ϱ��VkUB5�傅x3��32���E;�r�k!2��jy��7�3��W��7��O��U%�,�RSGd3��3���Z:�-)�;���2���Q�e�4��9��,k1�O�42?E��|c��l��!rH�?��	�=}��s~�	
�>V5�h^ᑽ������P5
���<�.ՙ�65os�b�@�ݢ^U��m���n�'����q����2����B9����^ f��t�w�����ح����Wn�9:��x&i��.�|h3�:W�=���%=��~�:�/�)�m��̂<��
��s���4\t-��3�kY)�2����A�3��#���1%�@\#�@��B}3���D�b/�Zȶf�o��!`��"PB�?e���;rh]�9�� ��㬓v0�E��ӽTG����ji_��n�U��b��RY{B���(���F�Ô����?d�w�LJh K B�a�z��b$��`&҂LG�b���]uђ.
=�<M�S.�WĿ�
�������x�<g'�t��Gn�S$EZ�~r�2�y�Gŗ���ԧ��a���u�	�$b�g��rP����>.c��ő�1`x_���U����\�O��-��{	�fSE�Z�㉈�'_�q���|W������Ue�/@&��{o�#p�ݯ����Tg�b����A�'L�K�nP,�g`>,ϓkc�����Z`�'܇�xd��	͸iG�/�.�|b�t��E��9������0j5���\��07i=i����E�3C�M=�^�kĥ����D%aၮ�
��,W��F�ڹ\���늋Z׹E��@;�h��C�AA��	�bC
��a��p���$� ��Y�-��ސ����j�W@4qmP̔5o�H �j�}P��_<q|���Ƭ�!^��9�q�t�.j#E�W��2G�\ɾ�q(�z{�C_)GM�ew�l
9�c6W�:O}@�er늭��USU�ø������gЗ���/����pG
�����3���4'
�����F��q�"�.���T�D�Z��<t#$�������/����c���H���辆����B��i��Y�l�S�n�>����
𴙜=�.,<Шe��+O=.~
]9��>c5�M���D�0�k�y��y%N�_��o'�'ՙ�6�X�~4�m�+>#���i��F�|�G��j1�jNG�Y�%�<.�ta/��mw���#rYU3��e��ß�N �p�L�����;G��Fa�� �~ߩ�^ƴ}��<aϦ��o2 c~�f�D�E����?��St�i���d�zz]�(+r��Z�����;�Z��W��뻑��� ���-)����UႧ�DDi��c8Q+B�[��]�Q���w4ҳ�����h{H%��y]n���������@t��J��+���*8ldꕩ��_篣��e=ᄸ]�M�bW�|k�H�x�aY����?+���V��h�տ.8l�b�gfA��"���M���>d�8���Ɩṟ̌3�ӊ��j���+��u��cM~X�vc�)��>S��,���'I��LB�<Kܵ͏<�54�h����d|g����������l �q1�� 뷼�r���Ē0��^Fg����C8����3EYL��z(��������4��E�	��9����������w�� ���v��A�D?J���&w�y�d�z˵ *�<�8�����}��,,��^���{�67���b�&ݿ�Q �Vh�̕p��x�;��J%s�����ܼ�� W�oiKA��*u}��U��g��g�o�l����Q�o�x�~e�i�^���,�pQ]��K��P%@FG{dszN/a�2%��F��_�X�(�c�8�Ua�ڐ�^£�Z���tع�mM� ��kۑw�ǟ�'z�L�{��� �+�QlWD������1�&b�G�k�Y̹���,s�� �U��K.����&>Pon~}�vSZ������􋮡/�~L���]��1����zx�w5���M2�K�h�o����1��CP���7����<-�u���[�07��[� ��LrQ�=����.rsQ��s~�1�B��Rڑ{����U���rV�^� �����3����R(�wZ�G��b�n�!I,�յl$ ���1%�d��V���k~�&ަt���V#�!g7�ؕ��?�3�'�P�Y�}
�5�H�B� ���t#�3ѱ�)8K�)����A����KTO�
3�@�= ��q��捲�>�����Ö�T����,R����B�F��d[���%۟�����T���l�O	�$FhM���f�x�):�8�H��~Y�&�+�y.UPs�oK� �~Xj��F7�۩U��1���ھgB��{*��6ُ~HS�"1�6 C�R��oG�S����Nbn�����ǚ��mq:2��9$1RL�s4g`gmPF�&��6�[k�JLb�����Dt�N�(�t�/Z��;��ص
�h&+/ﰸ��`.M.I�_0Ph�{,T���cp��yM]jT1�KH��q��,�����B��j�
4��t/e(B��V�wL�������|�2������T��!@��9�p��x��qo�9���p�3��3�p��"�C�B�8�
Q\���D�t��hȎk�e��Ư�#�B� ͜rݝ�!�W��r�V�`*�P�VQ.v
�䀿Bfީי)u������kh�]����#��rb��I[T"m�t����M�>$+�|f�D�-��j��Y�����}���AY�)��Ѷ���$n�R�lOa���p�C��E�ؠ�qKj��FӖONf�S-J�W�YVt��f!j��F��VM�C`�����2�V!;~���U��O�9Lz��nڛ���P��V�ĸ����O���;:�@�T�C�M���J�3�Ł�V���z�4��S^T*A�Z����߯I��a��'?D�R+F�T޴��cz�9c��%HN{�*�z��d�OΔ�x�&��b"xv��
d4+$��8A=F�,t���I���ЍD���Ǚpև��J;0S�O���z��A�Li�8TM�d�p��]hW�و�fe}�a/~N��R�+��q���Y�MV}te�eB/�* ��6I׀Πl8�>㟵I��0C�X�)��KɛH�&�������j%�)����~��W�p�$�4���OB���bA�=���pmH,,K�a�[���.X��F�}\u����0�.q`�ޤ<�$�GC���N H����TJ�;��ht�VE�;ۄX� � Ce`��@Uј[+�P�k2/B�˞@V�	?���%K޼�i��=��k�ȃ| ��{-|��<YϏ3Ձ�8@.��]G\SZ�N��>�XA�D�4��3�Z��� ��`�6"��r'��b4�ʹ�4u�I�|B�YQ(J�܁;$ˏ���c�|�˖)�K��0��8u=�:G�fk/�Uy!`��y�����w\�С2���&1�Br��+���������E�$�8���-��좠��bų���'x�{�;[��T�IZ�T/�����k��@�l�ڍ�^���Ps�;)��箙p���k5�n�]�?��ɍa]{�A�Ũ����H�a�G�!YI��V�����jS � ~j|�Byy�{K�Z�םsJfKvo�2�Z����3����||O��l��J��6��0݆��z�������Լ���*i3�e8%�q�Gg��^ˡGkd��/t��^���!�~�"���Pj�	l�����J4ψJ�tgH�Ͷ�����  |6�M�s+�e��n�6P".�[N���!�mܨ}�_�.�+��Y߾�CC;��d�'M���=����&"ob�ʠ4+4+;Ϯ!� �/�(6�J�-�H��-<�nɳ1���tz��>��軑e�(x��H�|�HISv�/��N�Ć|"bsD���I��5��T]S��j�2�c�j�r�Ø'%�^�����Z.t}C�-x}r�(�J̣�%ح���B|	���˖й�PvsĲ��^lT<���o2r�,�R_�;�e���g���p�R!tV���`~���X�@�pN���q�
C�U�aTZQ���0��*��S�&k`n2K�p�����d*�E�����^n,V6�Ƞvb�ͼ:�z�`)e�UJ�a~@Z˄�I����L&��&눈sZ����L��q�?dJ. �@-2@Q�yL�_N�#��)�}�**��3x����<VÙi�� U�Z ��4�Xf�ZE ���H%sV��:��sxcnwl�������x`�H�g,g����8q�D�;���P��iU�ј�M�,I�V��暅*t~u�WD=20y�{�Lp)
�.����޺޲�����V�þ�R9)BR�M���b��ͣ�"nKϴ4�EV�@}}���tQƑ�H�U/���ަΨ�q�p��8]9B��;a�>_�����l[I�ѩn�JLK���:%6'|�<q.��1�H�0p���`X^�]Ӹ�=g%�H���p�nj���1� �2�����tqQ�_ ��- �>�Ә�_Q W�f�wA@j\+5&ہx'�X�~��o��W;GZX�ʖf�����/� �4������n6�>�^�<�k_�QN����+�kX��@��X�����&9�K��P^��TC��g��2�P4�r'����Z9�;�z������VJ#��S1�I�D����'�\��fgt�`~7H��/�����'Q�{K���==����NO^�G��4yT0&�I��]F�ӽ+� %OQEuO�r�ZkcY�XJ��-e�ʙ�4�J�C>G�Q����4�6F���"�
���}�]m��� UY�5/�𱌀�B}8A���t�s�0�]�df��ʜ�g9V�#��L�2�;�k��6^c  ��(����#�:iNX���φHM�e���
%�H��e6�g|���9�<w�f.S{Ѩj�8jф�ø�/�2<���e�Y�c5V���O�����Nm#��@�)��� o~�0�W�0c�؞3�^;s�����E�7�e�CL�ڊl��OM<��=��� 2S��G6�\N`���Ob3��;��F�9�2�t*C[�ڦ�FFf<W	���!9Yjc�$�"���.4�Eg,��p%�š��%�-�n���%w�
��o�Mh>艅�afʶ$���,k��[�Ӕ�� ִ<�u)b��wt�%�Kk#xo�O�!�X`���Z~�X�1���j�V��۟T5�d4r5p�����q�;˕�:����sX�eƯ1���W�ɞ4߂��v=�S0x�(�3����y>���F�9�z���Ӈ֩�g[(	��#P��^[l�����Rf�dK���c��GB�3��Oˁ�>��o=�.��g�N���2&j�-����= �`Ed6X�Wʯ�����z�U��"�o?%���]oF���jef�gN�b��s`����.���b�� ٞ���|��GC���=9_��)Ŕ;uZ׺�B�b2=g�8����f�Ь�	��#LP���Y�
����U�}���˜4�����	3Tw%��p�Ejs��#$�Km�P6ᔚ�,���N~�b7
3�[�ǌ�������z捣|r���� �nY�h����@�k����+�LS8�6���m�CE �\J��A���xwkW��^�����=���O��Y4����JD��q�����V�I���i����2h���٣1\w_Y�Z$����Fu���X�u�6�í�񩑟�p�e��i����&����}�!��xG�.�,�� �?*et���%;���F&@>�R!�Z��7�x����x���|��*�x;�d7�uC��e>��$�����}d6�26�b*��R@o���2��qZ�F4*(1H��:����@rx��=��i�5@�IP0������dayq�o�--<@|�B�2�o���J(v�e �+�T�@e�n��H��jJ8�� ���2ю�؇��F7D�/�ܫ~����?O/N�L����?�k�y�)��d!��"F�؆�Hɐ.�d$��
�Ej���Q�nˬ���s�ҋ(�N&	��bhbA0�'�\�e�ʎ��;������Ƣo)���&��+VH�ˏ����^BDz���9"P��$���_;c���<�=0~{��z5�d[�~g��j	�5!�Ԃ�Z9>h��*�&C�uW~��������a���Q��`n�J*�
o���M
��r���x vZ}a[��Z���kr>PD�5\�E���%��Ri�T�c�L���.s��o �*���Yo'sD{�`ʀqH,W+����dۆ�͙���$����}!5�TF*�:ጟ2�L���^f_1�
n����\�g����S�ч1%P�Xq��3�T�����J�&pe����ߞ�dy��ܭ��g`�[��q0;BY=s�f�ĬƯU���}�o���L�;���˲��p�&���n��cpWM�s�zn�h-̤��(�C�s��Ú���d_�~�[�[갠ͯy8Ĝ>��in��ޢ��u���fu�l��������Pqf_��\ ���F�<�*�uVt���Ŵ�ZiQY'艛��[�N��vy�V��D��vJ��*��?����S���U��?�x9I;��ݪ�+p|�����)&Z�.g_�Ș�F�%0�-r
bo*D�~MV��Y���+�DgJ�X����!z���P�B *�]A{�����\\��k�'��ӛ/F?�2;v�oP�����Q�^����u�L�"�^}�/?����:�j�P؃ңq5�B�jj�	�䛆�]�bD� �[*̀��K�!O>�b�(ڪ�b �?��xä0�axse��~�n栌8m��J#ϩ����{��7�Ƈw�8\N�8[�)B����|���)Jϧ >��J�r�>Q8�����$� �զs��|��w{�$q�kꢀ�A�=Ղ1�'O��6ѝ0������N�N?4>x[�!luo������jϐD#�Þ�6�;)D���$a�'w�Z����_&��i����2�f��M:�el�0���>�%K6���obp�z���p<���C�
����]Еn�`q��M�d��P