��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk�����:@����L���by�H5��;\J�[��m�,�� B�%�]��s�,�.Z,1:׋�Q�w�]��x�SN5JK����\�W������'ճ��n)�9�Ss�>R/���A��x^;���t?�wF���	��T9)�Zz�k��޼��&nB�{�:�`1D����>���<��7G7�W�x�y�Ȅ���w�R�@�'��O'Xҁ�A�xqH,� �l�;�ds�o*��q'�。n�	�|;!7�?ͧ��Z�ܥ�q���DKH��Bz�˭�G��\��m�ԥȌy"��4L���[o�b��v*���۳�M�철Ɂh,�aʶ��2��+ȨGcZu���h��g)�./�8t���{���Yլ��,U�I�Iޤ����϶oM{�o�p
�����L��z���*��x�|���Mꥥ�K��?(
��g1/�=��r{  *�>.���N����n\hԻ-n�$Y��]$H�v7 zd~�6<�ò�]�9���Y����dp̣��%5ЮƼ9���~�W!����\�V�谰��[�K�T�\ɐ7W`��b�ޔV3��\�#���s�%}��I[��j�x�BE~���FHC�7�z�gN�2��BR��U�1���by~9B�Bڢ�u��UX�)�`�Z�t�-e[N�\ˍ�[=�,6G���B
(z�Q��7P��v�MbE���z�.�}�m�u���n*G��O9��鄱J���ȟ8gt�8EI�Y<��Q\3�Ls �9#~єԃ�f�'�k+�Ң�U��}�b���`çr
��evF��m��������&�+1	����A����6�H��K��~1�f�P�x���WR��T���WZ���<*>��[B}����cq�J,���2�%w�`�x�d.���LW��O�#���(�+�	*�1UC�&�8߻	�.�)�D���og�ꕒ�B�և_Vp(ِ>�;����pmj��I�C����h�`E���1���Pe�o�x��X����k}J��G\��ɹ�0-EF67h����P��r�(��e��A]��a�3�80�c�[Rq4΋lnÜ�UĽhb����|Aތ��,�m��Q�1���4?u�\{�k�>��W�����Z#���ۚ_O��ʃ�/Sj�t���Ī0@p*]��3��_ ��_�$����
���d��E ��w+�Ƙ�sl%툃�Z5�)\]�zbR���*��fi��]r��89R���̢��}z��~��2��ug��>��x38�@�7��h:�!߈�LG8N{�QD��Z�4��w�]��z�^�NQRV�6�NM��}�TߺȈ��ߪ�eIp4S�4��5�\l�����
�Pi(}X\D�Ȭ��!!��b`�������������l]|/R ��X�Bf��vV�2>����Ճq��U��^ӥ�l��C��g��lݣ��K�A	��N!�g�fm ^;Yg�T�B��c]8�s��k�b���^��t���C\��+��ވ²XB��M��w���zn#��C5)Xe
_F��G����ۢv6�RN�� h��}��}�q�����6gF�x*�$�b�0blB[!���mR</������ƭ�/�6�XF�B�2VY�9g� yNI(�?����m
������#.C�_����j�J�h�ؖ�ے ]��ڦ$�w�4{���i8\�� �?`�|��+cۗ�1p#��|˳bxfr�S�3�nK8P]�ٶr�8��}�����2n_�4(q��'v#���X��5����d���t���<������vNɔ1n���Qީ���eۚ�2+N�U�`ĵ�Y)����X��DP#���t�@�����Oo�?у���مͮ�[2(0Ǳ�������'�&*�����>\/�ٹų���D����Kd�,Q$ЊQP�C7eu(& �=����������v�5ޱ�k`5*�x
�[_�0#���F��/d���pSZ���V�]��B�Qp�����l�E�@΂:6sen��d����M<.K��e^��sI�g�8�6� 6uy �.��t@7�$K�"�9����)� �c	�P�bM�\��hd�ȭ#�����S��,�"�t���4��ʩv�)�A�2Y�-Tm]jF��n�{y�oo�Џf�2`��ÂT�w�^|d��a`%�7\�G{����>�J#����4x��~Ϯ��1V��x�Li4�~��o����|A|6E:~$B὘��]��I���!)
��we�퐰A�4] z���&nʻ& ?�*��:�gSxTR:��<��`��`
�HHɀ'�og9�;�|5v����e^��-o�4L��Ǌ��wV�F��F���~����_��o_�:�}	�N�X`�#&���οg�!�Z2ܔގ�d��9GT�wf��V�^����v���v��j�L6W3�~�~���'�k�U<M~\�9ן����r�L��&�+d�#�$\(�W;�m�s����s108�)E�J��w(6r��cGf�o���)F�mh;"��]
<+���O�PB;v�[�1�7�ꉲ�׌�Bg��\|ɾj��	��D�H+S�D�Z�6���u����
��4��{ʛŸ�����߲k�����j߽H@�V�k�k*0�)�:�Dx���)g;˴��kY��{��lh?����\ ⸢�dL����[���ՉQ"��'���q��[����cIN�}MЁ"�M+d�;R(�}O ɷ=O�E�a�nGY}����5vE����= |L1�٣j.�.K��Y#�[����Z���a��X!�^�`d��O˔q}��@z���`�3�Ϳ�L�Z�uG���D��`(��毲�X���1l4���eT�l����_C��/3�**X���\��@��19 v/Z˱��S\!��c�^�&�l&
����y҈K���-�k0�z3�O����q�.�T=-h)�eX��:Ԁf�r�����.8��Q��r���X��X`�S5T����r��^_�u��I��}Ď��D^��#s
����m�򉇉� ��[�V��Q��2p�