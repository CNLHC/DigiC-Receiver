��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���>%���wޠ��X�aq�c�|���j��l��Ϟc�!{�Y6�z��^mՏ���!T�T�?��.[����<�C�Z�)��79<]	�i���
E�~諟��q!q$70tU��d�h_:�����P��#��HT��9������x(��U�B�Ku�.���9��D�����JS�����<�׻^+(�+�}�{�"�.��Gx�Aѷ_\j��D����\P��͒fg;E|L�݆��?
؟��"��K2����u�����B�	�%B��M�h���l.��u`!��T����%����7���SG۠�P"K����O�ɋ���`ߙ8��`�w��d	+8dr�	nL�wx@�&��ه����U$�<f�+�&�M��k<���e>u/@_N"���΅:k��Z��k�x
b��͝�����pQ�t���;�,kӋ�br�1_n��K]�!σ��2S�&5;�9���K'E�J9P�\�R]�Kj\�?a�
����k"BD9ٞxd��/R�JSd��Z��|9���ގ_+�\I��Z��i!4�m��n�:ǲ���(X��ն��d�$eS�.�jk�ڒ���R�q���c&�aBȱ`E����)s�BA=�x�����Lj�N��s؊W�����NW��j�BJ��y[����s����;[żK~W��q � �Bŉ�z9�2C�}1ج���yXܦߎ�����2*}[U`�*;�g��_���u��b�w �m~?�Ʃ�Q�{i���{���E��2���#*f��(�ȷ Hi4�%�И��']��|B�ݴ���w@��LN*� ����
��a��&��])�U?C@�3?�OC�ꦙ9U��n�+V_}��
ƥݳDT�g�0�&K���'���|��%�B`!8��XVݣ[N�w�!_�g�,���a����9E�KIk�-�����<��&�YU=�b�l*]#����\OF�붵y*.��>V[�߳Q7��=u������C^D�Dy���J���_�\��T�M�\8��N���}��L��J�)?���e?a�\���3��h���OR����kV�¬)��?��6�"#�&L=��=�i�~n���z�o�����Jԭp�ҶPU��y
Ǆ(���^]�����P���on�0�X^f|!u�Ii�a;�/�w���,#,e���v����7�W�r=��Ԅ<���y�_�"h��1�C�5�g4بZ�Z��S���ux�˹���Z7*�����|1�]���PŶ��Z����Y���}9���s]�WEs��ꭒ��K#l�2Kn:ݖ���]Ƚ���#{�4y�v%�Za��W��ip���RE&��X+�[��p��n�a�����=20E�Y,&�P���$G�}/\��C��H�JV�2�׽�I4qp�l��{�����_q�0������;�\�N|h<����/��O{\L��1�{��]>r7k�:��ry�uX(��l��͒a�9Pm>1�g��s��nge4���p}�gi��z�=��vl�b�����?>P�ܬ��
�<�)�M� �vP�U:�i8�ϲ����w�V�1o����L�"%�J���A��;�U*$�R���]���A~_����i�7�����$e�i#��Qx�׃0�c�}��X��]��D���t�Z����{�%e^Љ��9k�f��X�==\zf�mv��Y��J�ҙ���~e�S�;�Zdt I��	�4
I;��Yxy>����WZ!��0:G���(����Mx��c�W���O��������$s�@���ߟ�����{��Ɓ��o�9�^tHN����3��W�B�aD{6�������qtP�E�߅���X�LNO޾����/:6�W�y�,ĩ^DD�
LIaZ��T53ϭ[K��u/��lEz3v�ˁ�Ԟ�h�N��+W�ip�����I�$��Ԙٮ�����ʹd�7���a�G Mo��� �y�yp5��]d���������n�O������̸�J������Z�$��;�>(��1��
��)� ����z���ą�oK�����-���!�x��	`]
��p�' ��AA��-m�^�������6��j��_������y�tUY�91G�C52�v�W��b��d��x��ԣ��z�VJ\��5����LU,o�Ise<��s�.W����f�@<?�V���cB�H'[m�@fQ�v#-=���J's���g�g�3���O�h�+N]��	3ܘR׊��k`�7ў�l��yk��6��.����v�U[�\;�K��X�j�P���u�Rh����FG.�}YvjT�>Dz���5��_~c�]�L?�({�J<��������(��>��T�طͣj�kB����4,#C!����1,�GAV����,�c�(���⧆���>�L::�Ql�]0-@��l�0�J�#���M)w�/Qs�_�n���m6��c�L!\f%�sh�v��^E�Q�#he�
�f�S�b x<Jr+��@W�#R�p�S̙>����5�z�bg�)q�I������E2�9�}RB�����`h��HJ�@wQ#�x�PD��)���b�̜������5����w1�61\] GǸ���0��s�E�/�T��K�-�FB��>����F�Ǐ��/�Q�2� Fr�.���EIu�����Y���+�#6z�ֲ,EN�\oE�W����e����t������޼��@P��ƌ�~�s!@	����wI�CX��:U-l_��N^��:�s��i��ǟR��i�]���(���;0_/���ɵr߈市��eC�����?Ђ�ɇN)���L�����`Vf�O�@J+���K��\�\Mjj��p�P�y��uB{BK��xl"���f{*��Z{�lZ�ge�H�6��}�ź"�{b��
�[�/����Τ��#���_�umu����T�17D�.�|�uʏ�kEH�|��ex!7��F��@[���'8���]:D��ֳW��[���B���N7���[Z>\���"	X?�z>��H��#��Ij�Z��nX�R�.�ӢQ����te۫bf�_���_�K4�0}�@M2���b�Z�i�A����8�@M_Qɕ�ċ���痆X���6�x�=\K��Ǚ�d�K	��J<��Ὧ���o3���	ԙ����y-�@�1�-���}=Bz��n[�cWp$�y*<֌8����5���5�Iṕ���G�5��0���t�j�?��X�#�[Q�\p����C(R3������j�#�����cGXw�`�
�n8����2�Fg�qLI,N���{��"�u���9�j�#[<��o�Э���d�t�,B>Ꞝ��K��*6P�v�j%.�JYy�����|��ZGd�H��4����Y�3v�5����f�)�]�!QiWNpx���q��1��� L�-�^�Tܼ
=)�u|��k�N�T+*R�׿��m^�C�O�Y\��i��0��Ơ	c��ZR�u��I)������|��AH�I:�E?:�2�W��m�U���
���"�*�	࣮^�uւ�yR2 ���;.�	=���������'�?�Q��vn*�f�Z
x/�Zu$"���V���+]�n�������V=Nir����C׺����!2ђ�הig&�˻a��H�s��Z���mN��|����F/@��+��Y�u9]�>��'��y��2����<:la�-�}�k�G9V�<�ƛT5G)��S	n�Т���!I�Y��)��U!�5�[L:Q����P7s�IuL�S���V9���&J�����+G��M����L��W�l`��`B�� `l�>�P���8�c��u��2� �*�;6� �и�ah�_��Z��LІ���Yw:����E�;3����E�řq�ҿ��t	�d�Fl$�P��8,Ҟ^/�SC�� �mR�L�(ˀ�K<Ӟ=��6+��M7�u**5���#5���9}���R tAШvJx�z����'�P��+�C��q�V����Z����ƣش����?9X�?�G;��h\Yw���4��vƅ4��T��i�RWވ��d�v(q|�p[��uc����
 4����1M��ϝ#V`��oQ�S{g�~J=���5�y2���Q����u^&1�|�b��Uv���VG�N�ğ�zw	�R��F�v��8�CJ՜t���IcG@��4���h��N�����ޛ��E��d`L�E���%��gڜ�+i�~�]|�*�@�p�)cm;Ȗ,w\9����CT:,w\�7�Wl*->����O\��Q]�̬�y�P������&���"�;Z�%����?d��WY�h�]n�a9R�;�����*_M:�*�t �P�a>W��L�Z�����$�i�3��ͦЊU7�6���ؾ�ڴ�G-�v)��1�٫F����(VW�RhQ�[�b"qGə����kGU~�Lw��j�/��5��� !�wN�$C�5I�7>ePVo�ba�^D"犐��ӛ��1� �*CO��_��ş�:/�ag�ܜ�C����6�N��(o#�T
vjj�Z�7������.���fl3����߅�;I����:ٍ�W���^��^�>�#��c�c���>���Z��w�4��˛�o��^ƌ�PUr�Q����UWm��n�E�\��E5ך�mUd�J��k8Y���#�yj�����z0cc�*���bqL|#�?��7L��'�������. z����Q��sEnwd_�HSh�eҊs�*9_�~܂�,�OB�I0�ƶ3����V�o�c��eк�hU��q<��/���S`x$�}�O|��\v�°X{�}S0�k�	#�ݘ�bM'���&��s��iF�����3�4I���	؋��ޚ�o�_CI4.l?�KtsBU�����5���J��wԵ���a\Xi�I��u�mQ~_��,\jĖdu��Xn,����h)��vD<ĺ���6�y��JӦ��3�o	�J�o�be#��t�!m壔G�T��}���	�ہ�<�Ԃ�2§!�z�z�!e���J1�z�t���m��I^���Q���)���x+Ga,�Z��\Ha��I�g�пG�!�0Ȃ���0�\#�Tl[^��z�bS���t�iS�D�x��M�<�I(3*�*m��Jy�H�_�d�y �a"M�O������^�3{G�!��GH�X鬺�f�$P:B�S��־���5�8q�}H�!�!��:!����ֈ�	Ї��r8O��p����
̘"/����I� �>=F���j����Ϊd�_K8#���J��C�����Q@k����x)���Ƴ�p��231�-6�7���_b�B���Am�!����O�Xڠ<����ь.T[-s�Qc3B�q�/̨BT�z_�Y��8r��ࢤ���!�����郏��k��'�0�f�(�����3�	:��FM���Cp�|bX�/������=�h����;�-E��>��JPl�u�?�����3�G:�D����UQ�T�C��I�c6a�i�+�W{�bF���_�Wc�͵�#I$�^��ꉢӑ<$¿��T�ZT���a��f�E�~�v۰C)�p�C.ّ���b���
.4A���g!�<�Ϝ��IpD�m$I����V�^����F=�����O~��#��R�S���+�S�*��Un�A�QTl癹j�N��Y���z[�!BCo�Rb�YYM}�����5n���o"�G s[��E�i����9�#���e��<�m h�;��@-}�����4���b�6!BRT!��
��5���P��%�N@Z�������\��Z�%KB�ҝ*��<��dŜ�4�V�@��f��vLͽM������N]�ꞛ��!��;�b��u����Β�#~�>�O���}p�#	jZ,E&����)[�eu���������Ԓ��J���l2��F2����h��h���{��q����k~��g5IX_���<�;�Pg���p�	6����5��>�`�}0|o&k
0�ֆ��)�������o���
����%ym�`��ņbƟ�A=Lz$�'z���V���sA>���H ��{ ذӶ��<FV��F�V��w�"�X9�g��v�j�������`�ߴ��Y�j��T#�T9��Rh��8C%��x:�B��iL��a�c&��(���~�L���DbaSX%9|APi�W�?% ja�{/Б�Y=n�e�ܶ�B��V��[����)>ou�W�ʸ5�2]l�3LKR �"�	n^�%�\yP�иe�f�Im�/xd#B@��)�k@�1zWy&=S��B�k*�I^M=M<�F���$nZ��vy�pc��t�ߠQ��]���p{w4F�<��աV�fM>�����nao�-�f�J�Q��-��*�	*6*����{U���Q9R7:T��P��Q���a��#H�4�N�W6N84®5ie��Q���BPV�kj�0V.����-��qD���a����R�.{�qh�.�f�
���T�D�7���#-�5t�)�9���l��ʄQ
�_�X!�q�wd��vu��!��{eCv��J���Y��h����?����S���P�f��G�
�J���a�k��k�3�@���nt,F1R�p���\K��3����C�C�o$��6�:Af���S;w���@6���87%�z��C���0�<v��$�8l�m&����A��WQz���_�[�JH}d��n����P�F)XA����%�g.,0a#o�� 4��-l�R��Y�Z��V�[0��fQ�A���ha��;h�P�a��X��T�B%�8�&q8���]|�k<��k����li�����R�1u.+c�Y���{&�)<�$�P�?��y<�)i6i���㤃�<B�"L#9w���K_虣��[�L�߇�Q�� �vk�#���r��X��0Tǅ��D]>	;���3��ǎlF��B��	M^�,G���rYXzA~��׎��,���k}��Ӏ����Ϙx������!`~��h�ܱQJ�&�r~1n��J.~�F��p�y ���R���i1"`-^��z�|��%�d����c����??_�&"��
�1�(��K�*'����Z<w{GY
����r[i#�S��U�ɞ��HjC�dͧ37��?�(�0d���A4���Ө�܄$��� �I�S%*/������!��T�?��8�l��A����>�S�(������B7/�.�� �rc��5�V�������K�>!<�����2(�����)z��8YT�M��N� =k�tZWt�x�c���E���T�2U�37����@މ;i�7���$�#˪��x������L�hn��L�t��P�|� A���?��	W�C�q7��rM�EIHx��T����ާf�==��i���7˾��ip*e��>,�M��$��+�Rk[�����1s�Y�2'��=���ʌc��0!ֿ���g�Vܴ��cy�ԣ���?i�7��Yz�n�V�{���뮮{��M���^V�U�d[�L���@��oDtQ_n�[d&F��%�U��Xc��K��4Q���U������_��&�
}M1���{�feǵb�N,)ݐ=ެ��;����Om��6����d�>�V-49�4��!�������=kv��ǌ�=y���]h�=Wsv�ǩ���;+�:���K%���{YW��5{R)�T�OOIIx3T�#*�D���1�x�V`��k3���+�9�Hi{\�T*ډ�	t�R�}z���#��i�\�y��k$1�%?��@�iGk�E��������,xi��h���ٗ/����Zw����j�Ū絊ܾM�A����;��("��lY�zhT��z�d�yT�"�@�=-�靈ZA{���V����C��'�9�I�d��,WM���,'��:/�ҿ���\�<��8������%����w�𭙞o��8F���������l�����h����e�����!���§�(��wh"��w�3�݊�!à��!&�!���0/��@����s8��%*Ő5�,�uc�Շ��S�M(K�2���s���>�ARb��
o�ay�M��ֺR���"{��O%��7�Pl "�.�+A����&�_�x�hrd��ol\f_`b��x���������O	����9�%P�4������&C\Z��Ͽ�>�o�C��,�AȆ9�0{n����Ԭ�1����m�~s�E����z�A>//ەɊ��s�0���^�$~������G���hjIe�{а!��@|�|����m�i��"��e��#.�S�?H��\�}�lQn����h���e���H�جW���RDR6ՍA���忞{oh��}�퉅6���_t�̒�P�T�Y�I.a�s����ā���As$�*�0����C���q��6�K}:���$iy��g�"��"E �t�	�Lm���%.������)'��P{�G�o"�/^�$hN]X}"����b�4�)�^q]`_���BI���2�qG�MC��wj[g�V˟2��'8(�.38�0V|`6hy����af{��L;��v��,�ZX9�������~�G�Ѐ�����{x��p�]�;�[�	�:=X`�v�"�W:e�26��y�射1�D���O��+�����t@3�"��D�	�Mo�'�2,�$��v��}Ign��ے ��lRO�A΄N� �_ �<	$Qu��7��i����,b-a(�d0y���/b�KXu��_ҁ6��PbJ_!FP�|��A^���g�1I�엖9¨��SS���nľU��'j����b�:fG�[c|�0�&���)/��B�ȞW�ꑫ%1�㔴t�*���(��ŷ�/�%̏g���U��}�(.�0 Ы�Yc��ɻ�M)h`��WDð�<f}ń��ͬa�G����h�O}���`Sp*|={Ȉ�\H:f�{R�U*۵[I�TɑFf�2ۖ�/��PsY1���i!c�5�H�׆� 	�q.���S��>�E�9�UT���!��.�.����BJJ8�˒� �����_Ȓ6���B�{����Ό8s�u��=OK�n�|]a|]+�|�ӡ��<b����N������)�
���dr�p@ ��F���M�f�@DJ����B#	87����}����W��w�!��H����(��H2�!��g&��t
��Mq K��JR���2b�����ϔY��H�|uu<5ُ���Q���EYm0PV�dYzY�%�2?�I��M��Jĺ��+�7ڤ4s�:�D�;y��p���Ub&ՊY�\)� j�{�Y�;�v~6�_��vVS�f��g2D&���<~�~����F��7��
51D�$�e6x3M��͞���M�v�A��e��?�;���ޠW7�����z#�4�ۥ��6@!���dW%&��W�p@��r ���.��S¿��Cl3js�v�@�����1�ĺlV��1�|����O���Ѿ�v��,�գ�P��/��
AG��KR%PlZ�Yf���w�ɹ��њ�O���^�����	q�tx�ϔ�A!��:O��{O�9�	҃&�F+�t��Bi�o�&��wV^��«�a�䍱�Ӣyu��o&[��U�	�y�2���g�}8+�t�BJ6	`�=�psL̈́˧�+p�sh��;�QT97h�R��`V�!� M�7���~V\6 69����/f`�L�|A����1-U��om ��[c�/"��t�Ғ�(�1�iB�Ł�~D� ��o�Ҡ�9~�3Nx�����@^��+��ϭO����wEu�!y��A<	y�<\��>>w38���k��>��sv�M2�8�Ë}�@r�#N��`�G��N	�z7U�6����֎+u^�v���1�E%�熜�d��pr/8O,[~�0�m�@K�­	���Tk����\}�;c�
GI����9v�RՕeRV�F_|?��&F��-�k���
�}��n#��WW�~C��&���!<���1��&��L��rȄ�iA����)�#�:V=��wMcP��i���ˇ{*#Rn3��@8h1��}���-A�MZ{��Q��}m0�GW���3�.�(���h"Nu5NҐ+{������ȠC{+�cSN���;�V<`��Q̣���P!��m��#�@���q�s�����9�|��<#���R9t��� d�U�Ee�F���r:������,Z��vlզ3e �G�#�R�y﷭�y,jn��/}� ��(���{d߫������5Q/�l��Ƭ�8�}� k