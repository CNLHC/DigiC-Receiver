��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk�㣪�����V��}�DW��RO��,�"Z�U[T0��A���z�3@T���H��F]�����,�IA�z*�� <��&Ar���G���;o_�z@��ƪ�
p\�6}܀R}�qD�ѻ1��p��n��ɣQ+��hV�ޑ6�2�����rm��>��L������f�gf��B��@\"���_�#e/Ou�H�6\�-3i<s�cBu��>�k�9L)� �^�0Y}��FO�5����
h��%���;��(��?��&��:T���X�gJ	I��j�Bf�9ŉp*�j��+J��6;�w�]V��0�b蕵�{~�~�K���j�LbF�[��{a'��г4z��+��XH�\�u?�Rrd�K�@�:��1�87y�Dp��?�{���G���w�y6)_����6�ْ!�f8��!ܿx��O�ck����֭�[��N\X�Xe�+rV���i9��ʧ�8�"�P6S�pc}$���A��ǇS����%��&+��vjJXF=�5�o�gg���y һK�fgSټi|_�]�k����޷.ۡ}O}1�l#|������;�Pe%#	s�%�I+�A�1�E>�E�&�]_�|Kz$�t6&�n��8��'L�#�Р1���!��eE$q��pg��r��S��2�<����u�_%m� �M���O�{ڼ�w{�!%�I���W�6 +H[��U�o���B��&���]�Î6��z��;��LM�؁:&���M*�;\;�(�B�F�5�K����W�Y�h��R�in��nK�r���h�����W���I��V�ϼ���A���>������:@lu�?_
�cR�aXq:�0��A0���E{M��.)�𭂲X{�z9�� h鉣訬�f��R��S��V6�
0��J��J�K��� �|�+�!�58K�Y��/ �j?�p����7xnY�5FP����u@F�_.�qg�$3�^�Ϊ�V]����яLJ���Z��R�T�g+�RۃjA�&�&V�P�K*Q�^�����$ꓬB=�!jr��� Q�*~��W���@1�殺��Z��-D]�q�W��;��(UX�����X�VM~4)�c
N�Y����>G�7��*�?��欄`D:�6V�����t�OR@�U�t��!�vUY�pL �Bh��j�炖��~���Z�6�j�ߧt�>��k�E��(Ȕ�y�w"�)z���vT'2)eǰ���M�л�M	���=�ZӐ���4e���rw�>�w3!�����K�z|zc������'6�sM8���ll�U���m�ѐu�F?xG�}��ǥ�\,]�ư$*�8i���(��˯�@b�����`�?Y� �"����l�Z)JWrZ �
p�e�a�%Zb3�A�O?k#�X���x��Ti�0~��g<�x��^���ϩ�Nc�C���^J1��Lŗ�����,�����1lNa��i����	���[ٶ�����b��"�ek�.9x� ]�X$熇&�=!�uO��̏�=�Dh�Ҥ���4�5�Bb�Ҡ�]�G��@��}�L�C�ÈR��Ѫܲ(@��Re/��C#�X�@�P	 E�s1@EP�$:�v�V4D��'���u0}�y�%�Ɗ=~ݛ���S��� ^���~�H9ي��[�95���K�'^��V{��v	~\�df�Ic�U�Q���R !h���@�ǔ��H�v}�>	��]�E��N,���P�\�v�bqsnR&�u�>���"ZY����~�oa��� �/���?�r��mON��)�(�#�ل��1�'Z������(�#v����
ކ^�t��]�=�r�9?1���]&�C�3�Q����떏�iͥH��ds�'�V�=�0�"m�H���4l]P��������o�(v>NUt�Q��uP	/����/�A��ME��vj��#%I4���3�U\(�$�S�c�X:�R$�[��|��Z����# ���;�_/�y
�=3R�[�+S+s�*I]{��S<<���X���*�ώ[��ڰBU�v��t�c�@l*�O��)ع$TUV/�e���5Mm)
�:&�F���{�$W��!L)͖�he��vn2�[�`r���r@j��u��j(�Hw���ĪӸ�z_��r�z�F�{�/��pa�V�zZ�\��)fM��HE�2�5]����Q����c�#��2�������B6��ǣ�����uq�)�
�@�׿S���(b�&�͓�M�V�[���77��L�Ts�9a���YPp�i 
�7s��͐;r����dMX\�fg=��mjǝ�w�\��̈�
��-V56�l3��E�h[u��������NJ��=>��F�W���b�����׉�r&eX�l�yQ��Yۉ���ˍ�Pf<XqF�������Dk������Ǔ�b��/%8��R��ߣ�1N����w�yc���s����+#=Jq)�ؐ%�h�Aጦ���Y�(qJ4�9p�Ha[}M `.�?�6��p��0a^�߳9%�y-w�1��L����a=�cET�A�{��=��؞�����R��fʈ��ƴ�.�|,��RrM����m]���@W��]���Me�5#-���7��˙�vAcnE�KZ�t�O��
0Al�!�cZ�@$�^�>c�,,8b�9YT�jF�[��Dsl�T
��y���D��Մ�������)|����V�>XT0K}J@�jo�~�5B��;*6��5pd�z3���qE��ne�o�A�l3���@8�ӬC��J1`V>
�I��%A@�U*��r�0a:��"#�wr�XE�C$�`C��CN�W, �ۅ���C̞t��LǙ���q��_����㓖�dGs��z�u��b)B\$ǗT�.��3n�0���Vf�;%ɉ]���K��F'D*��s����}|q=9'.�Q��#�Th��>H{�����z��J�wZ�9Pw��9��+��8�k_�_j �u.L	O�^�%5���bƛ�n^6���
�O�զ��g�V��GϜ1��値�)���!�������0�H�j] ����?�-��h��ղ2i2��:+}դ	���eH���@]z`C�U�&�_d=�(U��� \�����79��l���E}�b�6����N��\����G�닢4-��A�Tfx�P�[K|��g��L%��N�����qk�ၫ�%?z���S�Ҥó�.�u�J�F�i ���[dݮ!��;�I����9�X� ����'ڂ�6T4��o����kP�`���ލ��XN-�	��S�����8!�H�(�2\�����v��u|�qF��vT�y��E@�����DC�;G":Y�pu"(5|Q��5�LymJKH�������.��K�*h�l�
ex>M+��1��X��u9�co�Z
�晕Y*t��o�*��e�����T��7��Z(N �&v���\���+�[x��W��-�t1Kh߬�$	@���Q�A}<H��'(�R��D�چ,�в�~�5��٬ �2���d���O)�L�3!�e�K����Lk�g�׸��*�ʅk:���ئ�I^E:̛#�;�St�@pS�Lxʗ���K��r�{V#w�a��� �xayN��]9��W[7��A�A[��,�}�S`Ӿ�}��]�:w�j������N-��qO���|��Y��t�T)��7S�5R:��L+:P�$ȓ�{oy(1���y�@���>���V �i^�K�)�����|������~��˳z����\A��/��*���f�S5���Y	���Ta��k��΍��H��z�b��7���I� �H<�D}u] �:��[��C�7��mH�63�DDp�La�{i8��}QaГn�_�<+0-�H�>Z�0���Q#�-�5���*���.�u���(5�d���G�Q���7Z%�ǋD[!a����(�Um�U��7Z��d���:
���f.����c�!rNp�S9�����X��7^�����t����bM��${>WȢ�M�z$ X�m_��ٰ�=ɏZK�=���8�r$�`-��^��ԗ�pD_i��~:��(�'\�o5:6�Gt�a�{��hk��	�r��ލw���N�ĤL��N��4GW��KaHK��.����'p���f�}����v$;֮���h����a�ME�(�%��$�n���!
������3\��_�-�S��c���yO��W�A�+�r�Kd
��g�����@�����(e���IO�̩�9�(�1�����x�EA$n{�(o����!mV(��_�HL��)��-A 6jY-ɱ��#7oꨰ���;�AXwR�]�tIt{����tr�3���gG����
jo	GJ��"+Vb�-Hx3J��2��N��㓥1��Nu�ՠ��Gv��WU��6,��p�����N�Q�&ϕLr�GS���x����0S�ZD �kW]y&<�<�����\8���v$Q�T�y{��|�Da�Q��`��SmPr[&�����#P}�f!ٲ�.�a�=��C���j��V�C�֟/�ز*O���� 1�)�bݘ0���r��SS/7s2woՄ�Iл�[����U���]�����.)F�>@B�v�֝��K�kp�Vc�z���L3�l����F��R�_j+P_��a��>�ǋō���j����JQ"a=�\�s�
��=:E!BPN�u���F}��S{1�e�M.��HD�H
�}�ۘ�ޙ�)Хt�޶ 1��e�bK#���JP5�f��z$�(�<RZ��&:'����[�n0+��h0E�үZG�Gi�2 �$��}g����ā�y��8�� Sɽ��̋A~"�4F���j���z:�T`��b��J߄�u�X`6ރ_m>�U>����>�>�R�Z,m�:�L[�4s����aQ׿eɜ8|�A|ԩG����h+q���Ba��23�:�1�����n��f������m%pg�~����'��S���?�ӄ��1��Y����*jc�2�9�旐3F�=�h��[�����+Ib�4r#�m�/R3�
*���H�R���>��~�y�!0����r���ԍ5��	��0�Mb���Y����^'�c���'��J4mn>{a�Q�}n��.Q�t	X ���n=��x�%�픣�-k,���
Ȥfq\
�\"/;&�C�L��.)s�A�ɶ�i���(#(�����o]$z�K�R��=�gӄ�8��yR7�@G�a��f��s�J��ŕ�������7x�Oԝ3:o�hEq��97S\O�TR���5dF�6X#̝�_�8�Ϫ"ԕMqR�r�923�^�%��`Ӄ|2����5��3����^�-��� ����Hi��㷛��F�yK�!y�&�S��gH��8���i����q���ɷOiW@�w}��� �� @,���*��ph�Ȑ<3%h�tq���b\��8�� �vT���	�.#77���A[P��R)y���7ej`e6���&S��	mA�W��s�����L���Xꊃ�@P\������i#hG�׈�����,q�Vݗ����@�K��ٵ֤ ���.�6��م�o랣�uߋ+-��Re����0v�&>�4����Z� �$Rh�<Rg�[.��iG��ZR��t$�zܣ���C�Sz�i��-$gD)�Oݥ4���et�vV���!�x�?gS���s�`��P���Ћ��8�#���J%R�Y)6��-���AL��`�=@d5a���OT��r0rW]O��MU�N�wCo-���T�g��H�Ɇd�u����������#����㓇 �8f*'9�q.jd��\Q~�*P��@q�G�@�g�F-��S�i�e�騡�5~��{a�A���� �ly���<���C-�⊥7x��"�"�w16�5A�]cs9�Hr�L�������3����E��v^����w/2�4��Y����`؝�_Z�~�� �O<�A�*��Ʊֳ_5Sk7'�;ԩ�^��vŊ�5����}��� e�X����MG�[Qb)�<�t�ÿ�h�-ʠ�}��y�P��-;x�%k����=�x�R4օԧm�X�1�9���㱬��wџB����1mI:D0.�&& rM�ͣq�k�澍#Z#�B��|��;$�8���"U����'�#>�l��SZy8lX��_��->��jn�IoWZ�Dy׍�ǚ�3!U�pk��4� ��+����� dC|������*�N��ʇ��5Q�_��=�K��| �
�U����1����K�X�ש++࿍zj�Y�ɘ�®"Q&U ��I����V�f�K�yE�r�]}����W���F���|�ݧ?��7��������5j+��\)��N>]����*I�!l�2p��&h�P��d H� N�������_%Hw۵�m��ڶ���i{"Zk�����0���_��pOT��m����w;���ﲵ�8������uX�s���ٻ<Q.���7a��p�8�j�܍R�m�$�-Zu�2�3�R[/���UG�5�<�)8suƦ�����y�
+s�z02��3�`U���t��r���;L
�~�޲�ѱ���� `[�o8[Q�����@]�E
�a�����w��{t��H�8�Cdȿٳ�#���.�o����D��^]�g�m5�4�p�}P6Q�e:��7֭����p�ĸt�q�Ų�^<
�h��*���BHJ��)��_�n�	� ���܇��p��aVem��5z�p]�W�'9�����lR+0����%G���vě�7���gu�4r`͔b�$7f�H�Oo��O�O��s^at!�6 5�a���g ���W�r6�Jwq����N����� � ���4f&�I�DWr�{����sߟ�����c���;������\�fZ	r�O����K�F����`���I�\b� /[�}p>�	&;�'�A�/��k�ξ҄h��7G�+�}/�x�B�"o���4s�������##���8dGje&A݊�4���@;G�+պC�� Y���I�mS0S��\;ؚ�"#��@P�!�~�ˡA��_ &���e 	�Fk��}C�\8_V�]N2j3����Sk�Z#�m�����߰����2}�>r/:�6���y�>/sl�H%�d+���*YK�3$�Wk���zn_�cg�K9ޚ%i1-�W��ha���� �M�7\jǜg�+(�КxaGa�<9j��FO���CZ=���%�?u$nj�yBf�2�]�P�VʹF��K׍m�Tm�S��U���\�.*�yM��wj�W��^u<���"8�����i�L�V��ƕs@�^nyT�Os�	�MI��oX�S���uF�M���`��W�f���g�J�K,kI�������R��,0G���$^J'V�*ę�J|"�V���}<�!�Q��٘������堷B���r�K����n��bn4�b��z�1�xz�م�G��ڄ�4�B����"U��d�W{5U�� 2�;r�\�l�����0�oz;�v��/�9��bu�`������P͚n�oN.(˻ϥ�$l!�5�tP�!УQO��-Iً���;�"d����V��s �����ca��Z"&���Q,��Ӛ^�i5���������a0&�?v���k�(�L�3 �rm�Q��z!܃�B�\�J�/�v���$�!,��4]y=y�q� +X��iƐ�!�Ó�g8TFI@(��Ib�
�Ԧ���`q�:�Ϟ���1g,���.��"�v�OW�B5������m�!����Y����]��J�H�J�H�?����-��/�tMUp+0_���< �DAƩ
Ŀ,��͹�Q������Y�2�~x',�����?G��DĊ�8�Iߋ��Go��cѓf�r�?���Q���AHl΋�MO����Qd�O�i������9I��ES%*���;���6����ς�\c+N�8�u�U�qg*5�BNg��Q6fq�l4�r�ъ�~b�sV/�9a)��5���+��a9��H�\���j���H�lV��B�Q���e�d�����S��� ʉ�6�r��X���W�� ��`�����:��I�5n'c3��A�.9Ȃ���o�[?%s���)���m�%�6_����9��JX9����?HC�=�������-�|XV�-�ůPE��_�7��� �����dP;�2���{��}��ޡ4z8Dc �y���5�e|w>���_�<�?��n�r'V�2
��(�Z9��ݢ�Э'ǝFU�~~��m�P�XWO��n��d�M�KEK:o位���5Nq�����oE��cw �p�vgsQ��[%N�T�[t���0U���N$f4S�8}C�*K�°��%n;�ظh������h�"G-���k���YL�ԧ[���;�]N�Y8�e=�*;')�NN��W�BK�v<�?6_����ԗ��+f�|�ŵ��L1�������I͏�����߁Y��^���w'�q�$T��T���r�o�M���x�E��_�	�z�g�k�-�R��rZ?�Ɯ���C�﫱8>T`�]���.�li4����.+�"k��ă>AZ�+`bf�-�*|΍�Һ����k̒#��Xvy8��|Y��C� ��J�B�a�n���~���AvS��J��L��A1W�-]k�}lT��@W�r=�t���ͫ�������S�qW�hA�� ER+9�}r��b�798�b�=e�{��_���P�k��ؕ�iadS5wX�$�&R���D�I���'By��3�S��������:��f���w�d�=�}W�Ax�,?9m`t��]J���>�>T�^Gaཹ4�O���kf��vgǽ�7�KM����k����t6�SAla&���o��iF:�AQ�?@��
�DI�D�֋���^VTJ�N��5�n���n�����O�-�j�� �>"z���9�G�?752O�HK�Tcsi	˦�G?���f'4E��T9�?[�ʫ����K o3��������V�2+�LB�g?#'!�~G}�Q Sio��q��:�&䆠G:��|�lUI]PH�G~M�<�l˺�~�4m�fJ拏li�elנ���0s��a}7��x>��۶���H+����F���m
�nb~L��{`���~�G�o8(P�@:���n���� ��Y͏��~3��:��wXmy��Fd����	?������ʅ8m[��h�x���C5����;5{þ��� �[�z�ttԞ��Է����6����ޖ���5�S���#�;��S�*�}L���b�6ty��*�m+@l�����_��,@�hU��^��+�N��Բ�	��h��>���d)3� 2'�7��2o�^�=]QF�zCH�j�4���UL��wI�䆁a|�/W�k �5ni�`�!�U�=og����1ЭE�ܶ&�cϣ�����Ǽ���N_���r`�?Iܳ�F���>D�j�Zӏ���g\�9��#���h�s��Z��~ )�v�w>�vaz'�0Y�>�Z*+9����+&��֫������tgs��؀~<F6����M�0��L,�	��W?�����*'q�\\�2����O"�c-�	����Q��{/��p��ӷ�s/銒]��pX��#��=�|�sUr����>���󂱱P�rpSA�f`�X���>��.���|�-Z�^���j��9a陉� y���O��yarY��f`�\�EcRK�#�d�}��{��9q*�Mk3Ω�C���!�>�@�u�/u�������$5���FnPM7a��m�@z��p_�������M�J�� ���柲r�����F�Y�|Xڕ��O��e�<�(]�,1���gG��g[uSy�b��ulsN�h�HR�����6�vޒ��is�G�K75$J��C�e"Z�3!ݫj%���c�N��X�C�����o�o?�Q�rd��&ݔH0-�j�7�xn���})�+�C�ד� ����9~�! ��t�����U����[�6���/Ӊ��z�()$��Zd\�`[Q���0	���y5������p<�d�Sǽ�Hɏ�_-5]���/��8��ť��r���wŪ�ҧ?��~u��Eg����va�/_#�%���p���"�w�ZE��RK_�E"�2�m��)ұ1$)��Y\P	��r�hĦ�^{ur�|��B�6���I��p�1��H'��	h��e�
��i����r�1 "N/��PM�5��TUp�r��{T#(�[��m����b�$�V�8�oG��]b1̯t�ث�};k�Cޛ,����5^���n�����!���V?H9�-��&۲R�7;��{o3�ː۝aV�*�U��d�Z�6���^7���xb�;|�t�,	$�J�YݗX�;������1�!ro%�X�ֶ��On*��#�*����sl-ȟ�nuy�����Iw�y|)�KJBևn�Ga?��9S&�]9(I}gA�v�#��3ÆP> ׇZy��1;q��������Bb�����\ɸ��&$\�ـ��� *�aHsU	����Q��5�0ae>���H�_��kC�W���0���}��a�5 ZD��g��$:%HJ��0M��2]�u��~�q�v���6A�A��.|�ƻ�#�Q~[Q����w7��bG��]ҷ�Ď?"���Xx3�ҥ��w��E�S`S+�s�������Y�FY��L�m��W��#I��M����`��Ƥ��=ć�l��t��?�M����I5Z�vxbX�<y�#�  b�_�������`��k�i�'Ahc�n��Q��
D��62�(����)�D�ch�Fqr��h^�*;��<hir�|����b����6�M���P� �
��*}l�No �@7wel]�-Z��ǐ[ߩ
�C!��rO2�	��M�"���5�_��K�zG�cٳ����X6fC9���J@�EP&���#��A5U��I�z�a����b�k���%U����f䏒d>�%w�fV��73�?l�aV�c	������o���ǰ>���i�f.7�L���Q��P^�
�O?r&@U���K��L���Ib��(��5p�K*�9��vy�>:���r�5S�����WV������������H�D���^�I1�lr�����~���:{ʽ�`��*�:�3���RuѶ8��G<sT�}�k# �.#��c��I�;[�b�S1��~���Ca���@�������='Y�M2Ci����m�B��8� �Ƙ���T����RF7j;/��R�G܎'�3�=��g�]�F)}��9�|y�3�e��pAx���y~�TՉ�A�׈V�\WOkt�R���Em�eNiu�at�Z5&�O�]&������2Zҝ T�hh�y`J
'x�5_�R�Ȝ�Ӂ4���L��`v1ѓͭŶ��x&��r���́���̎X4f�ķ[�Wf}�(��S@�����q.	��P� {�p�3۾��Ry�[�mN�DD]mcѳ{@�>A^~�W��P��{y��͢�"yƵǮ�EAR1S|(L!�u3���y�A!��E�d�]ŭH���	�x]�ǜX�@e&�;*ģ;�9�ꓜ�h���܉�j�8)#;��*c.���L�	/�]!��p��d/��,� ��a�z���Z[}S!��
�z>g'2e�g����6rY��;ܘ�3�%W�������WX���n`�ȅ}��o�&Gp���b
�a���t9g��]�H��L5�
9<��|m�q��=���So\��kxV@�?��l]_��Ve��Fӻ-����b�~��K��u�Ƈ��}l�*��)���w��YsO�c��".���ք��9�+I�H��`M�v�����&��aW�x�B�W��4�u��{I��Gld��C_� �D��{���#����l����߹�Zi}���]�?ȿ�{Ib� �g��?<]x���$ڶVFf������1���$<9���%Z�|^L\ڨ��c����=���s���mF���t[� �0WG!�P��G������R�'@7��#(��_ww�,-��lp	��)�]������=P;V8���v�2P�;�8�P�9_����*KqnL#^:����@���T�����͹���0e�@��%?�^��: �?5�}mZ�����%��0'��s���+�tw�uh�J��`�����r�oR��
w��A����4�������#�:��z�Jn��,�NXh^�0H9q�>�� ��P���I�B_���^�Y���V�$��~h��	�_
�T$�nbؾL�,�/�kԦ�ɲ��~*�`�cdRWԌ�ǄlƠAMրg�p���59&k>�ЩC�FA�.~�~�.��]�@��z�
E�=��O���?4;c3�Ӛ&m����f�'�d��AUR�����N��E�k�Ь���O�u��-�����	���~����/bjG�;���Ś-��F�uiW���O^�JNc�5y����g8��%Z�.� =
�aKҠk��@�E�a��q�%X� ̀F�FaZ���g"o���E�^oW:�r�P��){�JCX��>����= '��@&����M���ih�e��!�hC�j�?��0���_�gF���Y��H*�?M�෕�x�e�ou}�W��	9�o�F��wo�G����m�ߚH���*��D? E���bHKs���Z4�p5¢f�#!���
՜`�tF:� ���%F�>ٰD�#A�2��s�u�&�BRHNw"¡/^�A0��+Q�	��~R7E.��\|c�ʊ��]��}y&)��Rh^��#��6� �+�1s�n"��4;�I4�F�jO�uV�λ�'\Ap�Y}&���6�l��Y��|�v&;�W�[��ݾq'�K2\W��J��}ROA����⡧"��`�bI7'<>+No�����[v*G��!�W�şY`����0�=�Vx�{��{�~�kU�sS9郂��j�)jX'�������/�m��yH 0@@�A�3	�Lt��K	�����6����^X'(�j����U�7&B��.#"��[�z1�kCB��v�OvO&��m�BM�o��1:�vx�SF�<���]�$��]�g���!3�	7�P�g����d��q_����C3�y�gv<�����Lq���˵���?�B+�,Q ha?�d��W�7�u���p���b�x�1��qj�P��EFјM%��$�n�B$��`� ɞ�R[���}o4�C�<T��^sXk0Y�@: �Uጾ�T�jh��X��#�	jA�ܡ���b��E��tT�3�#������ǒ6��Z��+�qG�P��r�@`%���_ZU�wI�`b�:���u��c��`Z��E�$��ۓ_A	��;�s~[�~,<?��a�K���8�'&���\B܂Jhv��u�^ݍ�P����;i�f+���"��'����/��)����� ��^�V׹i>�s-S����!u�,�j�N�;�����y����V��������:%���>=�&PK��:'���w�)
ؑI{[��\�,?�Ľ��Y(1�$ڙռ+���+\)������~G�10.:W��� �G��R��C���z*�����P���%< X���uMv#�|i�4�������is/��W��A/��� VX�%Y����G�=(zd��)K��On��%� �rz%�}Z��w|`�=���J	}�"}��皮�W��j"��ĲOO=tD�{�Ҭp����1�HX��R��Fy����Ys��^�gy|���L}�	�1
�����=��r��"ڧ��3�H�
��.6"73< ��=���,��	����/
;Ot�FQ~o�R}��	Ѿ�?
���E�43���`g̈́|7�Hm�/ۧ��c@
[U>ƺ�{3�M䶐E�~�v�	��=�)�%����g10;�I�Q��a�#��C��� ��������9Q-C����!��λ�������Fj7>��d�aĵ��*v���g����؎�8r���U��U���m3�<%�ڷ��n8}E�MKv��I�*������c%mSMfFG�f�]1=[�5T��s���Wz���� ӷ{�=$��KM��-;��=fl�t�̙�kh0D��m*2��?�Z8k�W*����}[�/`p{M�9����&���ܗP(���O䏼����;%6��x�o�Uw��4�eU��_��>]����2�f�j�.IH�?[i^E�I y��+��y�l�n&��������NE��
L���KV��Q,��Bk���iS@����];O|{�j���c��cy��0C����j}�ݻfAձa�1�����x�yW'j�V�Zk��UrMbf�A�;��?�h�i���}[�3:���ط�>e㚙;�3�����"�7�ά ��2=�m���Q�3���i^jq�cr[L�x�N�����',䖝R���B_�1�g{�.E�3+��S���4��|9rJ8}�:��xi�n�����ӄ:�Խ�-J
r�܁_j��V��[.���I�8�2r��	g/�<��o٩]-������-�/,�fd?������T���QS�w�{���EA`*_;�=�ü�c�?�U��oQz::�	��1c���y� ��?G6y�=���e�tJX8ף����w�}{<���f��(?����<��N�`�>㏌�x*u!NQ�����*�#�2b3���y�� �v11b�_]�� .�_�Jq�)'Z�b=����a�u�d>��އ���@�D�(���Ώ�R�ID��ʧ]΃���t]��3� �-���x-S+������ȇ��I&�=�n�����JU²�G���d������x�"�pM=�4@bX�'��������\u��l��Q�Mo1h�5ol>�I�7
_��L�7:2�7[c�����m�G�Ï[��m�=&h��()C�_��������z$2�,E�	����sx$t�z\���U��&����ֲ/��p�]��Ŀwָ��kG�#��Ĺ<�g�S�5�����~@�o��n<<GU?���DO�"�����~ot�u�CU�z�:~ɹ{���+7���������_��a|��Q��$[>yQ�x���?���u n�����H���r y^�!Iu�]2-�\��uCU�%,����#����\Q3�ح$ ]I�-:)�N���vtq��)4�O�v�T��������VW}[U�� �:GV揺ˤ��.��K@��EV�MӼ��9=���),�
C����_�Ϭ�g!ɾ:1�ar[�E�O�4�&����JU'q� ��/���
͏���,.g6uU)�R��>���]6f�J�СЛt��T{^�D[mS +)b==��K^R��%��`I��BL?��[����A��)����\4�|���M�2{���b]�A�&�e�~Y�bI���S�_�	-�˝�_ӿ��R����5��G�E�c/�?�|:J��Σ���
��t���s��Գ�%�*�h)�����B_F�,�0�+�e&Ѓ��j����Sk&Ngk�z�PM,so@t�~S(�w�&v�ŕ��w�vLu��U$��Uf��ϰ��}R�yQ7~.qF��J��3�mIL���F��1�("��$��+�%���X�&_�;���No"���Ba��	�1oH�Z{�#�Z��j}&s��D�6~���C��#��Q�{$O}k�E�R����Z���_�3�A
���YB��J�J����T����[��֕��#�����$�9d�0��&�h�E3����������<�&!δ�G�8M�8�=�kK@����3l��|='J�A93�?m�Ԋ\��NC��d�l�b��_!!���q����o׼�cɡ~� �	�9�$?����zRI��d���� ������Q44z�A�|�3�;�����{[i�f�A����q^-%��r�V�^��2ޞ�/����C�x
�tAc � ��ʛF�<�T��m� 5R�����o�Z�>JM�HIR�u���o������A��:�uf�x�����&�ax�"� 
,f���P>u��{Uj�����d]Y��aI+�Q1osO���$~����s42x���w���μ��rF��0-]~З��j(�~����ou��t�b����(D��KG�<K�U�|/�\�V��eH�^b!�گ����g�?m�$����{�R������86G�L�i����c5��Ì�3���-������l���.�T��v��Z�w�W��Պaz�z�W<G@m��q�5-���jY��};K?�(J%�Fv\0�	��[3���Î� �(	$���V	0�PI W��7�K�]-�'-xz�U��S7����`��c������;��tG�w�t�f��bu�]n�$�<�*u�'?�T�)��@s���%����������߼ÌHк��y��,�(0j�W���wV���g$ZsS�1�hb���ُKeK�PH'i�k��Q��S�-��(�}���O��.G�Eu s�k�&�Ď#�m��S��yk��D���
��gƇʥ�z1��`�6�vӑ�l�<Z:�Q�_3��0��H���cf�nBga�We�����u�c������x�����z���n����E�J�@V������t���P����������_И�%��/��[FH �S�Txsp���:�� Ïn.̔ol�� ��O�i.�L�~�D�u�A��6�v��.����}��r=l"{f����\�K�POSG&�2��t��I��o$�	}m��a!�Ũp׳�MY���HR�1N̜�׭�Et��e�-���ȉ��C�oH�#�n�-K2 �N|��9i`L�SP���J�r��cA�fߒwm�q=r�-2���s�_RڋJ�J�w7�{Ue.��56��R�ن���(�U<�2Ù��>��n��,��[)��{Q_�$�t9��E��V�OV��W�)�@G#p��6�φl�w+�tl��o����@�w~��C�}e��v����WbJFJ׍ÒY`�[m}SG��H�<o��H��Q:``�?K�gT�Os/KR���ݨ�T?�G^�mnfU堠�> �S��0���0 �#�p�J��w���'8{5�	#(�2Vⴕ�F�o��ǭ�=����f��v�{9Z�Ts�߮��~;����!XH�"�r)$8������*^#�lI�!�@�����s'6�������v�"�6Z쐀�U�Fu͝ޙ���PY�>Q3�6��{k�&)M�ˋgܛRv�h�ɗ=8�\�7�9H��V�˵r�ν���u��cq6�Е� U�|=��]��R�q�p5��D0�iҮ������r�)l�E��DQ����2S��"��ӭ��E��P�"�\�&4�Uff|����־�T�ݥ�)�s,�_p�2 kǁ�%w�&MS����]C�sG��Y�f�j�)�͆�g�$��_hdr�V	�Z :]�q��
D^)�[ڼn��nCw�G<�j���©��d5t6T��U2��"P?0їֽ��f�e����?�Q�~f�k@)�PT0�e�u�Ii��Y��"")1��$�d������*�(��v�&���)��\{����@0�a
���o\aN�P�)i�-�k􌹄�8�U���'�d ����Z�N�ϡ��
h/��	�X����:>F:�po���	��Z�&a���~�}���T���{0Lj���b>蚥�8S|��]����7�/�5A�B���M�k4���PG�
���hZI�&g~���,�qpX�`��ߨ��ı��2������qGn����[ma,�lt���8L���{.�[I"$K̰$��x��Rv�.�q��E�L<^I%�
�aQ�6��mw�uT��$��u�N����p��<���o�q%�g�)��,�a1:�q5/��O�����*��E܄� o`��,�H��X��<Wj!��l�aA�5�̆}tWz�!Cp���y�������g#�|��R�,�Ժ��D|H�������hcQ�E9��`��qw�F�&'�l�e�z�ɹ�Kb��)���q ���ۇ94���h�5���Wa`'@/~�v5A=�]�F<��$V�W��k��H�(����X�\�����3bs���Q#����-&����f��d�������)�)��!���g������_����0x�-��a��gz乶"Q���N���N�v��6e��_��-�̳L�6˗;2R��N�Y�T�2x(P<Z���{VK�R
z��fYan��ޠ��O��kf��_ͩY���v�`�#�k�T����(��(c���*�Bu_�w��
B�j�� �Z���ۢ5�Y�AT�n�����Q(#/�s�|������-�<M)�Z�����rT��k0���kL���Z'�@D.��i^��J�� #f|'h�*�!��yf�H��=���t�[-E`ji��'lU�m!	o��F�c����&f�4x�o9�X����~�+��Fƥ�oڦ�-H/N+�4Z7\�9��G���D�pt�6<��>$����"/Vh	#��r���kl)��?���
��"���=�OW8�������d@o i\8`ZU�`*�SX�k�Ũ��54/S��H�7w�rق���n�$O�Ώv�*�X��B�c~�����P�P]
�v�[��<�p��X�j�m�6(�j�|�������A�3d��.��t��U�?��x���
���q��U���JoM�h��$
/��YK�(Ͽ�1V�5j/��)����{vY�/g���W"l	h����y˂.'N0�V���T�XeSzzgi&<�F2-�;)�n�u�;w>���+�@-,y�%����
���3�gzQ���_]�����5+����X��O���.c"���)�����(���t�4wM~U��R�w��}g{���x�x�������Ym��e��:�ao�8�AH�dϳ��%�5���Q,L�11�x�R����ޘ���:=��ή��֑���Ř��on�ז}��#��N?a���B�Si��kR����eu�e�^����i���Xg���&\Q0��܆D��J��݉�㤹Dl�j?�Î�*�븂[� V�N���"F�E	H0��!?偨n`�]1��nCq���G�ℚqo�*2��s�%�� �&2������@�i�������ә���H�f��~yK+�>y���E
�E�TP��!=n��(l�\ۯ$��9�������^/�R_�`_�׉��)��]֣�����j�U�rX3;��D#�1˯ќ�N�&�i�<��F��L�.G��sXԲV��^�x�7<��	�5�#�����)�A$C��Hfw6)��K�#��dm�[�\��H\�����x�T0���֮���؈�3�A�{��4��(�Q�Wq��+饟��}TIJ����wvy�����sM��������&�B�`�]���@��R��o�"|�A�m?4C7"�I�ی\5��k���ž)�K�t\𝺕�&����/̠�ے!���!��
˼0͟ԭЉ�ZA�u�Ֆ�����R̵C�d����̐M�c�����M��˂��[0U"��L1��
z|� ��D������<���
��:���+�M����h�������n��M���"Rs����nJ� 3�"��1N߄02.Y^$ή@~�o���񸓙V��`�ϴm�M�x^'�� S潐s�{����Ә:��=��r��3UxqDY���:������oZ�lD�]����&GkI+�H[�lL�z[�A-�I��9�n����?�>�3$�s��Y;n�+��ֽ�~&@+�RX����1��f��C����O��u0D��E2˞�aR���-:�l����X�$�②ϊ�.T�~6Ep��uʺh�'��t�sX�OEx{�ܜ���;���/�\�ٿǠ�,�9�H���Ֆ���8���A�2F��X���2+8������2����L�b_c�ў�v}�Q�R�ENK؃�Fs��w�s�Ř[�"�V��$^,���&��+�����n�Ac�#z7.o�:��yС�U��ʵ�FC�K����G�榝����t���g{�.�d�0<:~z'���猱�T_�Z� �'\»;~�$hHAm��T��zc-�ڥ,.�.J��~�ҍtF���q��;?pMf5H|��h,��7�M��T�����s���e
��6p\B#�Y3��j�)�t�����F�g0��ѩ�)���
ַ�Zb��i��T��3�4�6ߌ�o��r�˜����~ϴ�I�D�&Ǌ^�>����ּO�	���jAɐZ�B�UtC�=^��Hg6���d5Q��G�����kJ=��1�>-��y@^�GW��9!i1ϛ���������)�3��HZ(SѾ@@���)����~��_õKjH�`����cm�`���B ����TY�)�pB(��}̰_�/�W(��3�A4$���egJ`_�m��G*�ݗ�q�K��"E���.b��{��Y�9��L9խ���וv*"J�b�����>�L\�S����@Y�[@e!Wy9�R�G>Y�]� ���-C	���� �t߉� �Y�Q9l�e���X�xի�0�ݿeA��S�b����]����b��ˇ�� �� ��S��c�����qo�&��R�@�"/���)��N�8��Ǵ8��5�.�E�ji��*��CڟE��xB��Z	2�ڷ��ǩ<o���m�հ�/+�+ N���zˤ�bBΟ�C������v�m��mGY8��o�3F�vq��'�o���1��7���Z2��K Ը�Ǵ�R����f��wͭ0�JŽ_:�=e;����H]��8y6Y.���ʀd�|��������H8ݹ�1��[�<���c��b��9��w��k���#�_�H�W2I��6FU�s�V���zP�|�d���i�������?Z	r��+��o�	|�z�7NN�� �;����+f
l�(E�\tihn&��۾��gY�
��H�%k^d����v�Z�?p�B��+�m �`K����Wy��Cd7X7�c���r�WMIQ3<�����G�	��f�i�"Rnc�CrH�l�7,��eU�m�U�� C ק�T�B�|��p�9�I����v��oV���g0;v�v�p7�̃2������)}(g�5����2�u��hvL���"�.�w*8kjݩ���Z��8��+hH�&��Z�7ˑ��hޛ�����d,3�_h���eC$�<�4���.�#h���21w����߳�ئ��İ$2�W��C�m,���4�`������C�ӥVU��
?�d�O�:�?V�]��:Cr�p���(\��W���}Rlm�g�OC.% 
�$8�,KäҎ�?�&?c�:'�c	y��������]��T�}�)$���5ɛk����8I�-�P��x��:0.���ɚ{BXݝ�V]eqV���6�e����?FO��J88�^3���b<,��0�B�+Z�O@�j����h�us���A��H��$����(��gK(�K�Md�ɍ�/�8�6��<�+ahu�2tH�yko���b#g!��\A-zuB37\�k��6�m�/rƝݳ�H��!2,r`0�N#�w��d�ٌD?�������no�w�+����'�����U�4/���*�\UR�����8#�gy�{�[��SN����+G��p�ޏ3Izb��y�],C�������*��1#��A1���  ����I���rõ�ї�Έ'��5y���e�pq�>��ΧK1{��jV�3�&���D�� �/x�]�#���bt|�g$Vo�^(��O˒��0�K�]�)�L�MP�������TB(o�2�wU�T�ŝ���8�| ʱ��Zu��N�0+���p�B���b������&W+/�y!,�b/,]H�p(�A����~cž�E$0-��e�ǘ��%��'ے_�pt��Y ��r����w�W\0q��nJ������o)����K�dr�j����'C��n�;l��jEz�GV�ϟ�n�w5p�u�5�����Q�[]�e#��g�Si�~ˮ����ֳO��ևle�U�|�Gh�R�֭ a�����P��cRo������PK�Ȍg`W�l`*��EZ�a^��R���[����P��*�[�֋n�u8J?V38Ax�O�D�$7J�52]8������PKg�M4M0�i���qBM�?wյ���5�wm'xj2�Y�9
�q��a���CЎB�fb�:f�}��*/a&-�!��:4To>�ϲ��Ι
���Jກ� Nl��u������l?���"�)�3{���ռ�ac����B��[��B�F\���j���@������g��$�D��WZ�qEp=�����K���r�[�F�D����P끾��(%TC���J8�ᑀ��2��� �����8�V@�ei-�@��f#[:��c[��#�	����I�ƴQ�Cd<1IzW�j$W���BaE2YVw@�l�r�:9������:����-�����4���G��7�y(����G,G��o�N��T�Z��J����ת}r K��*Ә�.M�K��(�ף�k�
>�2��(ѱ"��ߎ�����z�ò[oy�?RArn���`QK����h�b1֓���"/���w/�R��c	Z~���Ӹ��=�Z:���<���I���F��M`b��� �˽7�����o~d��@��I�Le�&q�?����Ơ�or�ֆx+�ؐ��v�*_�p\Fu�i`R���q��x#e~�p]�lm�
�R�o���F`�v̶hxՈoX�&� �ѲVt7A�nr�bȜ>�:�i��u3�D�<���P�o�ֻ�ǎ'�I�B����m����#��´q��1�� �0S�p��z��R�&� !���*hj�U�d�@�����҇Hwe���&c���3]; B>�9�G���)�M��1ȶ��S�9��lղ�7�n�d�#��N���K��፾Ks8)�\#GΒ�v�����+�}���2���5�P.�L�\��#}Ԉ�H�W�E��oa�Q��UDc>��/��5{P��*���Չ�; D>�����5�d�h����^���|&~�}1��j���C���<D& �Ţ�>�yX�A�6�nKJ�jE�ӎ�0�e��?Ч % W�9zwި��gI�C�o*�%:��\�.m����������K'i�2�ɦ��J0I&0�Y{^,�uye����wF��!av�Kf�����$-�>�j���
��{���I)N쯣q�܆+���er�w|"���� �h��)?)9�v;ܨ����s�A??�- T6?���1��
 )�8�ZQ�iEا��1�-&TCV=eA/dg��D�<G~��9I=%��}E�B�C��-�+��s��n���f{,�C�j�lDV�����
u���ݧ������ 3nI�K;�N�==�����)�t��� ��k�� C�����q�҆�6lm�p�'�}%�[QTtn	?���}_K2�Q�k�W���n�j��3��OaVLZ�P�������y1y������6������9w��퉶��5�V���9�]�JR��ߺ[�����/��{��	J��:n�b������9�2�/ճ��y��9W�s��T�C�2�c�X�;A"�HQ$[P�"��&"Nr1��/��[�s�A�I�	� ��;�Yi��3��{��b���k��� ��'8h�˅���́)��0��Ρ�a�Q?8@���G���r@t�!w��P�hW��mK)������H	�Ɉf~w\|i��	�#T�fF�a��]� lSL� r��-�t|�:���U���`��g��QV+�1t�>*{����Ȼǖ���%o��e��׊
���<�?	V� ���ءʔ��5��ɴ�^#�zD۱ʼp�[H��K��	����+�̟�����$(��C�[������7�`o�&Ck��N���Z�,�>*{�>V0�Xs�D�����D��XZm����G���x�W�b����j,s-��y�
�/4%�X	�_y5Q�IXa!�qR%���/t��)�*T|x��쀉 Q��Ү�v��%�t��J;���$��{w�RPG��'J�c�F�Y^�]���˂�M��`� 4'%f�N�mpk"х�M݁E>��:�W�(��A�O��_(���ش��K �뇁�!l��?x5�'Br�W;J�r��K�x�~&$���)�oU���he�� ��q1w�/5�ډ �HD8�<��ɶ�3Зkp<Ja��o���<����3|��n�cʞ�,�ʽ%��##Fgc�v����� �$�� Jl�Ip�8}$�~�(�IխW�2��)3{��t�G�%(!���X%i8�,��X#.���qe��Y���f����"�������7�zWE�Y�棈��{xlZ;��I�M��\�٬y�����X

�U�枼��[�T��l
Y��Ug}ӔY��S�*v��e�-'o�����_Z*.��;��R�F�����aS�E;c����>���L����^�5���e���[*�i�Ί.����sߓ9TN�G��.%4(�D�8�yBۗ����C�Ls�5zUAf]եh4U�+뿞F>�=�d'a�O9��M:G2W�I����\D$�F��4���	�E�Eſ"��0�n�K��,-.�o�QNS�$��uo�p]�6��fA�B >�ϛ]z�ƣ7$��~(�q�S��t��a������3�dM�Èߏ�1�
��q[�$V�ݚ�cQ;���lՊ�P��M�V�Fzٗ�����Θ��[�W�ú,��ǾNY�M�cx/���[դM�<�e� �-苃a�*�9(tt�*�5a���}M�wk��$9K��	L�����6���\{���T���2�z�7� �9d�igU�G���@�"<%Gtdj�۬�t?.�~'�8�@	p��k�蛌=�;4:1�A�}1	`L^����g!d�ܻ=w3�e�N�;�)�X^+*H�q�%�/�y�Ft�ζ�'�_�@p5��H�3Myb��*	݇��8yM�r5�=�#��c�<����Cm�ZC�W��E�B.ְ�*�zW�������,Ј�r�ۣ}E�� A�����T��~�k5G�x�^˩� ��9$�Y�a��Њ�}̇bo���u�U~* �� � �~B���v�k��'i�L�8����Ɵr]�����;�%
qHF�B���� XٗLT!��ܲ0w
�5H���io����CJ�������(f4	��Db�͓��2�܈�sX�+$=�v��:a�l3�?�E~W��F�ۅ��i"Ϡg�`cˍwd~б��՗�Z\r�S[��L�Mb�M����#&ǽ��us#YB��js��9)��}K��Ԡ��2۟�c1�:Vr�9t�{��E�u,�.�,jR��y��[�� ԴC>�m��{��y-�9��H��v����:\�Oq<����Y� C{�����]0�}�#�%Ҷ_�
Nuo������%2�G��T/=�a��\��<l'j֍�^���K�}��8@�+�}yMi�O��z��#)P'��Q�|�2�^K�z�Aܧ:�OIp_���<&�ќ���|0K��|)��%)����@���2�\V6��eU�Ǩf�w��z<��[��1��(��*��
]��V���$7�����I��>����2�"��YL;��5�{�5oNs&�?jtdQ�SӜ[�����@������G'���ޥ#��Ė�@�C��G��\r�ȇ�e��d_������U��󇤈	q�ߍ?󋻔�T�Ej�3ۧ
�\� ��B���5�ܺ�u��f�3��r�W��qn�#��q�4��RP�Sj�Q�Ҷ��n��n� ��H�Qys�O $�\��8��R܀������ݛ���hP)W�V��}��<Y����[��@�Khg�Օ�6I�� (�ss�va�&�r0
hi$)�Q}8!=�
�]����+F��h�Kӻ1����0^�b���^@���Ea�����uS+�+)``�h~�L�=�����/'�11F�5�1g�P�����C��'�m\>�&���"�`���~#��{�"g#�ygv^*�s\pS+?Q�e�""�OY��oG�?;O�/YٽϾ��Y7��
�CO=��	�K��Q\\<&�1�nj=D=H�m��k����s�֡R�x� ���W���~xk"�;�����z!q#0�y}T��c��)"��rO�t=�5i�l����PMg�k������ən�\�����P�^�@@q�{:�&�)��t����ú�wA�m����	�>M���aI��GNP�R�W �o���X���kc�"{&B��m�⛾������Ƽ�wȕ}b�P���8G� ���:#
�_�t��<��Oñ}��~BJt1��uQ�GIW+O��x�|7o�k��]��Ƌ=I�����c:�� ������b���L��!?�q:*%P86(���.�����0�X@|�\��S�BI/U��\cʦ��#���yF�!?<͇���k�E�U|����ڐ^r{Zڨm�:��昂��X� �L;�56���c�y�W.Pq���ڳ�3z:�Fą�4L��ؖ>cT�J�F�Rw}z���[Qm�CCt�oMPS��N�e7`�x>�gIȢ�K?b����������М]q[M��	�m��6Y�/�1�k�sK}��5�0��� �@����^�B�4�)��a�LM�
�N���'���'(K[D������B%��ܟE��r<dvh,�n��y�F��V�_��j�˻x8	'�oY��1G"y'� ����"X�(H� QD��[�]�q:����:��w����e|c�;l�t��T@*�e(k�6��R��e3�~���}�[`QIx�g�6���3!S��A>��Щ����Q���ܽ'�Lc�C�2��J�ܟ��A�i�6��.�?�n�Sј���y�Y�"�-��8io*�$��1�����(-�v�pq�Q�<�/ 
>g��<ֵ�/'�Trz	�!����-�����|��BƧ���H2����(UN�Ie�{�h'��C�c��x1gy�0t�Y#)�,��+U/
[ď�Tp`�@�U��V�F4��O��x�.��ه}����kօ8u�p���}~D��Kx��(��hc��*IjVXO�����
Bo4��TT��o��qJ,D<�x%�!�5���7��7*�����6�u�A6��B�=n��W|ʗ;g�zG]�?X�@Ґ��,
���t�"I��B[�<ixo!me�GɊ��v�znw�������]2�Yn	&L�/%��"~i�8ӳBg���R�{ ��Tr�;R��	'��;a7�f˾�V�tJ�֧�����G��ۿu���8�|��Z,R��wu3��]�0���];�d��3KAs�ϽK��<�҂wXC�%�[�d[I�j�qa�ԧ=q�+��T�r,�� W	��=�DD�+�7�5C�)���E��9�i�b�V�3Ovd�rU��k;�I�J_����ː���x/���J%��F���������j�q��qKءel)�YMCg�}�{��b}+~�0\��W�d�?�@�?(�7�I��R �7��LZ[$�"XQ�	t��ԯHc���2�cy �G\�Z*A�����.*�q���Ky�&3�!ӳ�I��n˦��*�GU�'R�D��AR*��܍�\��_giq�n(O�];��-������ٓ-H�踭����~�Li�\���:
9)&�G43��_���y[0��೪��I�<_�\-z]��dP�[��,WZ�\��tȍ	d��>���:���0J�����cI��V;ݝWs��������!�'f�Z���~<�U\_p��o�1���x�q�mv�hC|��7�u����^Uf�o��n�!��}@����'��Z�Voo��
�Jș���r�f����L��v���l�Qsz���<jb�55�d����JK'�!�:zI
�lZ�Y�Ҕ��ui#+E2.�[AU��Lz?� �q���������4U	ЋR��@��f��7�Έ2�Ŝ��ݛ\�P܁\nj�b0 �&$����aaF��V��m� ����_na�Ě�\�<2� �8��:��K]�� �>^�҅���}b�1�*r�䫯�X�M�:փ�4�B�-�T��-�mv�X���3�蛤W�4�L8��,�T�Y�\B�Q�Q��Y��p8>c���9$����SɤrD�q�@T��%h��X\;y�IlP�gԦ�&��Ьq���2��.����U)�:�i��[3��wA@�+�*�}��}��]S��U�,فl����o�ݙ��t��������O�$�c��X{ݏ�x�ώγS���(X�H��9M6�^��A�O��D_"Ț������u��!y�K�������=�r�.k$��Uyւc�.4��F�-k�W�f�	��e��X����:W��zFS	'BYo�1�������}Du�a��xޕ�K��?8I��z6jW��IT��O�lc�&�>������K��������o4��Y)�̛ h��~9��[�1c�"���b�H�����]�}���p�Q��.�r\��;_>F�\ B�M��zy�j_�� pz'"4�dKO�fj;?��I��� �����k���e��1�hD��:�)��][>ݚο�!Q�'ޡ�d�).Ͼ�o`��`���^�j�!���tf2,�P/onw??�7����"+A�{=���y�׉��y��QAGvlH!�.�9=Ϡ n���A���n�<�|�OƖj��Q�M\�-�����{?����"��d�B.'�c{y��ɸS�a�f�|J��;��y*^ea;�
��l�C�r'{m�~�H�c0ta���C'��]�E�9�p���W�Sd\��'�0j�]�!.�cJ��0Ƥ,^&bZ�<bgm��/~Di�*����@,YY���@�ũ�����5L��폽�GW�އѤ�z��
iM*t��	ʴ�|��]t������B�jY����[��X<�[��;����)7�x.���dJ�huH�CI��;�~>�@P`V�W��4�P�I��n�q�wf���,�lx�zQ�TX~�h7̈�'��2���)3c�P����[$��Q(c�9*��w%9V&�����x�zŪ6c�M�AH,��NWmk�v��Eh5w"�p�����z�C������x.DEW@�t
#FT[�J����Udqw�]��I��l���݉��6W��b��[޶��gxtN��Aҿ7z���CAg���[企:�Ӳ�Vt�F3��(��V��<���a��@�����rB���4 X���A�a$25��H�9�E��W��f�X�w.;)�T=Y�vr�r��q1:��~6�`D��㞺3grP^�ː*�|Ўۖ�ă�w��؀WF`�����{��	v��4w������{�,~*٥�k%��]�&Ӑ��	��4N$sQ)
И�%��%~:I��x��)�h!�[zՃ2��nkz��#}ߚ�ug~��Ó�)[�"��dO�͜�W�/ƒ%��m��p�(�!)��4f�6�C�>�v��4h6�S��|���Q�C4-��z2w͛������XzƪT|�`$�H����Y�}�| �Vڱ��P���D6/���F6 ��kXNc+�G��L[#��4 ��A-�ܦ��10�<�F��&$S�#�p{#[Yz􈰜�ֽ�}=nG��d�@bŷi�ٿ�j��b���49x2��~�<L>MC�&��`|�%LԊT��(*�AT��K�Ś{����ܘ'�ݿ��쥺�K��@��-�t���1��Y�[�m:���*���2��߄T��9�N��?1�)�ч���v�&�j��y�]T��\�=w(�QW���"R�bv{��Ǻ�kT�����q��� ���'���֮���Ly�;�d��Ƒ����JS�6���K� 	8p[��{�
+��5����'h~��D��iWa��Ӑ��Z�$���*KՍ��*=ʝ���(W#3��3���F�,�]���W����Л�g'=H����;Cu/��x��c��n�Ѱ�e�Ȁ8�5O��p^y�G�$|DlB�TERM+�\I`�@v����m͵ؗ���u� ���l|�2j����b>��������ۧjF��"�����y�Ј�UaE!�����S�ҍŞJ�o��+��P9�s���1J��p��G�v��sp����r¯}nu"�܀&�Dkt3�P����e��ń��;�o��kW<l�q��h1N�Yӄ;�3^/�^J�Śv2K������r�%@�����q���sܝ�X+]��N;�SC���L#�1�<��%)n� ��ԗr	�'D�^u�1w���诂c�u3I�S\�Q�́<����j�P2���ߒ���Z	p�%>1�&h��[�2a\� ұ�Wϛ��`���P�=?��)&�lo�A3W9�ȅ3ܫ*��4;���%�M��Y�^�x�g��՘J\l�3�$?��8{qI�'�D�����w������ɶ=�: _K������(h[��H(&�*�＿vH_�c�2�'��8;�X�� k��HO`�Z� �!�k����r%v��eF�[���T�#O�Ai�3�ΤO�
��{���$���*�{�1X_���#�ٺz+�sY�d5pMW5ʫ[���yp߇|���.�豘<㺷	�}�����fFu�q�~�bjV[(e��8��<�Y���w"���bxPez#����<N�P9��R*tRO���gc��^ �Dp�(�ޘߚ��,���qb�y{9���x�����϶Y��IK4����,A�\��x���QE9��6�qk�8w��ŵ˹}^?��5C�cO�ڮ��7�c9\���Qs���D"��s����}R��ԬB"�&f&���%���h�q��N�>��O��k� ���Q~���m��e�uR�);�ó~��^L��]U��ч�nM��T�O�%�e���"T�w�l��an	�@��}�-�+=Rr��D��Ŏ���
���2K��[��a����ཏ1vO;�6 �d�SG�<�2�*`�����_��A^x�dL�Cx�! e.�H}c����M�'�fZ�( ���R�z��Nn�{��=򔛈(�;��z+m���,��w���C�C[�W>�.�ojUT�"{'���|���P	��>�	s�[���.i������2��m��Ϭ|0��A��=lč""j�
I��RA������Z�ò:J��9%r���L�=�L؉R�e��&G���(j�C�}(%���X��+2�/�q\��}��#,��hڮU��j�7���el�"���oJՠ��vZ1�/��O]�9�>�כ6�+)���Y�c��<v3uی>�mU��\�߰���l��S��mω�I�/����~G�T�3�	S���9��	��2Z����5�MAV��A����#��2Z�
'.N��vC��8.3���e�kŁ;����e�ՂUa������s�s�:uaB8�\%%��*���ū�ϼ#�1�P�L��1;����UV��X�r�K����:�!�^n�oA�Q���C����]q�o�!�����{�Ɋ���\1�-�U�cIװ�
6��u���j���,�hU�����B�����TjnP
 -y�а7�V�jDh�H52��Q>w��f&��<�5���wv�����^�l$��&6�nYܯO2��>�;�^���ߏ��Dh��/T��]뮯��	������-�y���VJ��*���%	h�h�� x�u����봕��o��X���Չ�p-�F���M?�x��L2�@%޷��Sf��Y���������c}ͮ��!��u���������Z�Kzq�ۙ Ȟ�&��b���۵K+bg�� �$9�ʩA�=L��+�;۝�����A��Þ����?L?P?��,���/�oߞ^E����՗T�2��%����h]�h�B���UQ�%l��N��@e�[�Ğ���׋���^��u�ū��@-c���ݧ�).
�@i7�?ng�ؔ��mF�Z�V��i8�BXZ���4��.t�W�r+S���	��yKՠs�����q*��e#���c��NN����鮝�3 1��0F�Q=ۮ!����g�������z1'eI�A��@�F�f��H3��n���<�@>k�	�	�n��2-�7	�74��"�gߍ��&P�5���RQ�	�hX���ú��%�M|��;�T$m�E�\�_���#�O`]�?W�X�sk+����#:��o�_�:�М%�!�y��ZA64�R�?4S(�R�ܪ3q�&@G�5����*Ͼ��y�H��g�!o�%~��4�		�=�ܼ�C�����h�N	(�o�se_�Ҥa#�4���h���k=i:�3�ԜS��q�a�*�9�0�j9�6��{P6p��v��01��9t������j}�y���o�d"_��>��b)�%h�ҽO�x�wā$�����-���S��V)f���͈K��p�7�8UhX���I7��K[�{ 9pL
�"�H ����1�|��xR������=2���
_|�ہ�3#ʍ�����$C<�(I���Uӕ �
�:�%��J�@���
I2uw,�h,7���ſ�-I#� �X#��fR ������Դ���5��*Q��_��q�DFbc�A{|j�QQ��-m�`MBR��9?:�w��Gυ���O���^YCl��%|M�p�}���ͪU��,�;�Uv^%���j�vu�/X�(�(�=5�3M4$1�eA9 �C�:���yF�Ү�"��`����e"f$}���j̠0��S�g}	jg�u�$x^~ka����a_��Y�`�ʰ�@��R�H���e��lN��`��`�D�4?� ���K��B� Kk�5�M�.R�F�(L�=@�F`��3+�6Re�ԓH�x�:?��'�upw'n��=����Sc�
�-�ڨ��I�X��/OO=�]�)��J��eMR܎̀"�;��o�D��T��=�y���0�FmkrQ8}�`P� ��ջǌ7;�]9����͈οd�$n7:��E��ˈ NR�)��GMf����uI�"�i��gl����'^��$������@�L@�A<)2�5x8�R/>������k�ڋV#�ϲt�0��\I�Ω3�MF#4J�;����ċ�`*� ue"�|��Ht� n���+n�Wu� :^jW��J�`���Z&���9�v:�P�����fH���{@���ޭmlw���{M���x���(��A�J��xfM��,��Ei}b'	�{�&�#좺��������l6fx���~�&hQ���/,���� S�q*
3�;�w�ŋ�	{�`�Ҳ�#�ec!w,q�������:;�Wv�E��ta�t�:�Vl�yV�4��i!�2Zh�S.�ǝ��+����S�:�5�ִ�����7��W����,˷Yj0���8�)�`aQ+���}��'
�d��O���
�<���-WO��4�o�#P�o��� P8�̺��y iq
GT��L�*��|:dvrc��T?Ԓ�_�;�*.��=\;����������[�{��>���(�*���uxIx�E�D0����ŝ�l4$E.	A�ā���g�\_���#�1!7���.�?+��9�vL���XHH�d~]����wd�㙞^����x�F#��c�蓙	�K��F�TQP��5���U�;M��i����Q�(M��~�?Mf3�
��6]��zW��z׭qJ���SX���L�o���x�d��K�a_X���_F��_0!�io�/�-��%�iÚ�.�����7O4�s��z��HtՍ؀���	 -�@u�W�2��ܐ\�%�rƵTP��:''Q?`B��R"��-n՝gP�	�puO@ı'w�N��qe�T��r�E����T��(p�yo���sp�˨l�a�Kt�V��D/�Y����^�HEGr:$�
���	�OǭGY (�n��0���G2�#�;}S����"9�H����4��<E��G+���V���Km,7�R�)��VO�k89��q�Q�\�j��
ߏ�:��g쪆��5�C�6���%�pL���$�|@��x�7����"J̙�f��Ѡ���tm��>�`�$X�^�N�2�� ǆX� �t����q� ���܄�~�|#T��P:���[Q��*�B\��r����l���R��y�����m1',�x��!I<�#ٛ�TQ*���{��M}��J�լ�+�LA��E@[l����X3R��B�5��+4�D��lSˍ�/�b�g,@'Oн��N{H
ҙ1���>r�M}��L�Z,E_H6yԄ�5�Ps}�16���*R$<�<��иv������������.�O�8ګ��b/%�.k#���
��p�@)$������@m.Iw��7zN�:1Ԃ�N�o{�\ �Bȵ��%'I&�������hP���R|��a��Ȩ  �K�T|d�D9	��S�8�����r����˧�F/�Q�)sgtL~��+���J��!� %�-P�.����* g3WE{�Љ��I�s,����M%�r���5��n�J�W���Mt��P�(�HS� �~�U�8�h����X���푠��j櫓��)lq�S��
 �r`A�_���d���&#�y�sFѰJ�p������E}��(��i*�vU�({�SI�����^n�$�Td|\9]�H���|D*�ro�8��q�yݲ/�`Kx��W~��F�͂�(��1`;	8�g��^&>���F��z�K�Gk��e��!	�B�L~�V�]���&v5 �A�31?A�����>B\��r�� �u�+N�HJ�8�d��vK.ztl�̺\|�뢶eь�P�O�1�6t60a@�+��.�л���@b��Z������2�l ;�81����J�ւ@�4L��㴘a`F����,�C���d��u�[N�7�.�(u���Kg�-(ծ�$�b\�F�(9��dr���Tt�/�iX;A�>%�c���~���Aj������ �9*<�ZɆ��4o��Ej�g38 ���4q�%�,�?�7��;�뮐P9������*�&֩ �[���e%"��KF���U]��h���ѳ�������(ٮBG��b�p���h-��s��ZF��Ʒ����'�U�����
�5j	~��tkV��c�j<���%�$�$��R�r`�PQa-�,m߲R����R�6\2��(���%�T?��A��54��<� ��o�<����@�IZzF;�brN���9\���Գ�i�����_h{)�H@��p�yf�>y����c}M�?��$�!��kG��\t��gw$��Z� �kP�u��ʓ��jyˎ	�*�>���+����e�"��R��h�T����=l"�����5����M��uo���IOҸ	_)�B:RA[�/L��!M�(9���w��JX�[����Tv�~2����@�|����"�:t�%���=��PF�+�m�;.ܟ���&4�u�{���0CW�09{ ��±~�r�}j;u��M@���Y�#��S$"����@�-(�6����y�>=Q�������ݍx�̪�Ddm�C�n&���Z]�=ڝR�"�z�=QuT�R��3�"K](��d5U�z8�?y+b�� G����$�8�^�=��j��וG>�CL�g[e�.3�����@�Go��¡��;�abk�G��'�M�i��[�d�~v��X%.^�K�LDM ����	�YoZ��:yɇ�{nc2����֡H��pE�4a;�x����B O&Ş�?�����x3-��o��'�0N�dQ-�U�-��DzΖ��G� �ḫ�u��zg�0��Uӊ�o�K�4��2��+���˓S�k��bgu�L���-`�y����V�����3ߗ�\o-9��#4.�8����>��T�/���< X�"=v
s�R��)n�_L��'4͔,���4a��^�G	��žr8��~�5T�P������X{�	2�d�s)��+)C�u�q��,X;�;G�8Bch�|�����X�v�4}������1�$�+�Ư�Z`�vW�f�0 ���sڎ���[W�A}��(l�4b?�ŵ�H)��_��5�-�qf;N���)��͠&6�݊R�٫�eScQYK7ʓ��O����_Bn��h*�
���@MKj�}p:J�nk�[��w���H�ֹ�i�t������1]��"�&�~jq���;�"�	T�8��cZq|�rG��J���������A_�.�h���R�-YZ�������sr[Ρ /��7oi�h���QדZ
y�?�5�7d�j������f_W,�;h�{���[�Å*K�hM�E�Y��B�1-�NS�w/6�aNj���,>xC��^�G���q�c � ��������.�iM!8���cY��ʏ! 
|�p��L����������:�q��1��`�\Ǽ���H��X��54NI�I�������ng��Ek�ڇsN�Ƚ�d���i�U���3@lV�r��U��y"la��MX��&V�XMs~�����N�UëN� u�Ubq���(5AB��>E�fE�����>@���̢��G��ͦ>jw/��Gx��+��ܽ��5Lb����l�y�M�T��x�{�����x���|�.���y�N�1-w�0ճ����:�����p3��� T9�%Q�U/�8}귮v0�_�߉ic�h�19�c�au���a����hd�q�~5�D���<'�&���F����G,��Z��"/�ҵ��;�ъGb4�w���pJ~�=��?��sw� � �=�<�}���y�}�Ｌ���)p2c�b`��6s�0U�Gϩj�խ�����.A�`�Z����68���kH,�g�K�`�<�ؚ5yK�F���O���X��lT�Q�:��D���_�?&��G����O�#u�V9^dh���~�X���J�&��f����uQ2k4�5U�ԋU'���QHsr���jY�qUWn�>���J�y4�]�j��g�����1.)<�LYE���J6w#��)��t���5�#utg� H؃�����5[�s�K��?�����@����,�ٞ�g*H��t�ڷ��a��,�H\(�M��|n	�1Q�^��ߚ:ʿg�(rm-1a�:^���������Z���[���o*8�َ�dwÓ:G�$A�r�����qtSPD�#*=�u�;|�ıW�4�4���$hz�2�����T|��?i���޴�k�����ޔLj�����zƷ���?�;��UR�s�$1$
0���;F�&�KE���E<�߭Ⓠ���|}� �~��5Kd�1P�8�9�S?:h���f	&F�����VF���S�r@:�PB��÷��f�NS��kF|D�!�����گ�<�_�, �4�HRz4�<۞`d��H+���E�+$�C�t�o�k����Vq��bb`T.��d����!���{j�)�*)�2�[�+�Pt�5�x/ޙ���8�ȭ�^b2(HO�VHO3�a[u�f�lV�rZhh��>wmVX3ʾ�'������E�R�$��cx�U�By-ro��:��C���@~.�����~k X�Ez��k�A,_�@��ڵ��9T&tt��F�/o�5�*��Y�T��N-3���߱���p�=��>�{&s��9^�&�;v��Kn,��,�a<j��Y�y� ��-��Y��52�	(*Ă�������}s
Z�*�c�t���Nu ������jh�������d$�Yl	ׯ�W㦆f+�y^�.W�U�L���4��6Q!
H��SǬ��5�qC:�����e��E="����w�ـ"s�[����٧�����(z�k��Dp?��}3f��d�3���v;���d7�3�v�H�eO#U0��� !i�zݱ#�V��4��lus�����Ț͟=p��Id$�ё���*5���/*I�(R�q?&��bZ�]��͑�G�U�����I��ַ�;���i'��^����(��}d��)Soe�M@�(���F����J��Z]�ۿ�Y���Q�`�,{�˚��i�����1Ӡ����>_����R�9��A��m�{[�^cQ�}�+d_����6�R��r���}T赒C" sHlO>ļ04�	T�6$r!�u8�h�E���2�u$�����N�P�/Ertz	�eYh�GIg��TQ(�z��LW2�C"gA$2m�P���ZNy��qo�&���xeɀ�`"?����]SA�;�-|��LJ�q�v2{)D ;�	��#Aۃ���.�ӳ�Y�K��`0��@���	�K�m��xسk^��wjZ�E�4��5�Mdy����?O�
c^S�HwSȺ�@�k<�'���<��  �Y�6?9 ����n ]�H�r�����]> ��0� �^��T��̳I��C����9L��K�r�ώ>g�x�$��/;�,w�)>�V�F�5��Q����P>o�:p���Q�v�⨇H���Ü��Pi�=�,�ʭ&)m�+�~��XzM�\��iGU�*�|��� ff��Dd���F*�%��sZ�0x�=(,��B�X�Nt��mfz/L��5c[�!�������d��H:z�P�*n���M�E	�@G�������_��H��^p��Hn�+X	wF��衦�:u�JT���Ā����������\\�1�����E<�&0y����Nv:{U�'i'Roh�;J���ܸ�\	{���x��o�G��G�ìx�����,>ϲ������{��R�7ܲA9�H��Mf�5�r����:��d��-��xNo?N�`����=�c�i�(N��E��$I�L����)���0���/(̄IK����%��B${���3���F����8ځ	��ܴ���s��\��0o>�_�x�O�����|ӓ� ݁.3�5}�2���#�������"2%%���&��U�Yx���'
Ǆ�`�>�6�~n�$�ۅ�(�ʰ�HK���(;~ޤ�'c#T�2��!�Y�X��G�l�I9/�!K���~�{��)���*���	}�(t�p8�Gͧ��"�e��^��G
��T�tSS�|+A���1EW���Iҹ��2d횞�R�����r���O:aۯF{P51M��a�Gk/ʩ�<v���4T{><x"�_b�����'J¹ۮ�m߉��JT�=�G?�ז�%��q���I&�!�OH�w�?n�LĳYX��)���H�!��qâ��)�����(ì'J�9�M�!;�M/�૤:tmg��*I\'���ϰ������.�����'�$|r�z�l9��_#��g�Y
44�\w�����N4wR�E��KeR�E$3[������j��Nw\�0q������Igd���\��v
b���-:T�:d%
mު���Pc��*���駤d'���p��$�,z�E {��E	�� ���;ݮu�+�/os��m���K��^L\	q�U,�����֞z=��9ޥ�X��ҏ������ ��Zg�?��}�7�H��?l��8U99�0O���q�c��@ ���	[��y��%���8dr[K�g� S�4j�AQ��n�sܵ!�h�&m�M�Γ�"ܐ-;���l���{y@�#	�����Pm6���T��,��b����c��F2�7�`�I+�9
�,)���Vp_���q�7�AK���g��&ٓ,@L�"��o�!Kl�@{{&U�[r#jxӠ���IHl�4Y�K6@���0��
�'�3]Mh��_m�j�;�^����l�v7��r�>dc�-)�&%���ꏧYW-�!�F�ԃ(7�Zv2���M�%�좢�U�Y�65���D���v"�w���3^��VOw�;qc)��	6�#�ǐ�*5cPf�{��qH/[�^�-���F`լ_�R"�:��,+������ 5��7~&^�`�P��S���T���\�$��E�p��ˀ{I�HN��r#�$��=��'w�	���%JN��E����~^��L�8�KfF�g��h�	����1�$�9�P��7��%	ӼQ$m�ߖ7�:�-��������  54��GC+m<�_{^�a�ɧ�q0�p8��_����Qs�~v-V��
�ا�[��d\"�Z}��콆���ܥ/��?Wi��j�>!1c^Ƃ�*�������0�V���q4�׹m�I�B�wƱo��#jt�u���Aa�#�[Tzi�gb�dR�~⾀�(�/$?��=�
 W������4]�)�ϗGE3��� G^�t�N���?�g�k�ځ'�C�����訛W������V�{[�;�lW:a~�[m��͸K;���9}ؕ�[�E�=C��TÆ��1kzd�����`�8�n/��{'�Xp�#����,�]�e�x@{�]̢v0.�k�9�I��4ƥ�[%E~��z*��ә��ܑ8e�ӗ�]��t���ܟhK��$^/!`Kf�j����d=YT"(D(ۿ��q��C��2���!���8/G��D�	�vv��'$܊z��F�Dj0�A4��%GJ�ȓ��,�i�j�R��;�!��,�bsN$sY�^T<�p�g����ĭ���{E����qx���h�ʏ
=V#ɽiBt�X�ҍo���.yd�[����ִ]������3Ev�ד"&ST�ǜ��q�\����JZko�I�g0M��'��z�̰��1��Eո��t��̏�H�� ��҃w��gƛj6&�U��{�d5g�s?���IU����zs�Y� �rZ�>
�zt<�����y��9xu��6�duf3� ൣye`�vXiߔ�	��Zx�Bl�"r�'x��ޑ��P���s��n))���-��#rwMYnN���Eʘuon�qW�[�`��$D���a���BQ�2a7%�چ�幀��74�Q�m��⼱5�9���d���l�d���N�����B%V$&z�ɋb�X���$�5"9O9u�S�),#��v�E�j��H�S��ۊd��FL�5���?d��[A�C0��ǽ;��7+�h|U������-�Of�X��^Y���r���
��:�l�&+��3N�	ݲ=�XC�2��od�2!��ư_��:�%%/�VӁ$ق��$ذ����L �����c*��ob��xX`?����~��r������
l��։��c��2���H��a�e� �╗����y�&�2�]�c��=�?s,�ڶ��)��2�i����j���w[X���{�r5��=��<�����,����Zo�t(�-Ly��|�?�1i��h��;J
	�FVm�
�,v>+��w�Uܴ {����D̖��w����v����r������fP�����K�^�g㏎�ex����Gs�>��u�-3�tD �R=���|�]_��p{f?��.�`�@԰l�Wq�������8��.�|P��S�r�k͓�3#S��Uc���Ib�q������s��hFg�cN��Ԛ5�63\�%,��pC�g�
ƫp�pW�攋�����J�Z[O
|�/�d|�'K��^��jyL���ӈ�p'����Ƙ�/��hҗ����e����ć��r@	Ź+���a&`���I����*v������H�s��0������s�w6r�n��J3كj�W�L�
�Mi �u�H,/��T�u"�a��2�1�C[<���5�iy�2?�!̤��֞P���w4/?K����pE�H��h.w��q�b@ì�	�Z?�c��n�i�?Z�%�HA���i)�7�n���7oˏi\ޣ{a�wQN@�~0e�aƨY���7�o����'��� ����+��Y�����C:x�Z�N `Qd9&��,C�xxxr�*v_]�Dڬ�'f���x�l���/����`�'�R��'|E�4�"}�ݜ�rE0r�ʌ�mg$hA�{V�-�¨w�K�si�P�<?�����l�)S_篊�X�ؒ�ņ�iҪ�'A�9w�%�M�f��{9y�mq0���#;k�$\��v�{Vp���@�`,M�tf�W��L�~���?t�-�=É�i"�ϵ�Ԃ~��z�/�+�G��"�H��R�"^��E��?�R��.�D+�*v?�%YqX.���u3Ry�$���Lq�Zq��PH��r�>�v�4�n���x���Dxc�u�ⶆT��t,c{��&�������VN ����y�0m�����@}
^�7CH�a��-�RD6ƕ�I��>�	�.��TC~�a6��Zi1�QG�m���؊}|��od��Q��Z����7@�/�����|�$X�wU�F;,I}�(��E��Ji^8�oARG�ڐ!�t�Z.���\���|�H�`���%��������V(�M��Q��f���M�(r':>�$P���$g���LĬ8�^�_��d�����i&�[��ґ��l��� �r(�u��9%!��у�f
�M}w蹙���OC�S�ԑv�Ê# �CQլ8R A��b'��EH�<�c�.FȽ�y�)ɬz!QE�{�2C-|���!b#�?��S���$GD%6���Ee	�O-5zTIHv��u[c���4z��o�G]�=�?���O���zF:|E4ɥ�V���h2خGa^V��*�T<}$�F����݊�I\��v#7��9�����~djg������2L�C�lc�@����g�L��T��~�@h0������Z�MS���	�b"�
^`D�z�;Λp×O,-K$�D<h��X���N��0&�J���S�n���w���t����}�q�z�����Z��d�e�d�ͫ�aa��@�*۵��9����.*�/<���+t�W'H �ୡG�V����r��~�,-�K4�iEi� �[�����I�H�̞��lP7C>^����9�u�n��s58��F/t�S�f�.�Bb�n�~�IO��1� �#�o�A/���B�S���tB<4;���ڰ�<�']�?Q�l%���.k,�x�+��}����Oc�H��8��.�|�8�Щ}M(��S��ֹ���bW��]w ףY��1�����Ful���w���d����t��O-t�f��*-�G4i�������Q�f�d^F���9vOe�
~�-2w�R�����G�X�ǚ�F�Z��QZ�o�ۚ���~�u%�>k�%�X0R�E��0�Д,��#4\`Q�9j��vv@Y��֊�D��2\et</$S풪���� ̜`tA`.��Vt��T1������[^>�]2?n����%�A/{�i����UZ4 �~��	c��l�wo}��aW.p��17����p�<�$P���P�*`cUد&y�Ы���]P�p���[���¥�Eq>CX�h���k���n, :��*��	6_��&�;qXu����ʰ�|�[Oql��o0�P1�x�N���8�4�M��?�kj�$H*��,5x%��	kv�?����ֳ�����eBg�6��6빃B��5�!��Wa9�z���ܠ�0҆��'i����c#M��z_#�Uκ��X�N��e�jY�/f������ڣ��5����}�QŶ�-x�Dn]�W���U��{��,l@4=���^\aDe�7��j~����3%���c����~����)�1 w�Vm]����H���i��T��/�3�b��9�IH�*�"5t=,@��LxQ�,�I���x�R3�>�e�e��(&m��傀y��ͬ&��0�-�@�D����p�����l��;��@�I�w�������z7���[*��5l�ʁ�_{�Z)�Nb����T��=�*��%������d׼m��ǋԭ�Z���Ɉ���S��<-}
�c��v�JnT[���_�N�_�Ut����P��G3�sC�*J�v��)�
y�/�������X��L������N�@q����u�! ����u�h�ӗIJ�$���W�(�ۗ����'L�~�>Z�b̍����0�.��:��W�Y�� Cq�G�^�|��7dH�qk�\���J{����bN��(�ϤJ��d~S���~�^��s�5>����x�N-4��5��9� I*h��~c(��������/g� 4c�7Ԗ�uNXs�]�!�`��J�TF�&���@eI��r�U�c5�,��?e���n�t·:���� p@�e0�d.��a/�rqT��HS(����)��B /�,�w^Ujܣ�h��I><�C)���иa��c��02`�`9�a-�c*=���#̱�o+R����)�^�?U��~3�U���ؒG��Q�P3f���_�?�5�� ��"��˲��xi1��tFl�/<:�:?. ��O��*�����	��@�F�����ly'�Mc�e�1Źn���t���k	��
O<�F�..2��32KjYZw�8no�!�R{eJ~~�Uo&�)��'�@,�����i<9A�X�7�ٌ�Z�l��>�LYwOש	%5���Y���|��B@& �$���j����R�~ҷp���6�5�����T"��lE�D���5|Ms��t����'�k�{���r����^rR�� 2�Q�.��4׫`F�#���<F�,��_��AD�X�G8����<)B6�X��3�E��sX�ĀM즔^�A����Yv���M�o�C\$�3F��Zl�<m�Ȟ~B�d��*I#J�%"��I>��v`��/? ��U���ގ�*CMzC�G0�"^użi,p�;LR��i?���%+����,"i��l��;K��#[��I*,�ol���f�C�r�OfZىŇm�-���'������z&ɖUxe�T�@�A�OP=�[���9���>$O�ޓ,��}�M�s�\%�I��F�M�Z�he�šf�,���]�nA��9P���l�pZ�\��>���Ks��<�@�>��[L�)�8&ՠ�-�M��K�����^�� "���
V�{��'����L��ͫ�"��R�j�0X)/_Z�y�
��J��R�:��m�AH���S	L���2B�)j[�iD!��rآ�$R�uD2�����V���kyZ�`�`���w�׹�#��9p���`�[Gnb3k]t�u#�[�f v�_ч���)m "���6�nj�?Êܱ�ޚ(1S��g�n+բ�._�NX����s��[	5��#ng6��������{ �+-=���UwL�^�@��NI����j�9II�G�����;׳=nV9s��ْ\۹��'oOH����J�[	J�!��r����
�� sO=D#8�+M4��W��JK�\}h���d��W���Iv��jk/�Z���wy!`�>�E�#w�N	fmrN�M�Q�I�)
�_~�o��,cW�VtDQ�G$4\���IoKZa�Y�u1���_BRB�������kt{	w=#�C%�˵��Zom.?����KCZ��~|#�r���H��4Z�Ớ�V�1��k8`[v���T�.��U�K�1sU���ޠ�MDo��ۯ���mVf��c�jb��2�*aCOT+XO&����'��/Dk�ꎑ�
�،�a�P�K$�M�0h]$8��J�� �Z�uR��q�����:�����;�lyD7��5�w�l��_�r3Y+��W�$�ͣ5Õ4�T@[%��M���o�W���:�>q��A>�KK�.�=�ۓ_u�('��_Ҹ���~oƭ���,����SKE��,_F2��N�4� D��c���Ec�Y�(�L�ҩ�k�_~��}5�CjYf⢳m3&J����}C�r�H�:�8��ᗪL$D��5�=��>�%Fn-N*@��~( x�-&IOUS%����\�zT������,�H��ꥮ�{����U΂_�8�4lY�X�ED8��-�9O�9|�ߴD�i� d��F0����p/�)���L2�SxF��)����̕
O�0���1D�s��bQ@!K �;MIt=�essS���m�Y�?��6�L��������(U�A�vr5Ҙ{E/���5���5�U$���0ԋՑT8#�����L<ͫ������i�v]%=fT\�/��R���-`ak���Ƴ��Ň�+��Y�ϏbvY�q:��^�/&�����R�^ɗ���܂��)��yf��β�"p��,�)fs����߲�0�E��1��K��+"�,�w��Δ�~ ��&���0Ul�Y�DקS�_�7o'�_���������|�j�a<�9L�w�ME�}Y)�b9�[�T�DcZ`;��0���2b����8�u��-d}��s��^�0����>��0�6�۫�G$��#5s�cE����������#=Ώ�j��t��b����6� b���2�@U��c�5�i�|��p�ė\N�uk� ��V�����oq� ����6~w��V�������*�5
�.3�m�z�y��N��������ז�����I�wz⢻�?�\�
牭JVwFH7Jb݉�s�Ի������7�%׌4�|�(��6��<�|_�@)�pE� �� �W�M���x��_�Q����
��f����ɡ���u٦����3��;m��!}e�k���c��]�D��VA�ӡ�}�,E+���Z���2�Obz�js���5�[&M�<�+�8.�9b|�Va��ӆ����ȲB��Ǧ;�P���Dc��Lq�I�}�C����x��۔���Jg��S������3'�?/��/�f��$hJ���w�ʀ�#�q����Eq��)DЈ^������U!��7��2�D����0E�>�u�AZ 8+��o�����z��K��x��Y�{d,�$`4�[��#���NA�h��q4�v<�����}����H��!�����,�nB��=9�o��*2��e4�)j�噣��ꎸ�a���]Q[�PJz�kO��5!S��7 �jc��ysy�3boOc��C�IT��q�mEw[2�D��������Bk]��-j7yW!��N�����c�,�����ꤦ=X�I�Ĝ|`�o����j��m�A�	�4:HnH�c�
Q�艁��<�Dq֜�}�� �e&
%E�/��|C��"d���I�ĳ�z�)X�2����1�d��"�[����E��EXw�����<J�c�`���59<���c?_H�.�Z��RSK�ɕ@�;?��0, �̉�9�Nɜ�����=&��!�"y�8xbN��Dby���x������Y�!'u�No/a�Bҹ�A��9��Hg�3.0r�.��Z�U�/���R��xU���s ���'�^ �ݵ��ղ����#��g���]�k�$$��m���9!m9�?"��Pep��0����;E���q̩�6'�^�8=H�5��J�M6d��Xo@�|��.��'�~��zP@}uC�����sڍ��'\2��W��I�'ĵ����@�t9�?���&.>Ϭ^����az�'#Tjl�Ã�I����+����k��	c��RϘ//+k����JZv��_���' ��(Z�fc���F;�`��{�%w���2Ŷ���_;w�%�ip enP|7��$�ԕԔ��*
�����_a�?t�����<�#s_��m%=D_�~�z�L�낖C���J��b�Rf�3�3����y�$���bK�kY����f�@v2�KJ��u��ɜ�g��ˋw��j9�X�}���|�.,�$�-(98Z���7w��E�9��K�3��8�5�N,[|ܪ]���d������h�8s�|�p72�]��T�����y]_�X�>��n9�B���:>F�鵜��ǈK���7��\�\<	�q�
�[sxO��=J�d�� �8t"j��u8��p\9�Up	U><nLZM�K�HӒ�N�`�ь����8#w�"�(�?�S�CF�l�w]���5��?��osQ���4.uiq�$v���z�A�Ά۴�sg}�]ÔU8���M�?}�k����m���{�k���nn"�I���oĝ��k.��,�l`EBaSK����$��lN���W��N�1�A���O�ͻs2�m�}7jU��5!m@�=^3�@)Gs,i�$ :쐦���c�ѳ{��$�����a`�k��5i^�z��+o~���3��A��K$>
�)�K���l�\���yg�|o��^bʾ�`v�/���"��6<�W�_��N�;t�Ri��xD�K.�@+�o���s)F6�OY�aj�Z�?6Vʎ6�Zbh!���;�kd�P�j;�H�`(]�[��n�Se���~�����S��:{m���!��2���-f��ݠ�>x�Lt:�Aw7����^�G������1�D_���ߑ�Y��ЊN9%v�+�Vk����c|]�QZ=�c�۾U���p�.�a��H�D�H���:��mlz��fT�B�`kf�-A�e�Y���]�������u�L:kB��陎��<Ć��Mh�#k�([���0H��pv�s�R�FC"��})� �a��?J���b_�+P\���YyS�6D��-�����K
��WP~��G�Ib�2_�HZ����$�&�$�h�A�áe�
!����ފH|b�z��S�:wPo�n�w"�����o�y�t+[�P���~=ȯ-�A��w�Q�g��o��������=�f2A��o���LR#Ĩ�W��PL��B��A�O���]q����/�L�������ۢ
+���SE6�������2�i��Ai��Ɉ���;s�H�Fp�)���T.C��P@�j�x����[|�X�TKUK1�'�*�����/S�Qat��MO�Ξ��ĩ�NpxZ�����rG��cjt�c��k��5?9�����
6e�[8�BG��j���^�ȵ�����b��=�8uzy�������ghX��v��%��i�T�SG6�ҷ�H�>�h����=��̮����*S���&�duW�qF��v>졣���h��Fr�!��0��I���]Ղ�al���֦�ëtW@TGE��0
G(� ��*����~v��"�·\�Ҟ>��>�y�����. z� {���2�Q�E��Y��x5cF����J�=h�K��d�R�_�췼�XOAS`�#��Z���ϝX�(�Ӳ���=1׍�@���J}��_�~������
�؉j��p��zD7&�ԓ��Ďn[����^XU��=ʼ�<L4x�G�~9v����ڭ��+�2����o��f��s6<���|�+S�||:^���k����(@y6��j�*����T	%�����؊����\<���KO�أ.�rb⢖�I���Fh��I-���I�5��~�V�h�#9���p����5�FM�B�a����ΈEJ�yh�{J�>��aQɅ�nf��\��
ͿU�E�R[о�-R	�\?$QyV�Cj�lmtxO%T�5�M�:~��\����	G���R@��%�J��N����q~������b�i�H�z�8kٖ��.�]�z�#��Yx���AnR��
|�b�����)JlƐ�dKR̥��:C� u0JA�Ũ(@�]MP��BkMC�����0�p/*9��v�K����+�*d VG*�e�=�Ƶk2�^����Mm� 	aϏͿY��u��x��6�z�0-t�"ͯ�����(�wA�	��@	�t\�>���%yy^��D�7�+��e&%8��6&;.;,7�՝w+��RW�EwCv�њs��zH�7l8���!�Ce��d�X�y�3<ܼ�OF��q��'j��5�i�Π,�s�&h�^�j�N�w�uG%J����Ԧ�$�eL�!!��ݰ��8,��Ҡ{4T�����B'�/�J�p��Ntf����F�ko�n�}d�IW{-E���-���J%#�\�!q`o��hҩ�r����/�1��1K)
Y��kHA,�k992��:��E�д���lv�����u���uV��P@7�*�#�eL��~α#a���k��pǏ���#�#E85q���r�b�fc*~����i��Q�ߑ���Ț��M;��y��{0�զL1��(f(�r��+��z�����&	X+D�_����� �B+E�,ϊ�شBEA���8�;����w_�=����xhWm�%�����ȕF"E?�H��.U���d{��\Å
�~!�Vb>1�'��#� ��h�}i
R_�/��EQ���W�m٢V��O:G�u$���@s��f%o�+b;RA���x�zr~��%�֜�� N��P�'Ư��/<}��均���z�|N7�y��@oc�Cc��y�<��e��3�ƈ��X��UR��~R��zP[�$]����.���IeKR;[�]��ڌU��T�&mOUnO�0��K�:e��I��3�6F��K+X� t���w�sH�Rg�^��	e������D+_��+�(�usY
Y�%H�}p��_�IKh�O��z��	��aH�@?���.�zc�2�a��j�F�5��3a@qڨ�W���?g�}������X��v(��ϒ�*y3ٺ���d�h� �sʔh8K�oL��|�8(���<�Q��B𱛏27�6K�/��`�jRh�oc)2�ĸR�a�F�@ٚ�����"��q+%FE~P��U�r�1������W�~R>�<95���o��~�t
������������jL�iH��EojB�;x���P��N��Z
��Q�ԃk�W�� b��9�V�i�}R�����h��k���i4'�T��H���-A�u)	i{(��'&f�Eb�,r�	���o�Sy��	b@=� ���<[�n8�諍�S�

��y%&��?�38��J� t�˹����%����hk�N�@o�K7�j�=� �^6a���l�Bu!/eu:ʝs�F��F1tWa�P%�S�yc�5@�Y�
�I�������N� ��ݝ�uJf��&!UC����wZ�`�#�m�#��������)��_��٪.
` Z��^woG-�� ���R�6}=�ag."�5�.���W���=*`)���[�:��Ҍ�j0����t|�n.��>v��5����p_�bJ`�����v�2���Xsh�/�{[����g�;�c&j�U���&����$���[����Ci���0p�v��=���o8(�o���:� ���	����N���*�}�<��g̀��X���m)f�3�C��W��%�h��s��<����t���C���ґ��n;+ts�q�V]�C�o� p��yY��݁���΀-N��ӿ������#t˛1"6��X��3M`+asdK/�����Q��A�*1�q���Ȑ<�ѽ��'+����K&_4���`�exku������I���ո�_���dl���I�\��j(Z��=n�gEV����c���O�X2�R�q:F��b&�M��H�HLQ4E���F 5]O(���3������{6�D�/7�[R��
1�����(9�'D�f�N��(O�@��~����,�֣�~-�bޥ�%��$'�~2u�/�Hr8 ��I���\��%8�u�]�\�y\���s*�=��'�k1.��A1�@ѥ���M ����=�<�yWu/��Of�ϯ�E��'Q��yJ38�Nbmq{V jM�V�k��3\�!�J�7}��S�=Ǐr�LUX�~��p	�
����t��SE ��iz����J����	�,�K߶����N<�	�+�0�
b�4�z��N\m?V�o��K�r������`)l���� �պd���Dhn�@ש�s��^�H�Ȍ��7|_�T��s��E����t;���I��9Do2&m�:^���]'�tX���?y�ǰ	o���rV<�xXR%�(ñ��mY�9
1d?�M\9�����BF;�V��Í���8O��\P� �����7��傞�l�`����u3 ��q-��Z�76b����r%�;����[���X���&]U��.o��
w��l3�I���.�`����1)&.�6褽Gc�2�i^���њ��U�������]
>�)�]�)Z<kfB��~8��֨���#P��˹0��@� ����7��y逆�쮪EIl=D�O�х����Ҥ�w�J�l&�iͭ�!|G۪؇�i�eO���(\e�.�NٺT;e�ǻ���L:1O	s�^�=%!8�u F��e�P�x7f��*��J�5�ܹ��i)��m^������T�Q[a�
*����l��1�3h����+�w�vb�Z�,��aاO��~��ӗ"a�d]�ټ��w@,�����@�_�^""��x�or3
��ߨ*̩����������i��.�4_���������otD��&kj<�͎��3x�J�*ʟE���W�w�G�o	�4�����p���<oAa���ս��cN��������Qv=|�5E�7����u�h�\�]�fK��z��J
�L2r�;�q)u�R�&ۨ��j���N��h���W�����l��߿V3�!�H�.KQo&�Fu��[�XF�!/ǳD&�ڌ$]��oKh�`ܦ�(4�Y��H�Ƥ�A�?-QޔY�����u��/h&Dd9K&���\�3�3��CZ�\ڈ�cq����������'�E�6a�iS�_���(�?@f���]�$�-��������
N���6ѱh�ܣv�IN�ׁ��s�k6��!	sgU�ܴ��b&؏�(h���򖜃�S���m�_�W!$�#�	0���y���Q���6�Ā�5�ᵜ���sZ�ueXh�'k�+�db3�]#���(�I�
	K�פ �y_�cN7׿��_�G�O�T��a�����lQ�n6��EA�F����0�@{����d����c�i��X� �w���W�/0K_L���<��5���@+����ʇ7�5���ދ��䁡&$�im���s���ŌA�8��N�-��k~T�6�c�{:e�`��슀��QYڣ�� �������w������� x`����L~8d��_u5̘2��&�S�@��M�rt�i?	Ku�h�ko�dW������!j�K�d����4�f۽غr8sy�\�**����:E�ꚇ�����禨��$�W(-5ÕF�G�B��Z��t����uwJ�%�x#Ɲt����&�Q�,�N��P�;LR`�9�Y��/w���y�Z��!�H1����J���%�d	�u,z���][.����4fg/V;��$K�gP)!#����0MW��LA��~t*��hC�ӝ-J��4�ȃ�����ݔ� (�0����d����z�u�맿\���^L,�5>0�}��s�1��s����,�Ɛ��&lh�A�ʘ�?e��^�@�e����N�����4�	�a��PF�a�?�̌.�'��Y�2���~�n�(}G (�Tc#�D�����i�\��Yn,�೴B��h6�K���%	!_�� �Ruu�����Ȉ���qi�܁Ds�{�|PXB�R��摉�w���%�"�n�`���CI��$���؛�O'+�`��h���!,��҈tI'�!�l����>){_4;[��ۃ|~z�1*�/�ः�����)Z\��Y?!{��S�R���cV��B��ܚ(�r�.���5���g���q��.{����9��]0S;t*H4�Ank���p5Pt��_�ȑ�m����=ԑy+IS$��MS�M�F�i�wq��y˻o��;e( 
@J4���q*�C���}z�D(~2�[�����$҃�=ˉ������2��g4�Y602��3�Qjr붍��x���5X9��9��D�ֻ�[�]"���3dFNtx�Kߣ&�*<��9�8��� �����Y'Q/-
��O<��i�W���n'(�X�g9��=�!|���v�"�xe���X5yq3o��
���G�����CT|�#R����}���%�����׳D���I�*�4��b|*���*�n v�(}�NqC�J�����.ܪ�j��v
$T�\C+�����eZG��qV=��o�>D}&}�@ȱ�wg�t~N��I1'��l����X��	���8�ąﲑ��~5�@�f�WI�/	����d�yX��Ė#b\��05v�]gїձ��3Y�J�5\����:8N%V���@�[$�f��?�D3R�1�:�^���a���Nyܘ��ߗ��7n���❗{�A�&�ie�n�c6��I�}�����t�x�,�\����6UoD�Y,�R��X�B�j� 5u��T"��题0\���h��M]��K�넲��)��m�Y�RĢ:��<|@� �-�4b��� �S"G�`u2�Yً)	�NUP���#�6����ү�˚p�^I���X��m������
������>޶��pG��u�_����0s����q&硞̰������	��������I�RёwVX9Bܚc�/w;�~C�&Pw�Z�0���SI98��*6/���\�W\"�c���>�_�O����j!��6�������;V�9�L��4.�B��Ϳ?��%���%�;,�����r }�un�ۊ�C��0 ǶG�
��o� �f#�G��E������7���A0�N��z���g�e��B]�6�1�0�O9���'*\qO~Ȑ?����g�s��}��fU�ƨr�F��t��>v�|8�q�k�ͶQM%g�h�{�b�6@
*�;S��İć:��2~��"|}��WAh���.��a_��"kM�YgzP����SZ�	��&��$���~�&o��x�D���p�9�	��t�k.���X���s}r쪤��r����NTV$��c��&���^�X�ސ@.B�| nP�;�KsU?��q-�"��GO��>���̫�x"Y�$~�S8�>�8��8�U��#aa�;t���F��!��'��遽 =��hJ��ַ��^�3���S��I��f��[����h��#d���<�&H/@�_��<�}z>���+�>�]O�sX"7U�To�s�R�'f{3�@չ�j��"�������!����XT�"�G9�X؃d_�� At*�cz|c�,��tUi�����9%�R��kzMnƒ�w�豟��
e�2\E͏0�!���/T�B�Ŵe<N���<�8Dp�(��4�|E�;����^	�����_����/��������������F�~3��>�Z�1��%�0�g"&p�{�o���W�V(������,g��D�W�Ӱ�З�;DÝ�v��FxK\S�a(�)�XvukQa�S�@�˒+1�'G�h�G, �(iS�905�y�{\�c�D�w�X�2����+�y�a�jl��(�E�z*��E*�
���|�#u��*��2�YkIŸ_LfLvtϵ�
�3髩U����lq�r?ןs`��%0ᙴ�F5�I�����`�:F�
<@܅cbj9�i=�m���i"'�<!��ft���%��[�)44f5���K� >-h�Y+)�<�i��|א�+5��sB`Y�ɼ��<�RҠ8�jr-~&��ˀK���/���w�?@Rx3u��jb�0���^|���gs�@�Þ�P��[��b�ޏ���;������y��>��f�����3����m!T�F`+���ץ�$) ǎLB�nG��_����k�x����"���Y�ZG(�MY�^OiG�t����
��Z�!{�irC���2��DQ�y�����̷m�
�,J�,���QP<�+s����cwl�����wA�C{o4ɻ@.����@�9�&���o�ᶻ`��Rj�[ ��d��<�yP�Z8��m���*b��@,LN����5�1����xgƝ���%�b���B�B]詋	�n}�Z�)-��� ?i67ph�DK��
a!�����ϧ~]g��pC1O}!+<��$ɥ_��-���q�/�r#g/J����z��f��n	�(2�!Ⓚ�3%�ݗ�E�D�בּsq���H'�\���w鯰M���b�	#Ñ�qD���Fd���n#�T?A�i)��#v|a=�?[K��פg�
t�&NZ ��e�k�y>C&�n������2Qy�*�@�.+������
�ݟ�`)�D�=a@Џ~�r���e�&���,A���y�$�g�0� ��~�S��ߗ�ƬY/��+���3^(�Ģr���Oݽ"�</�
��c�Bǳ�UUN�肋f
�I��5޴�Y��e+�B 㕙K>3Y��Y��j8��3���qI̻�w���0����$�s�2�'�d���[�Kz��A-�|�n�q�'�4����&�x�r���(�?vi��F��U���b�V:#�;y"��5<��<"g�J��[��Z�c[TJ#���q�v
�~�r��5ڢtD���z��8�R������i!EO;��e�.�ݎ���ơ6;�P�&�9C~���7zs��5�Y��L[�u�����o@ʗ�����b���re��W1rXJEQa*�+dzu�:Ӫ�����%!(��<���܃(Eܹ�&OF�$
Q yy��mG��V��yXҮ��/h�2�Q�^gr7����ً��
�r�0�So\-�����Y�����
��z9��~HM:��A�]����_���AM,��Y�\\^C�e\���)�-��������I\7�d�b<D_	Z�+F�kk�,�V8�؆���/�&-�"%��� 78"�8����]�a�a0���#(hX�77���C\Q���`Y�ȋ���� ��O�V��O��0!;Pb�5�"l_����X�-#�b���W;^���6�,(ݳ�o{+zncEp����<#�UK�]��ظ�!v�Dθ�Tl>���~��
�<��E;���Ѥ>�h̋��. ��x�q�;��ٻ�͂�0�e'�u��l
/�L�����@���������ߍ	
\���y���K��C�ʧ5.C�	p�`{�J6')�BFZ�$��>�F���b�T��	�Zu!cK��������w`R��l�u8�Զ�����7�<��D�)Cw�d}�A)���|r�����\�a���{ޫ��T���`MM�"Z�S�*��M����O}{�L���pz��`�j��QQ؆�����N�Y"2F7��g�0���W��?���C(�^�Zı�f�+���p�ϝ���c�ԾEmۺ��7;h��׸S\ɞ+�ẝ8M]u�Kܝ�M������	)������Њ��6ů}�X#�:d	�x�4+8z;�M����gsޡx숱�����re�2��� w����<��ox�6A*s�������i�V'mz	��~��)g�I��O-�����^����.��C��*�y;r�q>���[f���/"�����.Ņ2o����C��փQ�.�����H��" "���wV]|�*p.�2�WT�PO�����q_��_*�j��!�Ms�}nw���o�}�Y�ܰk���R�愲��L�p	�WG�e{�]��o��EbF��~��*[G"Ay��x��(�����Yox����ܶ�{ctC��D��+��*�w����T M���?�<�4�3w?�A+qÀ�GKOuz��p����	��d�Y&y3���^uwe���f�iN[+�g��oI�[�~�c��\�ދ��O�L�A�E�' $Ж'� ��%�9�A5
*2��0�Y��rKFP�&���5[�s��i7 �D��8W{yyl����|yƠ�X�č��"��D<��T��6f5��a�:�W��%I�X^:>E5�֊<q�Y>P�T���<eA��QGk��H�x����]+������@���MSIc���+������2�~$��(�2ڧ�bYE3	Qu���^Vyu����q`�U��ОJ��a��Dh���d�� ���w��+���(�U�v����g
LDǽ��"�����'M��N�"�Έ�E�}�w*˶|3����ψh{YW�q"�=V[�K�"*E���t������}ܭ7���y��,RJ!�Ι`7S�pL���{d�S=�����d��u�"?����]�i��"�1s��%�Ϸ�~�r��q���L��`[��ԫ��E'8�DZŰpQ�}^�8-�
���3yR�"�_��(�0���jJ=y�#{�����9{3^b��G<��iy�-/���Q�����҇�� �նn� ���lH�\}X
����%g�-��69�[ �	۸/���\�r#�rrO�����7^�QOY������{`�;���?��9��&LMݡ��vPͨD?G9�6$g=�FWI����!�y}c��
� �i9�c��y�&���9����+���}�~�y���2� S���ڈ��o�OH^�]��&�Q�:���g��]����Xd���V�E0�Pl�P6W��1S ځВ��#�My\�F��L`6G�z� Z��)�_j��}^X��=�I7b@}�4F�so���\@��P$wS�UH�&�yU P�� ���7�"" �_�����Zs�Zʗ �T;JNk:��&{��gǼI�ӯ
T��o8H^��_��5q��h���q�Bv�F��:D�WK�4M��J:ږot9d!q�` ��������Jx7�r��Z\>b�a��[�r �'"\|���h�7�JV2����,� Y�-:{e�x�x�P�����/�P��߽g��}���_"D��lU��tV�=:)���w �f������*Ja�C���s�U�V>V[e�8����z'��X����oM�8������z�:�N'8�{1߲S��ʹ�����[cQ���a�mdX�b�,ڦx�:�!]yw�/2��3����?���v�r"�h�6�nX].'���Y��/܇��]b��/�����n�F����7^FH���!�xfj��EX2%�����Ղ��$�b`[�Hp��B��0����FtL�U����:&ڼ&t�傝��`?XUiY�B�XK����S��}2\��b��mO�� ����w�j�P�r��F]8z�9�|[?��?e��а���h�o'7��U-���y̆(Y(����v��*����5[�c�X`�
[y��)軾0MNXP�X:yC��\��J�r�C�l�Fl��\��(�k��J&�����.�0�?ycu`�@�
���?��^���:��N���s@��Z{R���� �m?�h
dR��A¹�
�*���r� h���K�:=p��SWy����(�������5��¼8lI��6��1;9m��t-1���?��L�+�2��=ߦ����o�(y�y�pʟ���D�l�T�z�J�#�bz�hM�q_�����	/�������(_��>�j�0n|�7�$��[����OKL�����U�/�R��Щ���D��p=x��tm������O�5�e��F�z�]QD*jn.�w����p�_�b�q<��퍩���k!�qA��駌�ϙ�E�3d��ի��UC��m���k��4��Z�3h��z��|A��/�PR�ɈJ`a���bb��E���%��RQ6r8W���'�^�"�N������[�m�tSӫ����K�P�X�@I�W*r"���ͦj��#�M6�}�(��f�Aӟ&{2�sI ���:D�)���(;�m?8��7��hjH�=�OkUm���PD]�M�I\�U�N�����u�*��ݖ
�F�@n�CKE�Y�a$$�S0�
_�+�]#���Dsٙ#i�^O��0#������B�ѹ��q��"S&awh��1ތ�~�څ}����oD�A�Aҭ	���;*uӑ+x9F��(����������W�>Fv!�_����K۪I]ĖiѰ��mm�Ә�\
 
��x��^GA��Yr�	�w�_�	/� "1c�r�/��nE�Ѷ5]9��)���SA�j�����>BS@����)���V��Er��D��=�:�ª��-�'�OF��a �����$��?���������V}\]������F+�ի�4�4ZL�,�:�"�) 2�TN��@�y�ʬٚB�3�}g.D܇8�?t�a4���hxH���2Ġ���c�L�]�����΂@vdײi��&�%��F�.��ۼR�i�"�;��<�XMh�d{n9�"��t��V�0E!&�'PC���j��6�OV����t.�0��nB�{��Y�\;Jp�˺#�=��8!#�o��@<0�>]�`�����-�I
q�L�����5�
��J�4�it�����Y�S����h�f��f����L#W�=�wq�u�����	�ypܾ������ۦ(Dx^��H,��ޖa���\�w��Ӑxg�y��wd��������W����c�~��2����rRz�����bC��u`E��Qس\��iRڰ� ��)0�oZU��q�.�
9�O��	�V������"^���ѥ�J�*�_ŕ�m��L�R�gv@2���Q[�㼫�C\��,M��4�dJ��y�<�i���S��!%O���zu�}E_�P��]U9S��S�vO�G�T��c)��_�)�߶��g�e{���-(�]����-{9�'��T(�8�=U��h})_�!?c�@�_͹y�ȏc�uӤM(Y�>��lJ¥2h�^6�5T-xΪ>#�7\��+��14���R��jE��?u���N�똓�j��T�ZnMP\�XXA2�g�?�(�P�*~1d�`7y�3覩W%�_�B����!-�# ��cb�U:�/3j����,�^j~K��AWx�D�L�Eץ7���Z�t ��u�̥V-8�d�L�Pi������4?7�μϑ����]o��XI��TP 6h��HA��hv�w�7x�Au�D2w���>���ӊ1���yC2N�?:��V̕6rjGFG8�|�o.;� �����	�(�ag,�	�~�q�JRh�����1���͊���V;�Pl�:צ�y/��<M-E��;�5eco�=!���������o=� @pm��W�Ŗ�etU�xrrp�iP�Ŀ�E�f�Uβ�g��ВK��~M���W(����AցGX����G2�*<�AZ���֡ߙi����_�'�L�\�+���Y�okC��[�){�(����ժ]�~�����H��ᗠ�ۘ�m���&؀��B_��G6�waIK�^QPWD}ܹv>��P�_�6l=���Zp��ʸ�3�,v�[\_|/�q��51O�!vzZǟ6�o�E���~~X�e��<��t@����g���^d�g0̬)d���%z�z�u�>�ZP]�"M�h�(��a�D�6���Y��k����ӐjZWU>���n��	}�z"Jނ�St �	y�;){���B�d~(�Ԉ�/��@������Cϋ}�:���)��s��m����[�l�uF��
2�8�svn�³j'�Q��?%{	%7Z��}���g���F)kuk��)#Ny'�^�_�o�����J�.�T�U[S��S�i�����L��ѫs�yD�r�ן(�!�ܫY~ұ�n�S��@W�`�+�����^��F!�}���E����syC=yF�/���(��^t�"˺�ʾ����F	������L��+@��X�j�'��8�fݡo:�����j�(b}��WI�s�e)�0�?����<�I{!Ÿh��L�yy��.�O�ހ<��.J9L��u�����ք\K��E�C;l��B��2	�u�^S��\4RhV�����MO	�A�$s���ɾDb}��;��hƚ4�zf�:��G�Z%�)�Z����M����'����t���3���M(D���ӊ�h�Q�[jğ�%����G��gq0�bv�P�!���G}G�x��/%l�Z�=�4&�W1��zbG�<)��u�pK�zF�l��'7:= m�(¯ci����H�Ŭ���Y���KX��#�>�)j��]8�Лx|�!|��*S�����s��yb�H�Fd��Eh(���aM^%����}�`̸-����s/���f��)/�t�ň��HB�SI�L���𧼵}Wq�1X��������0�]I�9�-��>m�I+>�4�sp�6{�,���8�����=
���������+=oH�~�O�1�$�^7O2�����!&c.질���#�j_L3:Й�[Q�P���d����S�U�;����`��e--S��T�ϊ?���.��O%g��@h!PU��j�5^��̸�"%|�^?�P�Ap lթ~1Q�+-w��_@��:\J���ǲg�#`�xi�q{��(��v�=��f6�yd��O�q�X����� r�T�T$�yN��q�5�mS����ۑy��W�LvaR��P�ǈ2���O>�g-����<����y�XO+YG��P���0�n�@SR�����X�US��s���8�;��Wi	�3[xl�X�7>�+�,�&���q:�Ķ���X#C�&eW�:�&�\iՌw�R�7Lې�.c�n��v�2�	�PY�V[C)��-��C�}�D���m|⎎��q�4����Gh� ����DؙL�o��t�q�)�/%|K�b<�Q�}�ެ�mA饄�L�#]0�MK'���G��'2,%+d}R�]B{t	C�>,@�˯{�ࢧi�J��F���V̷���Q�(�s��e:x��aЁ�D��m�d�G�f>��5){	�<f��Α���>P2+"������DIo���@�>HE�#�!j��5����Ζ�����2I��(��XнW�ZPEZn��\z�
�l�|�8��8
�Z�c�Z��d8?�D�؉� ކ����{�ݚ`��DB��ǽF�/��֫��|{����\��7����P�i��F� ?Z�W��I�U*�P1l�aS���5,�{�����qv`����^�-��b%�_pT��уq�`�1N�kol%T{� �J�&��Hv��q�M�g���]I�[�C���B�Y`���29S��7ڳ��e�{����r�)}����4��֣����Lms����ӕ���4��J˖#�3D�B�p@�q>q��涘�x˃ ��h��-K$�+ђg��S���ż>����{�f�J�#>���_Ϟ��{mv���=}���ɢ-#�}�� {?��#q�YZ�B5���1�J� #0����l�ܗ��2o^��^�q���jVd�8yf�~���ؖ�l*߲j=zn���)�Є\�.�!Z����%����+" b�K���^�P*[���͔T�z��k�)p.�QC�v�i���e+b��o�CE6t��j�p�j���H�c|��&qj�$��ђ
��9��`�M�b��5�I���pN�*�/z`���^�]�Ǣt�i@��솊{G����� �z��~d�����E�G��d(�az�G��bC�&f����2 ��X�w{T;L�)c�Q�!i�u�p��K.���k���fx٣L�_{a-��ڲ.	�<gY_^�y�t�p�v�M8}ﬕ7��? ��i���x~	ˀ1lzPpfN�� �Ȗ�҄q�Vd2��N���F��L�o-s3��k\��1���_0�a�8���q�p <~�W�L3���`�y ~�}F�q�P��g�i�.��k���a����t�� �6-���5
-B��&��ߐ�b������T������: U ҏ~�'���=�S*���M���Q�C�jgƐt����mc��g�YՉ؄����b
���zL�%0��G�Ŋ0��E��=�`>Z���MU��9�Ӎ�ӢN��OPv�n��a�zM�����1j�K���y�:�@��hQ*��C �`ý��HN,��ǁ����_!��U���Ul��Ŵe�v�V�F~5�fz�ﱠf^�E����8�P�~�� .�F�lھ2���ܬ+K�TΉ�1�|����l��èQ����>��4f���)fk�-�y��7^ב��Y�6;w�S�q��?�J�9���̱
�9I��� ����$���¬o х�� ˆ��\)��>����ɘ��s*!H��iaʬe����Yö�#f��"��i�:6w���*�t�b�k` ��%�b�[x���?^�?k��i��;�� a�@�l�9���7�_	�T��p�6t��	7T����!K\D@A5qC@֠-�7���O;
,V
c�`{��L�P��E/>�]U�U��.�*��'~��0��ѐp�5=�8��y��n���R�Ib�/b`	��9������I��a����kG�Ѿ� �X���ЄL��訵S�����͖��n�>_�S(��/{�ɮ:x&��˝��!��.�
rЏ�Z�r�;O��M���c��J��/�s��*��tx.�.
����a�H�Qf攃��n�cP�V��XODK P����1m7�����0' &�����[x��@�Ԡ^�X�N�w�[4�u<����?��=�j�`�|S���|���r]"�G9���':	BP�#�MiH�vSroj)$m����������i!EQ]�i�P ����g�!��y�<z�:RSJݾ<h̓������������=�@'Ih�G:�J{�!��ы���
 s4=�T��Bl�$~]*7@�X\���i�G�>I$��0�h����"���~�����������_�[b ��j��:�Œt���X(��n�by�v%���������;zY�5��:|�gil|����.�q�J_��)"�겘� �ٱ轕��"����z���S��l�B�zH=).�[�,�j��h)R��~�m�\va�p@�.��F�.�3
���-N�_��P��	�����Q�i���ɨ��i�n��	�3H�X#~��yF6�	��q�s�I�[IX�it�e\I˲Tiv�)8<��V4���4毬�x�g��&,B�ϡE�o��v�dH��HN�.�݂�Y⧥@W���4J�U�gp��	����j�IZ�J���U�T��Z�.��\�҃7������_��f�iޟq�S����(�������z�(�3\��`��I)���$�Y+���ü"�P��z^j��1����(k-X�V!q�C�w���ߚ!�����ڧG�Q]nL�ֱ��i�K���� �S��*����+�]�hу����;{x;r��6�Iҟ3�<��?�2�����^K�_��pz_�f��kA ���,���o���`<������WF2�<D�}���r�w^	� �.Cǜ֠����E5�tqЄ�ʹv��s|����6^l�7��8R?Grc���	�D~��g"�
F�]�irU8]��'��!�ލ0b�h�z�9�����Mg7q�˺����5��N���'��ep_$jvS������迍Fd渃�D�i'5�{2��Ive����2^��>{v@iϣ;[�y�1�)Hcc0k�li� �mdS��2�W�?�=����pK4',cl��ks@�O����
f���F��xk$;蔽VY=��89,��%�U�w��-K,d!�@I�tȟ�Q�@<�~<�����:ԉM�T�߱��@���\g��%�t��*#_�C����!���FM�B���
�2{�v
�Ad���&����E�4��JxO��*�+�����e S'��lM�/J�����o8G0�W虽Z��6�Jk����sߑ��M5�E�g�ʩ0��Џ�1��7��B�3~�5���g�Fp�b�u� 	���� {�3�'��hu���炉n	ox���|�dj]��<����(#ߚX���K��Jx�ӿ�ūf�}�xKr5�=;�|ds�I�NM��-d�]�(�6m6��x0��x��]S_8�{M�ꉿC�1N�v2"�]�\��(U�BX��n���)�Ln��D$y���<�u����&W8L{�����&��u|��ݘ$��Ĝ��U�����Z��揆�@��Pb�c���';6���X^Qª�/S b2�׀��.�$�j5��~J]U��/�sZey߶`	)k�;��I!w�˗��n�萱�%ӰZD��w�_�D�$8� ��xl�3m�/f"�խ2�y�F3zUN��s^�!�Τ0'}�c\�k��6~�˦�FbM��Ĭ>��w������u߫���h�bb��i�J{��u[�;�R���Ҭ��o��}�	�E~�)v�d	-OD2w��@q8+��0S�L������B�QGڃ��.��Y>n@�2�vW��6�h�|��b�d���T�
�Q!��nj{�qrQ��	G���A�������7�����0��
���*ک��c-E�z�P�\(-26�@#DH��."�B��#Q�^^*c�BU�����~�E3�Ȑ��O�A�jN^<���0�`5u+`���#� $���d`ly���[�>
����U@�B�-�=y��d;� ب��P!��9s�IWUE���l�<������WbOn#2s�/S���3��~��!L8��]+snDQ�����)�t���X*:�/��DM���{�p�2H�yم�kY�x���RǙ^�?�;,��E �R�=<�p����ԃ` 9~K�t���#���D��P���
K����G�fk�����5r��6�-o���٦٨���
&�5���I�����S�h����{��5�!ׅ�}�PZ��~�f�����h�d�����z�rHy��-jLV���N�-ݾ�cHUI�g׮�B�u�t���u$�ğ�',V$KL��$|�N��>�y�+���P���7ё�>�G���0���t�G�:U����n��i[V+�Y%�L`~��_8n1�b�g#���V5y��y����_:���:r�������X� �)9�-~��fƩ=#m2&�Z��F����1g��T	ïJ�YP�t����R�9v���h^�	���� c�~����E�q�?Xq�����~dO�������h�,�n0����#ΰ:,\W�emV�lX-���@еU��`�3~��jU�Z�};f� �{����W/\u��yc�ܵ	=1Q#�O����e~Vi�7�Ni�u��_�[n&?��ުX�%st�x:��?�d�\�f@��(��d���0����F�����tgS8F���c7օo�Qw�P��l	QY��2�O�-�j��,+��>� �y��#��۽���.e���W��W_��o�r�Cm�	q_�M���.�.lc#�夹��fԽ4��X �JVA$�(�z;�9�������R�G�Q��i ���X�x�Mn�`ۋ:��Y�,ͫ|ݒ��]�I�T��h�Kt㬸���2m�y��Ι]�VM�'�	�;0N��
�b��jB4r�:���9����E�oQ���4��|���c_`>���WF]�t�'�[�(�7��~�����s��y;�D�K��a�9BxPI:��PE��J�e5��t�yܵ4`�/H��M���h���0���m��5VtW��ȁ,(v�N��)7HՈ�6�U������#g��M�j664�5�P�~B��;�H0�	7є�U0;X�<(Ye�
Q�N����?��l�}��LSץ��!�ȵ�ٔ �T�m+%�7�U[�����\(�w��n��	|Y�y��$6/��h+��m����^T���� ��٢���+��z��!����Y`�h3ٷe23��P��Z�^}��Wߏ��:�p������-�Uە�];��t˦[@�w�y��6,E����c�_���\��/�`��ߝ�)�1l������s��i&>4�����>�}O�v��#��!^҂�` �}h{�y���^�j˓d��@)�1�&n��i�r38j���K��T1�Yj�,g�do��xmG���lA��M�v�������7:}g� 4ߵ�m�Ro]L��X�l)Ps�D�TzE��l���v��iUL��*d:�h��d �u��1�/�m<2Gj�x��Ǧ�"�D����\�,0�`cR[HW��2_m�t��Ze0�p.M�:��+!��\�)8�v�r���sm�|����׻��3a�{�����=A�Vs=�N���7f%XS��{ z���4�H����N?���P����p)��/�ܩ�H����C/ץ�.�ų8�n�d�Vn��Z`��������=}"{�)+�]��)�K���6���PW�Z�����y�uDC< �򵀽g��msؤHn�Ei�]K�\E�bT�X%��{/6t�OARԄ�tɆ>&��>�p�a�7xL�J~<��\�Tf��w�*��ړ0ɪ�>9t���Şs�	�ƗL�G�F�,C�&���u`�iu7�')ɀ�;�(i��݂�����7l�5�26ay���j��/�3�u߄�$�޹����x�ז���k�i�F��lQY�q��;�����N&�8�kؚ`!�/j��Ϋ2��7{u�d�(LeZ?r.�̶����	�x��|�a��6_o5�P�j�O�-��;�"Z����|K�l���ׄ���7ޕ�� *\�'IѬ����z:Z�	9!��`���M�><��=6o��������oWx�N�����Ӣ�H� X�c���9 �Y;�7��k��w ��/�!0Sޡ)>2sΰl���z�l*>2[L�dVduR��c�dr��hj��U�=b���/�N�O�C���s�{/��J�|�}��0�L��@����'"c�>���������zȵ}�V
/r�"Q���R�
M� Wd�q��]}?-]5)���b�{�a�I}�����e����W-%M�������X$-�G}^��1���B�Z_<(OMP��(�vp_u�]��Q���2���P�_z�~�^��n�̸�1B�+��n1-m��RG����x�i��/)�+}����E�а���N^
d��17���׬�3��ev����P«�w��,nh��]�
t�H~|�/ht]I��O��J�|�a��X�%����d =Ş�[���{�%��a){ȱv��[ۘ�6�ge¿�:5�7���UVh:?^�_�-����GYۃ�*��o"�e���� =�m�
���O%�A�X�;�{�+�l���7)4k����{�W ����)=f��bp����F5��s�����#��
L�2x�������]ݏ�	��K8B(+W���[h��s�K�Lȟ���\;5q���µ^o����n�w�ov�9�Q�y��a��e�o�V���b!D�ܷ����'g��)�E�|W�nkȮ�tT͐�ꑥz8Ɔ����]GV �oF;��z�j���=Ș���#-�{��3Z�
��,J1m�kXX�4]�.��/�Ǵ����B�Ԩ
6���$(=%l�ª&h�?��Fu�iOGJc/5�x ���I�+n�買+����C���S������1FLӞN['��g~��#R(DZW��~��3s��+K׭o�%�y��@�
}� ���`�9?o�NG��;��#��`����Z�:E.v��hQZlQ]@���o��m�[\�+Tt��ۊռ��+1�<��b��H8GZ��.Sgk�бCn+/sБ ��#kj�4V9J���V�{ ���&܁��T�LM�.��
����D��Ce��D���xe���\���q���wj9C1�靅&�u�N������Q_p􎽆�;��:����Un�E�Ҳ+�Mg)/�:�Uq��g|:��~s.�ET��-ש�u\�nGdՔ>B��� �P���-?A��ϙ�� Bӣ|ֺ߇C�,��_�&r	m��բ�z��[`f煵]�3�R�bPChrEɷ��z���(����*��X>ؠ���΂8���Uy���&���_󏻃]=�G�.L�w�?㍆qȠE8�`yB�6zU�y_h�M�-���/n��Y�T:rF4�ᜧm8�i؜����|�Té�����
1nۇyFF�C��#��LHN�?�S���)�Ŏ�?�\ʖ��Y[����O(��^)]g'{	�9&C�yt2�q�z��"}��5wo|��dv&�]�ܧew-4�(���=F�)>��1���S�Hf������O�mD��0	
�������:�u�2(y.`s�aЅ��{�~%�Q9+,Pj��M|��$~�3�x���1H;�GS%��f��:�ǀi`�<:����J�F�r7wX�\�Q�� �^(sy@Y�>6�I=���!�w~�C��"7���#��Xw�����e��Ó�����9ʧ�����)3�%X���������ѕ��D����$X��a��|�4�ű��M��:���i��'�)�ڣG1�P�&	G� r,&�y� %�&��E�"q�$��v1+h.ª�@S(d=u,I�?^���mp�/:HO��4�%F�0ȵ1�?]����G?����t���kbTߎ����g���.�IW��k��3t9�4���a�G�ֺ�C��%� �Ҥq����K�?�u�gT�wACW�����'�ǔ�-��L�4<+���G�`�B�EE�˩L6n�l&C��٨m��#$�M�xnQ�	�c�i�y��R2J�K��K�_,k(�_pP��������PBb|=��t�M�1�.�5]�I�Q ���U�AQ�&[J��l�qg��1�[�k�Xs������ݼVhg�������dՇ�8�@�tG��9�!�[?�Ks�j6��T�����8�R�-��+$B�����H�DV��:�L����,���6�i��������f��I�"��$��/�)��r�2>�4u����}��:�R��	��F�m�k���u��ķ%i<&�.}��#r	�I��l%p
��G0G'��e���`��T7L�� �d�h/{Z��K����C~�FV���P�>� R'ב���F⋖�U��@����������G���r�y�c}ǘP}��0�����[p�L�{��fؕK#��Gwn���\ߥI����Q�q"iby�A�U^ĩߎVأP�����P�mrUh�孴l[`c�0��C��Bō\�Ǡ6Z��_�ҞO���]��]��4�!�����@Z)�&�*lo5O��b3�p�+�j��7p�,�}�9?�3��y-ϧ�x�mK��F��FLj:�@�o�mNG���8��ͷP0�F�I6�;d��xi2
��Qؾ����@��i׫�{�Y�D@��">��N�4����3�����f5}���;B*j� !AV(��\�^ܫHH:m�Ϭ�����jS�o�"�Ln~�K��lUk�c����S����SM�%�5�64O�W����Bb�Zh��D�[�H}���l� ��%Q�ux���o��V�ӆ�=�SD��W��Q����T"�0�h�U���0P	�u�%��GT�J�6q3� �"�-KI�>���w�G�?��0�r.j�����֊�w�%����Ƶ��7�0�J��ԃI���-�qi9C�5��h�����YѴ�>����X�A�I�['���H3�F�1���� ����q��I#^��A������JI8o�p�?UzP�,Y��$OM�eզ9r!L$q�Y�7���h�,�`%����er_��nG
ց1ݩ��P�������
n۝����w��	�����FYgr���P�F;���{��Tc"�9rU�����iz�_�큞bmgƭ�Ͱ�m�2��桓1;~B"����:/�F5�63��ז֡��W:�=hl�9�`3�ڙ|�f���(i�U��MxT�E1�S8�kK��Zĝ!�����
9H�3�u�6O^K6�Fj&�p�	Hʇ0 �-��mD�`��q�8���˸ap3�%\X����vn�wNu��Kjp�ܪ���e�H��_��ߤ4�_?<�m����n���T=���Y�ߔ����(��<˭����=���(��Ig� JCc|ՉoH��F�ᗃ	��
�
�>A8����T�'8�y�k�z�����t2�9�ν�XQ��u/������WBx]N�?���͹g'��S��zu<k�Bٵ!.�7��rp�`�o�?e�[�~Cx��|��Uj���2�*J�g��&�g'J�>�$8�ik��d�?q�ǿ?y�W���^u�|̍���ĶM>��GVzN��[-O��^^��G}m^q˸�M���aB�h���>�p�	�k1B�)A;���`U���-���8��3��j�zU��>�>�o�rJkT�^F	|�S�Э0����H����%������ݫS)�DW����q{?��(N��E�Fs r��O{��3ؗ�i_�6�ns2�i�����L��jr��v5m/Q2�U�R6s_�������y٬5���|G$�[QH&���cR�|�*R���S�c����g,��t-�v�
�5g:9U���I�R���y�uZ��ck�'�ЄV���y����p��Y�;��W+2��?� ����A)d�5-R�w���Km|�wiw��uwJg��nRB#��${L�>H��A��4P��\AT�`��c�z��4��
]Z���L�T!N�b���4U�݆����M���a�B��&�+"�/�@���"3۱u����Jp���N��cv�#�"b�7A��AL:�Mi7�����v�wЭ�*�X����s:�B�]�:���&��H(b�T�I�Fq/l���f	[�T��sS�?��9���b|=���p���J�V}3 ���y�,c�i�r��_����MhD;�o����[����q��>O�>��U�qy-"ʸk��)Or� �E!����*
�
��Z��2�e����_PJ������?�"���m��Xj����'�u�f%�7�^�����)�u����$5������P{ڟ�Z���zp5B=U�W�[>��
�fbԌ:�H{��m���]��)m=�%jMI3ӊ].��6�T���U@CC]Ɯ7e����/����O���6b]ٌn0��t)%�Va2?��T�_X��2>��\|���q[$���Ntn�-z�-�e�y�/f�~ߒ�]p���B=�� F1T��$���C��~H������|�>%/U8��se!��/�mvV�x&���\�pG����ԋO3���P���w,���CMU� [-Vr���CP�W-�Ų��c[�ޣ��,�
8z!�?���L��h���}Oy[�t�Ǫ������|}��<�G&߮.�z��4��
��LR�2/h�?�D;mY��9:;�9�O����_5J�Ѱϳ���<�*d�r�\���GZ���(�znb�ܼW�,��j`Oͯ�B����
�J�5��g�!�C��4&�3�O��� ���Qj�_){c�+L�e�Ϙ�Sf5���i{�g�w��F��!����ʞ��ӈ�{Z����_�y��a}c�@,o���:[�9{czhB���+�[�{i��V�V�g""m�ba��SH���j���y��:�s�+�}���
8�=Ȫ�C��{
gZ�Qڄ�����b�E_"&�3��t-FF��"$�NF<l����o�\M������<G��X�xd)�.>g�j���UՖ��x�T�r�e��Sg{�bj o�C��/�_yw��ot����u9���]1�=C������0��٣�t��[��!�1��?�E�����c�8���Xj΢�u����m���8����X�A8��a$#��V��$��᜼s��F�ɔ�B�����Y�\�O�I�@Ĕ��B�0d�1��.�J)�Q�2m��ؚ2�/��R4�w���Nе[
���hY�a}�sCE���?o��^~��9��h��Z>��H���ݵ[ y��+�.{\4w� 4�b���u�i��cK)��+R��_���5Y������j6���
�$�5I*�o1�s+����#����T屄�p41�ʉ��ɋҬXH0�P��U�����,���N8�xK#�|�D��&��Dp#4"��YK�:�̣�-�s�>y�O����|�7��]Pv�!�HZ�1������#���fV��r�Q�2d�>��XU�$`�;Kqm�˻��bwA���ts�ER�Tə:R��-��lhv�n�b�6M"�.�O�(H�db��Up����g����0Zi'�~ގ6NLOԊ�Z��vi��6��}.�����̊��6���������;�sLi�A����t{p�+�(E1�4�T�@����g:��.�(@�!�i�_���|���#�c�Y��"I��Ћ\уg�,�.���1!JG]�?ZwŔ0��|��`!��Zd�8Q��>�nˉ�D�u��pnk��z-Oҩ� �N�k�UN2e��/�7��~D־�D�z���e�P�^��?��4�ٌᶥ	B�d�aEL@A�*���Q��)/���	u��쾥ޅ߀^{}�i�C��o��E�E�F�����
Nw������
CU�փ��l���� �5hЃ�o�{<��/I�E�X�������KfMJ�̽����D�b�I��j�E'p�ݒ� ���l�n.H)q�)�h��y�37�-,<�5���	1�Q"%)N�/R=���) o��2�����LH��_N�시�P��]o%wY��mm>Xhv(Ĉ ������#��j���)��f�[��]֚��^�D�vX#��2r�?j�"+��n�9u���������r�hQ�����O��W��im��K��Gb���W����v᱃����Bm2��F��9ak�}����p@����c�cq����E�P&��Cx�}3�.2�VR`jx��*fp�7ie����Z�7Ӹ�oH	���ä��Vb�_�wI�=�V�.�F�r���ay�ڨ�+[�U��)QF���xi�yM7-O�Zl	���#L�ӥ���AL���'!â�\����	ZP(&�F������bn�螂�ý����d .���5���cf�����F �\���-<��F��A,߇/���K�������8�}�A���6�����'A\j�;��4E�""U����)���t���9cX?E���� �92�{�֙^�PH�7t!|�#�L���}i�a�K�t�u#�)U� U����26����ċS���'�}	wE����ʠ��O��,,Ȫ�����ގ�{k����z�=2B����
����`I��� |����~���&}��Q��L5*��l���&�j�������N'�}�Ah�LH"���Zho�zQ�&ޒI�g6�yƬ�<�]m�q۱�����:���}���p:%�E����W�7'Q+P��㌼3}�'G]��=�1�H��� oS�����ot䢗���'H��R�;q~�e�����YTA��R:��/�$�M-A��*��VJT<���P
ϭ[S�J���T,��mƤ�Xn�8�ҝy��jX��S�aE�Cn�7D����G����hGe.����74��ṧ޸g�A뱥�t�gR��8�K��.YC/"*C� Sa!��G�����7"E�3�p�? ��J5�=�/��DG�7�R�W�]���fξmI�;'�1۳�+��-Z�u3;���PE(�Q�\TǾ�Qd���`^/�&)��"k��(g��&�N�SST��n:��NL����Yaں����oEa?�=� Foo�đ���
�X�
�x�V�I��"��0HrJ�o�+M����6�|�V���r���$=�Wĭ
%;��D K�x���4�C�f��b���3�`<��Dyˋe�,^\[��HPhtaXR��4M�4+�_�EƧS(���:q�躦������v�}�
�3��՘	("=1J���tP�|��p�X%�'�l��9�C�x�������©�9G���h��H�X�ݯ���/a�=��Ë&G�s����'����� ��J�u����mW��� �T��0���Yɱ�dl�`$����3����.vs�5�ς����z�g|��/[΁G-.�7�-��ZסܝgS�6g�ʯ�}���02p�MV4�g��P�f�p���u����`�^d�W�� (FE�*R5����A�8�m9ԕ3u>̆�'$�VdM���� �M���F�Z��k����L�S�8��g�d���Ōr��N��@.�MΔ��\�
Jle�qU �
�眳��ְW��ԩ]���a='��zn\�8��;�]��0v����KÙ�Q��>�Q�����?ӟ<��h�%N���r}X��`:���O�*	�4"Np�_��޺1͐�d�~�|��]�J�֬/y~��������~�P������z S�x�U���a��� �YҦ~5�D_��m�Hm$9��M'�b�d��a� ��FYP�b��?���ȧ�
�:��2d)�h�`:ژ�Vض�ER���TC�u_��2rY����4 ��Y '<�{��}�t����J�s�[�B�Ӻ$��B �<Z�&��/�^��l�ٮX�[����x|H�-r	HKz��&\�f祯�Ci}����OL�Y��_�]���㰴3�l�GE�v5	t��!�vy�I�+$��WW&�5�����O����k_,0�:� ��x	:C&�y�'�����r�=�����9lg=i�0u��[�eI���П���,�HQ D��uv�qo��͛�c�� ��W1\2bw��i�F��5[KT!�Z��T��d��4K鸇O2�`1� Q�U�í�SA�6`jB��ɷٳAqI_`���������qx�FO�[�3�~t��yfJ����w����x� x�v:����d�� 4`�f�.>���d�RnpS0�w�{���R�a���:������BŦ7ƧOA|�tZ3�1�
�o:֑��c�0��2Jb��7uy�ݞ�$|����rPz̃CD_���3����qt�8z�����βf�`' �� g�n@'�g[[v����@4��9o�Z��m���de�Zw�7{ῗÕ�J��w�	^b�^��/Ԝ~��̞������Dh=�E1-�ۖ�%^T4��u�^y��QS����̾��/IU�;�A��N�����������cm��,�gbL�s�3�۬� ��B/���]����1�$������R��@hv��x>�4�M�t9��RN&����q�����YzB.y���Ŗ�I����_��dgR$V����!JZ�?uOe;j��g�%�%t�ҫ�N+�w�h�d��KmL�Uy������&ٹ�ێ�$�=�BK����!�B]��%)�U���J�F<�,����;�
s!���v���j��x�4��kD����@:�z@�b�3@[9�x�*%8w�e�S���*��u�7�>����Ѓ��e��#��PG�-�tN�(xa�#�Qt�S�~�h����AMc}82�ijT=ٝ�����3�ˌ[�$(0�Y���f?Da��Mj���G���}�畈��ޗ�{�-@]Dҥa��h�'�Y����Ubq$�P��D�|<�\ڂ�摳�L���9����tE����2�CH�	�������B��{h�^S�ݩ�=}�h��A_-m�~��<��}�H�l��\y`3eNY^�C+sF��72���k��{����ߑ4?ӎln1h��`�<۽���\. +�:���뺲3�.��s�4�>��!2g��$���|�+ \��_����A\G�
� +� �.�(�@VށǇ�q)�|��+�m�;������D[�T^M��Q_>�{�@*oR?iG[a����&�y\$1��C�hk����^�8�(�A�HZ�5c&�aY./�#��UŮ.$}N��Z��Nw�{�&{S>en=B,�i�k�;��w	�4�k+�����׍�D�ύ��i��X*����HF��к���	m��bh�S)�_�fJT��d#��:��y�|U���,��0�R�H��Bv�j�]�`��3�4;��t��.%�~�O�ٹ<ĉ'X�	�4�<¨�$��+Vz��EK���*�/+OD��CJ���c�U�P����D��.Uk�c��W�Z0�"���ey����f�\aK-{۫���`�t�b���O��"le��:Q�%r	�f��,~���z�h�L���U��a��^�w��쳣��J�Y��h$�Vk4���
6�h�H ��@Ր<y?��(������i�K>�����ף�|�:(�����䕪ӑK*:K�[X���,�S�I���6)��L�nF�nc��ݸVd��d;0,��2�ANGp�	�E�Az�둮ts�
�K��d���޲x`%���-R�;m)e7��^t������}Џ7=��@jɟ���\D׾�м�_�`�D��Q�!y���q�_���zq��i��ԛ5�s�nQ��`���73Hl��\��wr_]C��n(G	#�|�*A2���^b@ٗy��,�d��w��fוq���Z�[5bd����Ԧ,�\`��;�N���{�P�O���[H��2���}4W�-^,���4*b�	�l�����~�li���I�g�pF��=��/���M� YN\h�=;u�T��=�(� �rϊH�؀��@1�L�f s�jjĘV��Y��p��an��=zu�+�b�5KMo6��
��0�ˢĽ�Ja���x��Z	49o��K���#�]"�G'�Ǜ5�$2:�v[:A!��hB��0@c��,&��sb>��À<%^���L�%����T�{!�Yc>mJuPo�p��9lɨqP0"o)�,�L��՞H�+ؕzz�-������2�M�����?���e�����{!�q�J��5��ʜ�T���8���o=�	c��%��C�,�"��xe�Y��I�>�|ȣy�~������U�d��3�%
␏����!d���Y$ E��[9�o�"��HU2FV[����"����&�������9O�K���ԕ7��ۿ�������ɨ�:��(]�!̍-k��G�5P|֠�������0س��po;�N����lY���X��nݺh�X�9;S�6�.y"m��r1h��'o臼�9��[_L�r�:w�xԸ{��Y)���+2�С��>�U��o��;����PVb5; ��9{���b_/}|�#�Ak�(�\+|5����)�5��C�Oh~���9vs%ǍC}����J�7n�h�"[Y�LE�U܅tI(���K��ui����O��	L_��Ϸ�y�@b
�^�v�^� �.�^�+*N���1uϽz��ٳ��~fG�
�ĻJ���_X���Ab}������RU��f~z%��hb�B&Je���atltl�ij�yN�i�2�%|���$
��h�sa��آ��K�F/�>"¼M�LPF�%7dVl���Om�����yJgΛ�����O�����&��:D~<=6��7�`�ꗕ#��`��
xJ��zG���X����b�`���Yr���dKWS*m#����	�ޯ�
����?g�U�r\:�ǫ�v���0?���4��)�i�k�`4�}��̎�XNϑ9�r_�f*v�ҕ��Ʊ���	ll1>>>�)i�-��z#��W�5�	��M��0�?h���!m��~,Q��u�yG�4��C���X �!B�iOP�v�Q+5n���c{؟N�pG|�f�����ҋNaQX*~��f�^MLeU��鴃n�(l<���!���{i����EZ=���`�Dwx��]�#�uI�{�0Y x�RP+���g�DU�
a�n����*Ր�! ��w�#�HI/��J���댈��yGM��V�~X�F�����Tae�v����h� mMx���/����w��=o�O�W8J��b0EX.р�y
�D�NK�n%cT�����8���>sALmxۉ�[����sv0�>,�lsꫧ��*r���,��VdS��rb (e�`��oQ�Z|������2_b��J)��?�a{Pk�J��k�n�R/����)�b�I��Eߨ�I����3x��{{H'�팣�K�ZWZ��]S�Y֋WX&W\ R
�s���}�!6�S4������.y8�ҵ|tD�|y�I���p'	n� ����i㣥V�Hy���s~�F#&�(q�`��3פ9�kL!la�֠�Q�X�W��؎4���bt7}c� �u�����!�c���O�_r{_cj��Q���Q?��UG�m��Z:�s?G��2V�m<���F=��dЕ�`R��ģ��V�7�A��V��-{�L�N5����y��hS$w��*�&�,��ƻ.�a4���\��Q�U�hI������hAʳZp,!���>�� �)��8������c߈-���ylh�ͧ��U9?̍��jd�O�
g{7<�w��/�ӂP ��
J>��4�˃�[5���=20�vn��Qߟv�I|��m�^�@!}�+�o���b'W))#��u'rZ�j@vl6��`0�` Gin�~���s�tU$Q�N	��\�pd^��x7Ҋ���z���E�Iǃ���"x����&e����I��@k�1�~������ɟ�P9Z�X6�zX<��^�J�3Cw݉�������a.�M\'2�J\�i�vD+�q��zh���)��n�^p��t���ջ��az�Ȁd3�a,Sr� ��d�`��x^��?�����_�k]�g�C��w���R�)��Ǥ��-�ʑe��#�[�'���w�^am�l��W���}��L�
r֠���:꺑��߼�1hh���x�r�9�
�0��)�:E��ۧ��K���u���_9Z���~+&��lB%�U�ݥ�8���}�AVc˟3)gb4E5�voۭ������3\a��G�V�#��ʍ�hG��=`�<�&�N��ߛ�'�����rp|�sVSy+m�UD�����~ݐ������M�=��!ߘh���x�hH��pc8)��)������ga�t~g_��¢h�_��g��Z&�[40�dX��h.x�Ml2z�m�QU8D�#P��\a����jAq�;:v�{@bz�ވ9]��עٔb�:��9�4�$�U7MM�b��~z���}������;IFy���.T1C{�GVX�J����UpL��
MD�#�v�8��O�C��Lu���5��9{P��`;����>��3�Gy�����{&�3P�vK�����{e�= ���*��Y�΍H��\��#����?k!5�>�x�nd�\�Lq8��\���l�@=]�z}���LC����?��g�V����b{�N�A7isp�q�0���*�{$�y+�3j���xL:��PG9���R��~�4��s����G���lua�[�ۥ-|$�Z9��K-,}J
 y�t��x��	�ss��r��~4x�i�Q �Z�4P��/!�7p�ףr4�G��I�ņ�4E��#��-#Z�vB���@e�8a�*��-{:�T�"��*H@��o(��g;O���]�p/5�<P$���.nTE����ګ�>	���<)V7){4�
�I�_��b
WA���C�f&��Z��e}e��!��T��?�-���%�.1�F%M�s'ץ+��\�e �C�5��Cȍڄ�V��a��
1eE�'O��ۜ'Ru�O� ����cP[����X]���$N�\�HT+NY���4��U)e����S<���UweX���{�V/�}�l���c�t�����$,Y[����_��嶰��N&ߟ���
��nou��!e2�����ښo�"�t�`��@�ӱn������Lgo �Ȟ�t�X�
�E��ʋ_`;����,�<��`*���$x-��{�U��/A�N��x���Q�͓��q9���֛���)E �Q�=P6M�D���7BNL>{w��Cf��?��>JΑ3�\!�:��@	��4 *����f�aɂF��fB��/��":Ґ�_>KA������X;IE_w��׭H���Q0�0��f�I�0�C��Q'϶���-�X���}Z��V�HG����B⻫ر+��o�� �}w�6	:f�Z���M�w�ڠ���������S�R*�Ar27���uU�B#=�.���ɔ��Si�G21v^v��r�|]'�f����q��f��D�������y��� ��]J�u{u��3��q��O��Q�$�)A}�%�?�tz���9��%�%���SBh,Ղ/����,�{_�#P�`�sy&1IO'��B����v�-����;��
�����N>]���x�5��~�HEw1��o�K	����@���|����@Zڔ�)ڕZ<�h+��G��{O0��Rfn��k�IX砖'��iv�O���� <`r�g�\�]D˽ᗕ��/�zaNٮ�50�i >^̏H8�-��wتJ�e�e/R�JH��kl���j+`���jC���&��9m�u�e�=%3����/2`�:i=�?��;:��i�I�#g��,�$$�;>^i"����;*h�o_	z���_,M� "$�ߒ�
D�F;�5�fl{3(i1*̌0��#�;�R���34G �?��ձ��"�K��8/
��,�¶���4^�7q�8(c�f`#w⢒��v�(��g�Oh*�K}�)9?�L�[����̻��@��]���J���:v�%��ù�\��!N�m.Y6oB�i�q��t4S���7��}�Ɲ5��"G���N/,�\d��V��q��H s������,�8nRqЗg��{�@?���Q	�.���Yd�m�d����cj�Ec#��>	d�����aLI�E�&�?�Ӝ�(�C��1��6]��9��=�}����9�ʸre���JQg���r��$z>钰�ê��R�Ŕ){����|O��Ղ�Jѷ�(���u���J��aK��I��8���*߁ƫF���*l��m6��*��o&��j��َ�)�y��.�������`�x\��g�WA�C��( hJ�˶je�l���[)��ow���׶Yę��{y��I�R��~�~3�y�6�$��=���/f��i�Yg�YZ�[��YoTPp�O��׋���tRuq����"rN��K2��OO�|�Lq����hq��i>����h6$�uA��3��5���G�!��g^���6�heH��A��~��ze���|�8�ڢV8/&�t����@�&�|	��]�
�K���d�}���f >�4�X�KLB@O�
��{:v���OB#I�_:Ю�wg��7������rD�R[���3*W ����w�Q-���.����[2��{r��D�p�#����Df8�sYk�x�.!�>��� �\�y��2$"i>k�<��!�T��e%%\������ x8z|�����$C��=D�ڗpy�`�hOh҂�x=�)��F<2�JY�źÁϑ�;�|�3�1�0�!����)�b��s��f�fg�9H���C�mh�P�S&����@ݏ^�q����BppE^�~���f� ���) ߰��5��!;��>dZ�����@|^F�*�8 �!�zk�!�ֶ�-�^@����y��6a�4��7u��s8�����m�����yo��{#����v�hQ���{��*G�]`��8�=�*�+�cp̩���A��[g`�ݶ��[�l,)R��h	H�/L��9��q�^]3����. ������,�
��V����v�*5���b-Z���$|Mk�5Y$��IO"i@�fFve�BR�W�i�)Lb[P��_%a����yM�[�D#�l`H�I����^V 2�(����Rb_8��&�(���i��چ��	y�[�獬l���|�����CgHQ���&���E(?:!�y����́w܊��$BÊ�ܩQD��-��*��f��t<�/L���!G��������p�Sx4����d:�w��Ɉ�Z�Olx�T�a�m�V.�vAZ�ȟ��EK�0�_�x۱|n�r]�c��1]m���sҎ�W{��EUS�X�x*���NP� Aw_����D��>|�JV�Fcx�!������o�OK�6*������4���U]a�Ho��!l5Vay=oeZ����9J���n��ռ�MB5a̤�n.��K�Պ,�]�9B����`�X7�l�\��ߧ8ܟ��~H|[@$�K�J�{t	��1
���"���[b�@�숅����Q�|i��M�s��:��2i��M�,~&��N�nA��O;���Y/����xe%,��*b'k$#�x+�y�!� !��P޻�_��q`qzȝ���B2��y�'�_�b0�E|W���Jb����T��2�����g�ӣwIY������mp6)H�x����>��"�,Ũ�.F-V�x7�;;ުo���Ц5��2�����+Rdo��AƊ%���t��Nm�Fgy���5-�Q%�����C�-�'����r�>y����2,���aQޔ�����E7*Q��|J3�Y�$�N�o�Ǟ27��s�#��~�b��<�`��N�?��J�"�vGA& �"�3��@�"}���`�1<A�𗫰�ó������I����pbu�[K`���;S��EF��6�ɣ%;1N'd	���������Q�px���Y�&
uo �o�����j���D(/����5��aO
�.�b�R��]�����E$�ca,�N��H���ԅl}Ծ��:�f����h�;�4�9���f�`,��`a%�E�w�U���9�8𸣦ܭ��e��H��9���e��p5t�3syG�"�PUH�R��,IǇmf{.��u���ve����Y[�ڌ�����y��z�y�	p���rvh����k+ߑA�$q]��I�x�s�>\mG}`k�:^E}jjp�^F���`+�Okm�H�������m��0�k{���� wu��g-��V�D�[U_W��m�t���.N�P�׋%Vf����΃�(�mGɣ)���SI_�Z����]�V��Q�ر6]�{�U�@��$U��LP~G��͹hΨ������'���(�3~��Z)q�������,ٱm�(�}�r�{.3�q���"�9���P�c�le�/���~�&�/f�z��^��&vjw?��0��l0%[�K���a��μ80:�}�nM0�r.�a����Y����Ř�}M-X�(3��0�9��	�0�V��t�=HoZ��|LM����i]W
33@���p}zG�Wډ��k���5+�	 vWJ	z���ˇ��� /���K6���U�ۖ�)Y��򈻢�*#�7�O>�L��ǘs��2�2�J�O�2��P��憢�ÖH����K��맮HD�Y@��|�����q�;B9�*p{JRM�auV��bԬ��aYd-o���;o��;8hx#��rm9i@��?�x]O(��V��㬾6Q�3���D�7Y�7�wMyM/�^�\�����d���'6���7���GC˝%,�7g�����Y�֥q�8v�tv��G(�&���r�F�Έ>>��Z��@3��7{��0��=��i�ˉ-�)$SLF�;�mO-
��T\4L�"0�ǆ�DB4-�I�a�O}7�K��[���(�4����$�Uϡ^W��A�ԌUF�߯l	['��<g-j�_��#r�]����-&�킭ۘ�6��㑸�������adsZL��5�#�yN"�B�8D<�&I��:��X�)2�o�Q�l��0�,���c�Fa u�K��/"�I��p��=C_ �`�=�q,��G��- �q��2��VݕU;���؀B0P[a��O��>�,��z�/SF�P�X�>�B��Xb��jڈ�/{�{��E�|]����25h��*a^�:4r�C��(R@딻�w���91�؁��i'\��"�S�WsO?�R��A�VP!N)T�X1辽0(&q��ٷZeCh�擶�|�(�>K���K��^H��26��Le*6��l�en�A�2���ۥ���X1bk��lWi]��M�����x:Z����C���mC��+�%��Y-��%4z�G��G(���Z*�/�ea��F/��&�3&Y�<+�)�d �vJ#���c4�� C�
i4L�C��L7pEߡ�6�K�'Hlxd`�y���NU��у���m�m�#̶|�m�f�}I���+�#���1�I�MY;��vf��/k�&I	�*�(<���§N��i1�(Q���k8��&�e���]k������U~g�U�g���e��!��s
`	�onە�]�z~�~Z ݥ�sr=�?���^��i�LQ
23�5��!�'�"{��~W�6�1I��GpQ�����Q�-\f��j��$�Xڵ3*�7k��`�<jʲc�~lpYāߨ����:q�#w�(O���2�D�NS�o��CS����#�蕓��"���)Btn[��9�&^�rx�S��Wk
����ĤXy�t2�\�98���@yj+�a��bj�ϪÌ�Ob����ٴ��@�Y��$F�YǞqr�y�=H2%�z��Td
��_՟/2O��3r�ԩ�8Y!H\ ��I��5T��P�e��Z� ����Y�>=��Hv�_s��))�����՜g ��2��Ԙ���0k�.敳���p,?�$���u+��>t���Μ��F�Y]�{�� Ф��gϿ�{��I�:�����^��UD4�B�A��5���`��P^��6���$�l(޿��6	6-���+��� �ög 1o���1t�f5��#	�Ț����q��\�+Ygޛ<��0�7�vP����ǦL<��@O�|Cބ�w��ͼ�D_��Ķ�f&˫��C#�lWʏyP�Ρ�eҏ�%�%jEn>x�Y�c��y���a��6gB�eg��;��z�94�A����zY���RJ|3�@��6,m�A��f`���̮�o�����;N���?xZȄS3)��jxS\t�P��gO%�B&�_�!V���Q`���.	����8@j?�J�-J9����BaK6`;)b:���,@NƐ��)��P�*_�Z.Jk�*�u�G��,�]8z���*#�AAL�k��8g�5���<ap���ڞ@8�T���ծ�K�z���\��q}�x[�%��n��R��"���X��
@gT�PAɪ<�Y;�+U׉d�m]������U[�Z�f1I����_�����.�N���X�_̼K	��G��I�R!zUߡb��%P�8y�:���R\�k�mE�:?��U����S�=�e,7��wli���CQ�*�4�7&�A�i,���4�E	.Fv�%�n��#N�MߢL7g>�
%���ߏW?�"\�@�p_��kR��p  ,P\1/IwgK9��}6��˚��Q�<dǍh܏ǀ�C'�u1@���뎔�L]g:�G,(��w<%�X��A��@.�пk!���������e���3�F���v����ޙ��zo"K�4���`�
&�;��P�vu�@��{ۀ�(���U��n�h�V���?%޳H���s�G����k�2`â^%sq���L"���r18@J��.#J�x�b��|Y�UhҾ۽ѐ�����^�����6t�-�Ƕ9���Һ��0Iqmt��%� v�A�O�@�@�[�=*���<��g/�����AQ�y���~�����bɢu��P<AA��g,��vͤ�_�rR��A��)$.JK�CN�����(�֡s��?�0�%�Qo��Ҷ�U#�0qw�1ÉP�:���rh�_�X5����۵�`��P����`s�8F(^P�V	��R���^�΅ �n�b�mY|��^yX��f��Q��2wQ���qm�y�m��C|��0}e�2�~|c��;}���0�J3Λ��h̐}�SM�u)�D�k��)�������a�F!����R� F�`n?��K�u}�*���l;���B�9��'�ɁOAz:j�"O��=������q�8�y�R}7�&�-@#(0� v��=T�:l����4X
��aǏOПk��r��n�v��\Vwi�MjE�^`�R��>k����������S��N�O
�)=�؞$�V�0��'Qj�C��0K����M� ��ĥ��Ai�	;�ۭe�Z��C�q��[B�j�\{�� ��b]��6s_�0�0�����Ry��m)�XκC��HU8c��j$m��+o:�cR��A)zF&o�쩤�Aǉ��-@�[
���z+�&F���u�Ym��D���(2rYܙKV�X�i�GUKb"�=��]I0�-KW��lTE-��g)��VfN6��#�G���nύ��t�R�d0����t=��CŞ�o��|�������3б�+f����iP�䱬�ln����LC�3l*И��-A�6�ȝn=b/b^8���;�{����P��q&(��2�CocH|~����?�V�>��ׇ9��9 T�{�[|��[���,u�P�t�h��^k+�+GL�H�f������ �F�����3=�|8Ds�ߵ��j�Y��ޒ+����6!>�8�B�4O�`d��KZ��k�T[��p�G���ȡ,$�N������*�O�y�M�����e��w���9�e��t���ٯ~�v��C��)������+$�UޫL@͓��}��W��ѻ�����u�6�RZ�^�)��]���&�Bw��W����FQ<6m��2�\�j�����d���x�\nZ���]�I�kȷ���V	j�/��J�e�z��1ʣ7ۅ�K�"�8HT� ����s#��t���VD(S����5t!��K�h��%�D| Ec��\H3�[-�t����0"��|��}p��3�Oϊx�-�R����EA2	S�JY�mD�K���o������b��6î�iU�/k-y���^:$Ac��q����y�k�Γ������'����N*�
q"-��aP9EZt��'�c[)�����)�?gv�j���%6��J�J�"��S
��6�Gg��"9�|o�2�*Ŵ%M��t�4
��^xc۹�Β�S�1*���f�������%:�q�5����e�G����q!�2c�U�BY?��[��o�\�}W%�����e艮.y=��,�H%��r��8�q5�h��1��NSa���l�"�dO%_��/�:��0��$�����f�:�/�m�Q��q6 /oG�$Hw���w2˓2�_�f��$����Hk�(��ʹ��l��'Z.�K�텠�p�'�u,kb���C���k���rX^N�,��O���.�E�e�[�#�fA�]�\d�
.�l��X�Y%�,���� �l�G��5�HR�2L!%����0���
�$��\��p{}�{D�X���N��o��6�s��ԶV���Vm�E�bP��%q�h11��������K.�^���	o�gE��u)IG��#~��t<�ĂN:bpx!��[:�i�F�FH�����7ɹ�uX�-]UX�P?�7t����[�9�錉�_h{���%��S��Z8��&��06V��ip&�<q)���Sw�f��'�����s	���6�2Y�ᙈnT�hv����H)�cU0����݃	K����e��h=yj�6,�����=����Kp�3����Ƈ6-�g@�o<ki�������]����TO�<�[(D
(#�[聿�å�{�T^�|k�3uW�F��4�ك��&�n��YK�S�L���OD8��(�Բ�D��)�;̻{k�+�����x,���c�.72���>�o3h�N-]E��
� �(�hsPN,�^��&Ejh;��l�Z��´(�l�́O�_����Ʌ�ԗ=+��j��U����=���-9�)38���
zL� ��#�D�>Q�p�
.�Nzc���c�����*��c�e��yF�k}�<V�����
 T�m���$Z(v�,\��B�v%��U��V�X�ԕ��o�I�U�MRn#�/��I�����)�H��+8��vY�Dp��3,Z������BXk�7M����S��+�U&�����=Rt!~�<�E��}�r�7�DD'hG���l\�/D.�i䒹R���x�"�r�}��-ۥ0�>�"p�����F�;�e�b��N�_�u�F҅�W0#�F1��Ӷ�e2K�������8�>��~L�O�h��כ��r��ڶ(RF��Td�0T7;��-*H[U����#�0��dJ^?����>��$���BW��|@Ґ��̲oFm'�{�$7J��I�MF��{�FZ�S<E7#�L}���a���/s
N̆w�;_֞0*�l\e2(B���S$�-�kN�9�q	�`���n�o��S���� �}������h��{#��X�%�G����C� l�.�fEҠ."��}����CPIt/;���Wk�7��gL�s|�R'�_�G)�5��Ix񔼠��s��
�.��s>v���j�='��Y����;�����v�"�i�y6��~��wQL���<�kҦ��6hCc���;E��F<���_#���b�i�ۻ�䟆�������ڦ�Va�E=B^�c���q�^Ky����Ȟ]q��+	Cţ;{n���[j�$�Oݾ�:M�ϋA��,�|n8&-��떏ý���0��)_���Ɠ����#r�$`��5A)�C d���Op����b�.|;Cy��e�n?se�-�ƃ�9��^�/�u����6c��O|�O�=�:�������
�گa�B]�ZhS���ٹ�AW	�o����g����{8��E�7.�`�4V�)Gd���#6vC9S��`����߮�&����ftNX����Q��S��B$9in쏻~�x���kT�ip��eV��u_������mnz2VQ��bT�Ad�������'�?]ب���<�ZK4�)��6�G�I�+>Zp��'���&R���³��<8�� ���M����v`�]���^����f�Ď����k����#]h}�՘	,v�-#�����DS�����O����:T魴�Sx	�>�0�:��G�8�^�aH�A�H8Nӊ[��X�Ey�^�F�F��^,�p��i8�)D�l'��n{��u�r�B�c�9I��Cnc��;����7_����qn.������0�p{m�;B?��F�,����� *��_%���ֱ(t�{W����+o�������A�1W(����3��G+�mCw� �����C�iG{��䦔Oϳ&=�Tר��ZZS��v�D�"��NH&���1�1�%���rD����,- ����XQ5�QS���L��[����� B#�&�0���Sњ@����΂5��\|��4,,7hȪ�����6W�-׸|/�m�J_��
;�F�(��C`t\����6����0�tT7���KD��%�z���=����"��̷4�u
�3l���@��1��^Z��N�cH�v[�\nK=q�%�M��y
Fޑy5s���Uy�;����K��y�ʸ�2nq�|�����TO�'����Љ�4Rر�t��A�/;���9Ɠ�=��
7��>)$2*Aop�Fk����;���v���R-�06�3<�������M�T�#5�Az�4��r�H#,��K]��;���A�1뗇�3*ZV����3).��{ᖄ�D Q�G�G�7?"0���j3���M0���>\j^�⃃C�?�͡���؆�;�9*+2��J�����Q�2I`������|"�� ��$�ۧ�A��	n�p[���L�
�×w|�<�e�m`�\�˵��@��X�������U��&�U5Y���$���il~���-ٝ@"B�5�^�7�!ve.���~��u6�кgC2�Sn�)�= ̆;tf���nm������.4O8m��^�3(J�}�|4�<U�ƴ1���K�	`V̹�,	��T-�δ���[NYE]Ł�X��½!ϒ�G��6M��S턗g�<���~���	2�D��Y{��h�B�����?mD����2*X��\�����'������4}֒�sct8�#vc�B���ת(�ӏ�WY�c��>����)O��#�̴��2%fK8C�d,|y��DkHe�^ ��	�Ʀ ��{����u\W� � �F� 5�,��#T��?M�K�:���Ҝ)�Kxa1,xc�r,��������W����L�� ��ԟ�[ȳ{D�~�_4o��'��P9�U��d��Eev���q���*��g�/�%��1�Cȿ"# �!� ����7�B2aSi.F ��9���i�|N�U�'�^ix�RWE�7�ʬ=�"ܩ���_��y�H�xZ��g��L�O{�I��][��WA�P�;�[S��" 0�������6%�^�.�B�����w;q�����iTH��&��PXA�ȥ���+�ߚRf�t���@p� ��F�ϵ�WBu�?�$�o^�?�����Nt'M*�#&�2I����n@�?�&'�L(6�!���#�D]�Avׄ��Q\��MY����:O���V��FK��C�;�Lђf/���;G`���̨��{Df��F�[�)l�9��O�f��oW�y�=U�Ė'�t������u�Dm���Y�I#L������,�/�)�jCQp��$52�
߇���i;��`��F��Ԭ��2;�3q|Խ��� �=����P��:�+*/�M,u�p@*��{.��)7�cC��_��!U10 z�'�`(_�5k�+h%Y�����#$h���$a�/*G� ���'H��Us%̈́����I/Ƥ� %j$�޲�BQJ��Hh�ֶ�
=�zZkQ͠��"�7<��:�1A��X/��&Ԓ7�Cu`7/	2��ޯ$��=��n�hs �w�<n�.}]7�-ͭ�&�`iN�5�2H��<��tS�|s:R�2`�D�s��0�b����e3#�Q��i�_�).rv�n�!.)���PAb�Y��t��;��n����w���cA��)���L���%>�=��G�pAۿm��n�� 3e�����	�['lhB.�[5o�|I9sq�����p6s�v��,����$��s��O�1�&��b��Fr���� @E�W�ƣQ��y���荊6��/`JK^�I��|KK��Ǭ�����HĲ�Pus���{���NL�Q@=�ZPF�0 �@Q
��t����-/I!/f�;�	�Q1?���w��2�{x�IC�ҎW�{������b�f�h¢�g�{"�G�v1G-\x�Q/L.��--fFr?W��߬A	����p����:�'�!�ɥަ[("L?���g~�p�j���|��f�!�æ�~��މ*r�S.��18�Hɕ��6v�?�Px�s�6��=�8����b�sp�'n�D*�=vz0�	Q������q|6�@���1���h�kY߹��oj	1e����L��IKQ�eAg�14&�Jw���a���2��:�]J�Ŝ�@�o�2��
�������8�I2��^�R �����%^�n�v$�����t:����b}C�95���g��;MݣskpZؽ��I��T�B�T>gģ[��5�����`�_6h4$��/����41��ce��L��(��h4%]��Z/<�m�T~�@хʏ3�'N&*�dw)	sn	2���n2��Fc����űZ�\�����^� X�LPOEٶ�ANj��rUX���]֖�q	1�L?��
yH5o�E���"��sp����Y*](Y2U��8�~G-���
�>�iOCr�j��Y�����~k%n��6h��H����Ņ�s�Ƥ&EYj������g��X�l��i��E��y:8�M��hmR!�flI'�6R���s�Tm�t���1��b&	B����
>bE��j��E��F?vŔ73��m�ׅ�_�^�j
 l@����X3�g�]%�Ă�WM;>�WF3��[�>ʂ>�(���đ��!��K%="��Tji�.ң�D`���_�@��E���Pe��3e���	]�P*B'��=X�7����M�%�bN����g�b0�v}��>��� ��:�g�#^E-�s���Q�s��,�/���*��;��xZ?�3����eO��1��7����F�m>�]�a{B���kI�9�.����$lV��Έ@&4��K�!c�4�K]D�U'y�8�d�Rrz�QsJ	E�z��O�~2�]]��㕫�H(�r���*��Fhj�ec�:�A6�0�����`�f���
Q� 9KUn���/R*�?�?�,�NI����؋���˂��$�W˚n'�����T�һ��~L��*εn��J^V���]$���Ǉ3^'B8�˳�>c �3V��k@"��oj��Q$S:
�"ja��_��%�����=���C-��ր峬�Ŭ�&�,#���)7S>��=�/�ͭD��Ƥ�����[PL��nݎk�`��>;h�X�}�Ԓ������!��dZ�)lݛ�E���i��#��
���DY�.��ʑV��\��cWo��rp�����\�V���c�q����._9#;q�S�q��!��� �!y4iT�p���;-!�pQ�O�U��B6 �\�U2�d�{�Kkb�[�m���4u���'
�
��^ؿ�Y�����=�/�e�(Ɔ>�i��d9��J��R�$�k��M�O!t��<����$�~(�ɾȇ�����5x�� /�!�22����K_-p�Ӟ>����/B���oгRY�.�(ĉ�KA���m
��͆b+���Œ^~�S�*F��I�&��f���Tj[����}L��LS4�����T��#�W��e.��%ةG蚤�;@2l��"i�3��Ėe^C���~F��w�@x����ɉ� �{\�#8,-b���#e�����K��Q���	�$SY� ���j!�v+�M�y7���okD�
nH:=�� e��%� D��"��%��������M0��a'FW��D� 3��25r���Mh�Xs�(�����؛{����Yrf0nG��kw#��W䞊'D�6���!����4Me�C:�c�gV�񀳇;�m-�6� Z��2�Y�/I	�@���α�:��m>�6�����o��[B�\]HM�r�=o���w^"��K4��q�L/�(�DN���.ELi��C�7��qe�qo˾�����3w��_\Et�6\z�%�?-_��
�Ye���@�/x����0���"L��"V&�,D_9?�=@�9��8������dh���ɀ1g>s��
�o)�9�0��
��2�����a�s�P6�,t��\g`�Gpj����?�B,��7����K��x'72�Z={�y������5����3d�M�}�c%�q��ĩ���,���dC׶.ɬ��}Þ��� <���b�u��ɬ�Y���	�~��V���1{q$}0��
��ߗ�@�@�BhN���V��9B�1j(�o�f(E��>Qjϋ�<�/���ok���DE�-�rl�%�{���q��`^��� ;Οn
��n#�ՉX��� v|�/Aن���(y��7�]{�� ���w���|��m�����	7�#�m^�[�X~�d2���v椝����X����F��<��}�!�( t�#�z�N=,��Ӯn������ϲ���#���-��Z2�v�ͼ��!��H����GiaF�ي��%��2��G�����9�4��L;?+��X�e �,��_�b q���%~E`�b��hKgw4.�S�FU��J'ˠ),� q�bbiU^c�@�R�|��e(��~X�#5�+_�궩�ё+����G��R;;�%����g����S��9�������z�Ħ
[R�=؂�]�Xf�ŗu{��QΎ9jc	���2���cnQ@����ڀ�㫫��Ebj����!���US��.p��ss����+��u�H��K|�^w���O�@����*!��q�R�v��f�m��������[�u�j^���}~�;����;	p�N�v���D@�W��њo����H�O�ʏ�`���r�j���]��%�t|_�7���v�=I��M/��K�x�ݢ␮�7�]�{ĬL��ڙ���d+��p�1��k�ѩ���� ]��y�+&Ś�"�f	�2�׹�x�aшӺ4%�mc��v�#��b7������ݸ�"mێ�4:`�N���)��e.6��G���
e��	_'�M�Ry��7�"��=ʆ��,E�Ic�쉴b�)�Ю�V�-Mx��0�o��o8����$ȡ���(7��sxLjR���Q���!O6�}��;�ˁ��B��]����\�.!�`�q�E>�|eM�|�-{/L6J��/�ށ�z��\+��$������ӥ�?S�\����Ą��f�N)7a!.-�_I�2�Ї!\�H���i>m��Q0�8����+�(��6�RS�?��@�U�r^9�k�l�
��8
F���7:a)�z�%_j���:�$-�Z��$��\{�����О@P�:�Z�)���q�Tt^l�w'��k�~�h�w�b	��z�.O�˂����x�"�7�������GY(��M�7�T�y9��v��y]�T2�w'�,�us�M�cV\�:���ًY���li8��M��	A���&9`�x�<�[��ٿ$QŃ���暈��:�Y�/�Q"�.wġ��n��!�g�/.N3�J���q�y��%�����QR�(�շ7U���ܵ?ՠv�c�!���fa9GSm�Ke-����ŵ�����'A71ޫ4�t.���K4k��>�C�ϴ#��	��5�E.�m~6,N���ۖ.1G���o#�ӦL �����=�m�[U��=��*ur#���{s�y�Gd.n*�r��d?o�銝�%�d��m(vd,��" ��'K��Tm�p�x跗��2���Y���|�6N�m G��o���{��_�{Ae9H�Hn��]-R�Ӕ}ӾÑ{�;(���%�v�]�]^D�������A��Ž&�g?#]�Chʈ�>�� `;}/��j�<��)!���� k��y��Ή��KD`UB��?J��Ve��RևfH8~��6���96�9�1{`6Nw�.#oɔ��� d�Ff��U?�~j����
�y
�IW�8���$�Bss��K3b��断e��"��H�OоX-).YQ�W��&��d��;_6Lb�R�lm�|� �)</�}N��� ��ט-��B�#��������a����Y�|�f�.p��#���1�@��������	d��i$u����y)��{Ccx��c�,Z�c�+S7�5^CO��:�B݆xz��&�6��,�=����[xz�Z�a�=�1�ԙ{y&VnӌlLi/�V\O)�{+�$fR���J��ë�̈�<l8���\x��C�"�ګ��Ķ|�ݬD��9�w����~-�m��gC�־��ٳ�j
�$�g�v?�����U���L�`�O��������Au�U���/2�9���y�S�	�7��������9�iUb�/�({��V�O=?I+�����}��M�J*ݖ�#������n���c��9�`:��6��=�
��{R���J�8π�[5
��h���{�7^��Fv�-�6m�i����<��|�t�|	��߳>-��&F.☌���퍟�_�7C�D��`��AT�
���@�*�kad�qE#���Y��a � �Io�ji��1i/�q�wDɕ�C��B�����y�����;|�F������\s�����i�]�o7Zx!��;�2,?�/���(���>,X����k�3�)5/�^-p����J�������ZDxN�[��PSY�6����d�v�rs�SZ�0�+/��Pq7��!�� ����S�����'�F�/�Ѳ�Q�gvye뼨[[bR��CD����� 5.$|�:���j�>\�'������!����/]�fjv!�&�>�\���\�v,�m� f�N�tu�>�"�t���g���͛�W�e�s�ގ���y�Us	X������$/.7�s���UO�&>z����6�B&DP:�l ���⢁6i8�,�C��1�3���x,Ϗ��h�mGCL�vm	';����9/)�0r�gh^9�L��z����phv��`�����&��E����c�V4��s����$�Db��/F��D�"l�$����ը�Yg�N"]zO؅���y�ض}��� �H1S8��yv�ou����Ep��^�]ň+~x�ȸ����S�� ���OX��\����)��٣}!����r���b�@!W�����Q..��G1�K�\"��[�<1B��T��2V���*��P\��� H�1� E�j�Hӯ���UG3���̌��E4�o~)���t)i.���G%Cҹ�����<�ߞ!3�x��Z�Y",5�I�;Rf�6!��+2�M7���6�-���	��lr~#* 1D��8n���]� ~Z�������Xxj�\p��x�Q��Yv�����XU��	`p>������x�c��Wр��T��I�e����[���@$i�8�`Kad�Wu�aFv�H@ݯX��1��y������=�$��\ރ�ݬ8���;��@4A��$6�q�D���0=��e$ؘ��-�9}@S�����s�T�x�,a4mm����Ƈ��8���\�,SfXZ�-m��oOBJ���I�\v*-m��w��
����"��0Y�� -.�n�ct.YI�s�w=��,�Z���*��p���X�ŕeA�I��Lh*�?߇!��l��ʶ����K�DT�B�GR��E� $5A�l��!���)�f2r��J�@4>�o����.2Vȳ��(�:z[`���
>b���,t�¨����vm�F� q���|_D�*�L,����/�AH�Ζ�k��}-�sޚT��rl2�+m�o�����#YP�Rؠ6=�
��HǗSh�w�oF/���bX#N�VYѿ%�C\h���6�u��Lj���5��i,�w����,-�DoҲ�n<k*=�u��-��U3?K�Yן��G�E�cz�r��;)�U�չ\�^�������v��<��KmZ$]�#.@<V��n0aoR�&��w�|���beԼ8�$�=d �|!Z�N���P3f�A�ZRl�K�G϶ʧ�SܢYv�'�6i�y�=M?��+�{X�ԁiZ:7MH+\��V�Ջ席��J��;�$u��|�S�p��JW����F�d�&�SR�`� �*ٝ��i�}� ��榃��҆�Ǉ � R�j$��i�h�7��ȷ �;4�{�2�4Jz��ng��6�t��FН�|��w���^�����{�tε����VJ*ޫA�S�>�����PWx�N�0J񜥄]BR;���c�y�3�G�� ���{���z�Y�?��ҟ�iȤe�47p1 ��Ope('o������� o�=��!M�X��i(R��$����Ñ�y˼�h`X����] �6����؇&0|J�#�L�b��C>jd��Z��X�R���i��l�t��!s���y��˸�ǲ+�8ת;Qe�^a�X��>�r����µv�EM���{%V8���b-,�E_fƄ6S�͟���eN��[��?1���^���sB;��>l������H��e3[�ސ?��泌	��<kO��~��A:K8�l���a�.)K�՞�q]WJ�"��?!����Ì��4xK����?��uU�v\�sw�Q%�j�U��htj&��߀Z'lDN���������z_���,1�Ĝ
���%>nW�xY�"�(Ƚ��E'i�2ن�TЃ��2�pe�~��@ql�=oͱ��(a�8�@�8�@kF���� ��m�.ЬR���	_�%h�u$3�"N���kB'��Я���wk�A�̎;굛�X�j_����y���1S��.|a�آ�c�R@��¶����1�~��H�7K�=���.\�mW��	�W�(���G�G�����L�*�v��_`oR;�*U�◸�Sn��TZ�iI[��5����<�F.��wԬ{�6�A�"ޙ��;ep#�b��2B���f������U�A��xMmy�}M��ZMrC�~�I&k�Hx54C;�i"̶��]�`�]�X�����"��/#�Vh?G*���������?$|���k˔��@�U�,��J�.��-DtP��SZ������qeiF'p b��N����pg)�nI�hݚ�|�{�/�Th���b���T$��r}�s-��i��Uk���p�TUeAQA���_�/uO�4Ur��g
;�
(��!�X�]a�SqƑWJ����
�ݿF�tv&��3C�l��H�'��*eНZx�Ū��㙹��J���1�ާA�G��ʹ�
-P�[�覃����{8���_���c�)6����]/�q�WN��zD.���e<t�j+E`�0���rg�'��{{y�Ly�u&Z�ǧnG"+b�d�R(���m�j�Av�Զ���kS��O�a������ӯ�>�=�kZԂq���C"D���}�xD������B��Ǆ��x~6�-���f�3c���o��7O�9Rq��]m�7��j,�A��0	E�1RM&��ꃑ5`�dxo%S^���:�s��2��4'��F�=!�	h��-��c )|��	e �B�$��y��+�0�q��~�@�ɸP�0���~�!��4,���f�����W��(�^X�.nH��UA����+��̰���8���*�d��+�wB�_����]������O���Ÿ����f����FϦ~��>.̀�āah��7��/������x	�&���y��If���;!;�'�dG�e�7�w�6���5R�:��:d����`p'�(�QNQ���)��Z)��3x���� �g	�\�b��oV�d�o�F�w��<�`/�)Z$�l�4�D4�\�#6�ڀ�W�m�YA�|��vS����Z"�2.U`���
bU򌼊����rR"�Z#����A]�+�g��X���0�R'D3��#��p�޵�T1�L66ݵ�hS�	?�evd�(�]�dH���Rm`_g����/+C���V��U:�Y-�1L��!Ő�?Hz��d��������7��Dz*%5��XK�sغ�|�
�Y�5	�7\�s�k�F*Y�-�gaa%��qK��V43�9M��Z#�.���������oc����b��
D�!�cN�X�q���L��z��&���o�Z�~��4e�냎���V#��7S
n|�&,��OÔpa��L'"�Z��*D����>��_ ��wG��x��ݯ&��7�w��y�	M�&e*�?��I/{�jV�qL��f�Յ�s��:��(FQ9\�z��4�4�� &D��`}Z�7J�rؼJ�.�xs� �jE�����_���_}w�G��O(m�B/�����|��U����r��˲*��m����#BP8i�#�횇�;.!�tXE���6�����j��g��^-	OX�ƽ����v�nk���Zo?�ۭi ��ec� qR ���i��ԕjH"�c4�m���˲H�گtB޹k�@D��dm�c�S�k���;��E3
%��˄��~=�ס�Z}��)n#a�/����He��o��V��@8�Y 4n�|��D!��t4^�p�"zK��s�'�	��*,4�[���c�n������iT�+�4�éŸ���*AY��s6N��;0�1yVw�?+	��^ʡ�Az-����g'�����,�)���EM�>?+�R�Դ�@��5y���fjj��|�M+���o�.?��5�&�!�r�97Ly���>D��W��(�a��f�l9�-�6�Dm�hT({�
����-|�
���lcQ^ �!c�4:w���Xetڠ���iO�$�֬-֋��7!0X�Q&[F�z�����d�a�;fdHJ=�Q���ؒ*y�w��'/�8l�r���~���cC�-j��?ۧ��{r��8�(��l�g�g�8�¯�J������o7����n�\TV�}�|�m�n ]Mɹn��G؝w�*��"�C��6YT��qV����c�!3��;�
iD_6���H���([b��|$��ڤ���������j��o��X>�n6'�p��!��#�����4~uGǩ�(��r�i��Ȭ=�㺵i�	�Q�_�KN����J6/i���5%s�d��I��^Wl&�%��@q(�=3}-$Ty>���0����]t�L��U}�˝h�d��}o�NQ����3qX;�P����s��T�n$ݡ'�Z�X�S���9`�C��z���L�.	�k%w���:���ʑ�7��^c�* ��,��^x��1'�^�n���%̊���
)������K�as�Y	>~H��W�d�q��}���8P�U�* ����20�Ȫ�M��u^�+�3pR4��jdƯGG�0�Nakv���֢�����mp�y���^C�#�K�o�v�|HV��k���łoć��۟����5�o�>(�Y���X�Ҵ2Ͱ��b���\�؟��(+��,�QE�8��B 8�m`rq������ŧ���nV���ǅ��ccϖ�����%�&�@Jp�y��_����nOڤꅻ1%^�?���N-�̄��Xte���p�Ɣ�{ı�Gk�L��j�~�brw$RS�\�Y��e�M��x�[f��B�f�z'O�(J���"w���E�FÖ��RѼү�jmZ$V�Ã(���}����λ�J����s����k$$�95Cc�7��Ί��L6��
��;Å<��nXX�����m�h��x�Bs�c5D���}^�d�teBc�i,��f�ǁXc��Y�P�.��ӭ.�R�T3��y�>߅t;0:`��G�K`[iZ���)K#捥�)e��Y�&�U�8�8^�� `���V�W}J���Ӗ1��JK�>$��Gj��6@k��vwG�F�m���=$fC}��|��{"�A�}�wA�<������]~/����J�@H�2���s/,�T�<�̮=�9�d_瀶ڼ�o>�"}ח�[�d2���[��/LݖR^�#�������H�7�J�8��<���YWR(9�L����N<��ɀ�]�	BI�����Zw��/Bt`��gs�Ǿ\R/\u9��'�I��L%��AHMO����}�����	����:
K�Ǒ�hN�'�hK��,�a"J(�"�`Q"B%�?~�c���|�fj�1��6wTX�
7'+�F��<0�
b�OFw��=��19�;@�ý<_�"3���c�n��D�*ZY{r��?��v8�����\�"j
��v3zc.?�U�F�ϗ�������S��&���3�5��J9���,��K	��t�:��#����/ ���'���a�S=��BY #j�3Z�MYm��������qt�:�� �7 V[������!�J�@�c�����P�!lU���VϠ"U�ټ�k%zV��z�J�r�i�����TKnT�y22�5��ai���geL�1��<Zj:n 
�#�Oj�.�f���.�6<�E���[�`-��;�[�H�?5�"��#9�����%���=����6�����r&
d������w�-��@���R�oxZ�)�,��t�����rFd!��E�4zȘ���S��������ߤ�֌n�,0�Q2�®I�Ա|WdR��8M�4L��TkA=��*��IڒD菀4nej��Hg{
i����
ޞ|�nF��s�kH�@�j�$����?�bu��@�	�D2�,��4���t������� 2�%e��m��a��76>fޭQV��L�h��Y	���e��bf#��;[�b�?\-I�'���&�������ctڝh[�
ߚ�p�;8xr)%(tJK/��i���iOv�EN5�?j)yڤ@��_�2l�wj6%G;-�I�0W-�T�h85�u��W��g�BA�K[��N�4��{Ҁ��ޠ�ZMד��Q	�]��	(<5Le�HGڧ�+eC���f�-�ؖ���)�,��;�����%��J���T�sS�Bm�rb��	��d0��##.fw��
d��4����h�T��f�Dh͓�He58�pct��Wo!�	�����*s�E�u����V~�#ϊ����i�H6{V��I&씙u�ùvhlL\�,��QsW�XN�8Wa��k,��*�:�W=됇�a~~��Z�'���_[� q;�8�୲	����wj�Ik檃��7����h'��_٫�cp�=:�)u	'K��v(f�L�X�hf�nE�j��E���mE���u}���N��������C��x[��V:5�N�3�s-��JP�YR��1���yK�n�l�@վя�2脕o9pU���P�UB&�5���u���#"���[���+���K�{���bR�8L�Z�9���(+�ABwfw��sC�Y���5i��1�:��������_����	c�<_�Ld$#;8�yS����L开
�Y^����@�B�����ˬ���z��ah�4�}'<^p��bz��3�=�!���׸�<3\׳<�(�GXɝ�*;�s3���x���*���н����͍��HQ<V����/N��_JO7�i�ig�l&��6�Y����u6��j=���
󟌾;[:�I�j ��v��KD3�3`�
�9�\�CrČ�B���.�E��X ��ωD��e0^2YxHvﯛ�x�Ɠ�@~8)���ؕ�}�<��傦�^��V.,Z'��ym:UM��X��E�d��P����ﰇ���ho�G�#�q�e�Υ�_6#�D8!���ʯ�TmX�OM�[��jmH�2����y������=-�[��@�g*�-/�$F�N�	)|��kk&� ^S����d�єx�-�߶v��R�Ե��c�g3�VV}�j�5�,�.�W�,�l7]� n$X�E����X�Q��$�ODvc���>���eF��E\ִ�ѥgxÕ���\��4�Mv�_6ނ�%U�ZE�2���3�mߙ9p�� 򯎘�[,�u=�	�W[�lB���9oN���ku��]=���q��͜~g඄���Ѡ�s/�!rA�R�g�jrf�����c��U�eLj'��X�$%��}aH��z`�Dr�d�-��^O���M@4�LLm�6m�����_T���1'xF@�����qd�!��o���~0��&{ӌ�8�O�}ٱW��K�����=��J�����M$�#8�*�a6*b�Q�e� �Y���_�O_E;���,���Z'�:�}�^U�֌�� fX�����V������t'aL^�2߂��~�m�d�4��tO��y�q�����e�N����#GD Ir���O�%g[�E�kǔ�5����%z�M��@���_ט�CA)�X��xj�	�C���^� ���ٯ��V�uQhsǃ�aD���>	��Htv�% ���X7����6�E׶�f��\o��65POy��}��w������=q�ͱ��_��3?�9)&P$~|��M�0����̡�6�%� @��m��ki68o:��䇝��ֶ�X�A���Y:avN�Pc&HC�,��mV��\��ɟ!�o����l����n�+)�ő���nLM �o\D�w�E@���:!w�)��M�*ໝm'�h5��I�/@숼��SL5H�`׳���d��P>0�_����!|
����f�KXX�{�ɨ)E��ɽ(5���Ƶ���w9^z���k�9q�$J����5��T[$t�Y ;}�#qy=�D�~97k���U�m���'��!�������E{�1Ox��Ub��i��0�֟ ���6��ˣ�Q�4��H(��c5'<s�q.��.����W)��HE��i~D�:+d���w����^`�j��Z�:9�:U\HQ��笄9�Vv*�e{���`Z��	�"*��A�zP��wSK��������y����LG����
�&��&ܚv{��_�����K�6���iO/(�>�n$��{i������GV᳗�pܔ1�_�S0�B6g�04�>���g����*]O���xH	�Aa��:�y�7$&� �v+�2;iN����~��Z.�S �כķ4�=iʙ��9*�w��XX'w�?���#"�@	�(��6���у}Itb�2�����L�F}�@f;��F/LP��+�J~�\�z&��0G�;@μ6��]?�9�$m$���I�<���X���ˆI#���C���m��;��_6�������v!~	�:N	*Y}��ዴG�({�#.%;i�����jBWZ)�uӞQȊ��^jǣ��J8�"�Y_��"&�3m��/llKޝ����re�I�22X���m��2�b�Z�x~���=�N�� ���~���Hv�+���39�n��6pJ0�12%��_�+<z���K��Fp��|0��|S��v���8z�y�7S������R'yi�%�i}� &��������?5>Z����q����jujIZ�,�N�L6w�>�����,ǅb&TJx�)0��W'�q�>�q���y��������B>�.���	gꎤf?<Ɩ?�i��/� b~+�������N������w,������4��/q"�,^{�ͅ齡�S[�u���=�5�H��0$2��6ߋ
m$ˠA�@�gvކ����Q#u�M��s��L:_I�
��R�e�������ct&�P-����c4(�G���3���Q�~/�+��g� /i!��a\�-�1����G���RH9ݓy�#@�q*/d���u��hyNP#�b��
l����<6�6"v�0#HFЎ��m�6��d���RJ+�e(2��ۗN��O9�V ȕ�>g"V�s���{[���j�b�З��9�y=����z�8���7r�A�B!������4"p�2l�(Ν���v��1nU{kgh@\������S�\P�����x��p��܋���Є^�{6\�J��؍��ʥ��9$��z����T�F�%��\��J��RO�R?7��̄���c�(�%b��x����cv��yE���]�%���5F��*�;���#��w�F���3)��jį��9��k�*"ϋ�W{�%�}�6��]�]Fj�l���-��-�\�Ȝ�i�4*~�瞲1�j�|�m���Ź�u7�%��ܩ�* lVn.�29�R������?�+x�D� �8���\�9��a+9��t�2gr�p)焵l껮��Uٷ��f?D��Z����"0곔��_������P)-U��5��F��X�`�{�B:nB���,I�,;��h ����Th@�1���'�J~��_
��^C���5�R>�AdH�X|�f�w%Y~�Q�ф�b�o�EEX��0C�����8r�Q�s���ؠ��
�|z���~����fÅ�H�y8o4h��ߥ�o��k�[��1�6�"!̼�ɤ(��(Hs�Ԩ���Ӝ\�F�1�)�=Ծr������e����{엦+���m�V��ͣ��_Q�F���]��!c9�_��kg�����O��g�+Ӑ��@�7�*��D۷E�r�*+4%C�_��ѥ;��*�<$��P��� ���8�W��Ɏ4�߄���\[�Af��c����q��n��A6�U�������	O��P��]0���<��N�(�,����aj�D~��9Y݃i�}rP��W�)z�e��D�Il�P�����C�U��Qpȅ�-�_KP�l�g��\xMA�&�	�	�a۰����x�Ԕ[껾Z��ߵP�v̂��n	D���q�Eyl�i�z�z���m�F�DR�	���/d���w�d&cMx���!Zq@��:�3ȟ�l$\'( j/�
��*U�-�_V�_��-���wYꌱSiS��.4M���3Z��]!���	�z�b���>����Ϋ�&{W�:F)p�b��"�ԥ���k��.����k���z,���� ��7A1�~�V�D�$��10{��*�u'�����X������짿�
��L'�bٿ��iH�^z8�!����,�2~%Z��n�uz�� �)����������#�9T+Ԟ�v���TԶ!���0�;��G���N�u8��t��Dq]�����@�F�/�$U|��� �E��%N��v��c��D��U�����U���5X��O��II@	�|z�CW�G��h`�Q�z�$�̜�p���H�U�ߪ���zJޙ-q���_k�rݩɦz�
�M�8 ��]�T �`.�[X(ϩ���댒Tv�di� @(�*���(L����B��Ż�*0ߥ�^
���~V�QS��Y3�h�q�O�-��>Ǧ
 ]��%� ��Wv���m�!���nQwc���)K�<�����t���a��>����D7�z�����G���B�Q�S�y�04��h�M�n!�i:?FI��
���^�4��o&��Y"s�p�XW#TR�A���`�\�ë���
�l�~r&�!p=�]')߽uJ����g��+��ld�>��#�E)|D ����^���z Qi�_��#��g��ؾB{�Ya�X�^���Z�<�ؕ��3խ6��]k#Q��IR{��r�M{�J��]X�nˍ�(j0����w��/G%��:�QY��F��Ypg�?AF����p��v�8��]%��ZAo7ĖXr�\%��Z�Ǽ�U�Fn�� Ծ�
x�r�}l�޿�H�����XO��d��P��#���
�P�ۥ�e�Q����r�c���y�Nڙ�<m��f���"*�噬�D�qzMp�|Osa�a��`�B�0� H�T$hs��J�� Z�Hb�Zin�
ߍk�|���c�9�(�;C�N�R��4�*�O���-mZg� �}'��ޱp�ݾ��sR���vE�3K�%�L�w{a?���6t�p�����@"�I�W�qP�?l�-�R{#i���䲀�P���4����ֺ	:��mF�w�ւ���R����'Vg��R�����"�"+J{�P,(a�;�	x��B�-%�������A��e.�� J�j��l�Ȑ���71J��Y�������h)��2#�]Eu��O�]��0fY�,*������6`����zJ��nE)dLbெ����'��2.���o�_��Y�Ͱ��/��8�
��h����Kp���\��I��� �
�I�	�n����e0j�g��� �Y��Ў��X�μK&���h��t?�#?p���������(NdH���������ذ���L���3��ET�yD|�zs��6�rv�H�bm�ڴ}�Y)��	�ς���	���D��;����bƔN�'j_1��nk�Mg9�X-�[p�/q#e��`�WolSѠ�2� ���L��h��x
B,�J$P�ybF��d��Q<�B0��j�8�{�c*z��K\�S�F�82O��g&�����.I�^NoϱR�` �SQ(��~դ8����\��i��9�_����i��!���?�o��J=B����y�v��갸�t�&��23W�� ]�F�b��{�)l�xAh�t��Z�T��U0�V)||ԧq[M�h��̎��2tBO����i�ut(k6!1�8�'�	����_�'OLڶ�o���N�F!�<F���l7^�^/�de��N2�d5���k�`l_%�J'V���6�
ۅ�ɸ���҅id��S�a�ȗ~G�����Fw�fC�eyK�Z�#Qљ���k��X���=v����CWP{3Fp�k��d����q���_d�_f��LN|l��N�-&���I%�/W�� a�Rډ#���������n�� $�w�TS8�z�]�Yoo�P ��'B��ō+xoc	􉂎G���iW=O�ܙ9�NZ���pP�]>Ô& �E�EL|�
ښ�v^gU4KDK,�d��p�?������yr��*���M-�� gum067D�v�gbܗ��m�_
�lI"צn��왢j^�������^�GG
���ֻ1q��/������)��{A��{N����5�����V��T=��<����*P;�A��8Z���O��K9!���h7���=�ղ���L�������ӶL!<���3�g}��n���-��S����eg �1
t�l
l09��
Ց�>R��JĒy�y��c�"���Ϸ?�r��T����(�2ٳ�+o,�A���ō���h��%���:�����yH�q
��y�{s�#L�Y+uc���r~*pC���h��!]���"DF��� �!͚N�u-⣼&�f)��`F��q��U+EP����o�~��:���B�y�M��YU�Ip��:8ղ�g?�,��Y�lW[���J	������_�(^s�P	L��3;���| el�� X�*��oW�(���*𓌂���>Ԑϟ��p�]��_g]��y+p�#d%��ĝ���^��6�ߔ���53�d��xn����'��dN�����=�t�h����e�m6,���g	}��
� �O9�dX]����E�ˮ36o��`nj�E�@}�����0x��_ao˧�g
�	���h!D�.(Ic�-$\9T�Շz�c(G=8��/!=�f�$�h5 fC�_��7����{hg8(j�7�5@�A�f�^�-Wu�D�sLȓy�N'�Y��9�_i@h��+�L�9�w�7��ʜ�N�҄�<$-��jH������G�K���yJ����̭�+N�E�z���[�D(�PS��Z����4��t)��#R��t�	�M �ۛ�����(��e�JG¸�֜өd#1f;�/]'���w�l0>f_viU�������d��9Q�{P��/�7�C�j7����`��UPq�ے'�Ù�ym��:A��4@�ܭ/���O���+%�I1.�R\Q؝��,�h�
opZ�z���e�Tc%x�n��!�+��=*��׬
�I�%�T�rb�o~$>��-�c�{fr~kx4j�|��t�jc��c�ZgG�L�$>4��k� ����~D�?oC�i�}^�H]��7�6��v����Rzzm��\A�Js��o�°��|>8܆�pZU�%7�$��B����<��$���~	h�[���Ճ�0�эN4�A��XpqQ}�+{�#�:�_�g5]�a�8k�Fǋ�y�jIrN�Qg���r@��W
΅�kr�P�{�@��c/�A��(�ϻ6п��Ys6�u����I>�1�K�E�8\�.b���Ӭ���zb���߹��M�3f���S�+��n2�P���ݥ��+�m�#��V�Ur~�����GQ�0���'	I�ZHW�-���:;�Du���-`�r^�j��#Eh+cf�����?������/�����A��kI�N�+<�:�]�� �	D�{�J=�w�Ld��d����
Ü�ij
�Q��Հ�G�AO�i�p  r^�Xi� �4�����~�8��M�ɍ�-I�]���+��5��
 0��Z#���?�P�~��ω��߶+�����j�脔�	��=��d����$�]<3X�ұI� ��<'��e�U�nWK�����T}ʌ��w���\�VJ� rO�Y�+NL��xs���0��"�{]*i���;V04�f�k:ֺ2��"{�kQdU�1�G����>]�.ۥ�%/d	̈x��I����>P[�u��\�l�k"����m,x{���ϝ�WJ�<�G�K94�O`��d��������0P� �F�q,2��^�d����yq�#C�;��@�)##�����2�fդ\e.&��+U�{�|k��hM]��I�^Ǟ���h�v�x�r��r�x��|Z����d��a���?�Vֶ���:���4�}�g���y������Ā���&�s��JF�9��̜�C�l"{���-A��i�U-dg����^���
sѾ��.�� �_�V�Q����E[�N ��-�;HP��0��L	�~��2�@6��ŕ�5v ]j)��4ߟ���M((��l���x���HL���^7�4y��`}so�B�.>6:�䛙JZ�
�9�No4����i��
��ю�����W��Pٟa}�t�F��--�����U�Q��.�%I8��k��X�'��G��QF�v��$�;WqO҃ �iQ�i�,n��d�n�S6ś���k!��8{�|O��0l��x����󷆌���	�S� ,���Tn9�{�!{Ũ���c��'�G%I��@���t��%3N#/ �ֽ�w���K�
�ݞː�19[�i�kd7����N3� +nE�fQ�8o�c�^��$�9d�a�9��4#�����䋾�sNQůT�W<���D缌�f+��L�ZI�[GAO�~�j���U8��Xx�g������t��N¹m�J4�,(Oh�3�����9�˂��{�B�A!����T���t�:(ʷ�)z��E�Z��~]x$�)s��L���Z�Ezf�yޏ�M�r/� E���s���2}�W��D?/M.�5��Щ�^�~��g�%Ls�B�s�)�8O�m=��.M�3@�p�~�sگMQ��v����C�0�J����|��#�O|�_�)y>i
�J��^ŪKJ�-��	@��bg��d���[�L�T��~(�I&�B?5��Q��d�Z4�e�ёg=�kt.<�O^J�#��ˠ�W�j�x>pxr ��]�Z�O^��)H�_�/]��oޝ�x��_�v������ݪԿlDA��B5o*�l�,)�.�&=e����+��A��X6=��s��՝0�vs�H8�j��wk�3F���0Zy�0oNs�w�:�TAa�4���eg�:܃�s�K}SxTt1�g�๵QuM�&[(�-��Qy	>m�-\���6%���ӌ~��/�̟�U���l���c��k�Hd��f�c�>����퇡}*q�����w#2H�;����˅h�!�b�?&e��'�P�{��A��h��^)��g+7�m\Q o���S���-�P�=�	��o׻x�}wl�����X�Hد�P��w��bJ#UO���6��}p\ f�۽B�.�I�ް�K�L�*6�/�ǣ6Q�PK ��`\o��@����P�8Aj��<C��SZ��U��)�I�<x`G(��(X��<�ơ��ۻ]t|c9Y1��7G��teK�e�4��`�|H�@wZ�u��͎I��f�mƽ�X �*��Ba����MJb�=ݻ�U��K.}j�h��f���~�AGi}��^�}�6��3I�S�L
ϯ�2���f���M���4��(�ȹ���fY���F}/uI��8)����%���5����P/��
��a�$"�bdF�7�;;���"�a���\Nr�J;0լ��H���Q	�M��T<���4�b�'-.ݭ��PU����d�`��Ǖ����hNw�x[�%�Q����ÿӏ�R�Mg��?]��d|ѹ$�����4�)�
�I�m�6�PA� �Ԋ�z�[����o�RDc=	$��p4Yr��z�o*�dD�/�T��3��ϧ�׭=�[	(�l�۾�ܾ�D3V�ѿm��d^9Cj������81FI�����s>������KU�SO2��qkt�t���nB@Ej�x�2��6(�'�4֊�@U��p�7n��(R)]���
���bFJ�H�*;c|���j5��1A&�l�d� �)ŵa�h��"+N��:�|���b���:��ʔm��j�K�
3�TT@6V��u_T����>�C�A;n'�r�.�-Q�������i|��]���ϙ�=�������ƓZP9*ܳ@{��>!��z7���7`����g�P��+^�����Z��^(�H�BNP�k������EWM*|�O����Č�f䢡�4�Y��'�I�G��O}v�.��F�^.f��1UԴ?���4b�fP)\��3�aF�]�}��7�%�W:Ȏ�~[���+�e� #j��^�D� �0��^Wa)�v,rB�hn�s?�w��pq�<���6u�T�d���`%ކ/3�%#Sj�q�I�8�2��^��k��2E%h�B�DP"O���)�޵%��A�,��y�����3�1\аƺK%�'����*.-$Zw'�
���Wk�P�}�=�J�W��#Ԑ��g$�<����>�V:�����SߐV�W^4iC-n��,Z:8�?FzU+�u�T_�H/�Ş/�U4�_G��"�W��DNQ��oD�'��|�;�ѽ�$16�F�D��
;!faB���!�\�?����p{���K�Ul����ߥ���ň�d�̩�u��8^���K�n�6 �ZT�{����9�R��"y�2S�j�w
����W�K�J>���e�\����`�._rp�E��|S��1��M���b$^5n�=z`�q�����k>K�$���V�սE(O�S��]r`�j�ǲUf)��<:ۇ�.ϥ����Ar���6d��E� g���%�)ckW��Ԃ_�� ���m����6*���u	ږ�e�ѳe�S�S�¬��qW�I���r���p�ѡ��2���.ٞ�]�����V�����J+bv7���d�+_0�&�����l.���u�y���Na�u�:l�TcA�g��$�wr�gR�Iy�QL��=0��U<
�H��-X��%� �v�[\�ʪ/=v�Yt����_n��f%�-��U������D��+���?ZӚ�z���~��'�c��W'��#Ɗ���z��Guz5�4y2P�۰��E���vΰrV2{1�}�3h�u��H�F'��bJ�8ljl�Ә�:�A~o��{\8�>�9s���ļ1��P��x.��k�5UB3I4�u��1z�&v56�M�Md����H�8q��9ޔ��)�Gd�j�I�>sO��paz@�D/Yg����P���K�Xדfs�NWV�W»g &�]F�:�~$F��_�,�� �s)�Y�3?Բ@�sFDS��֬_�%+�b�}��4���J
��\�F25p*�-�V�֎x�Ε뙜�v8o�+	�a�����\jd+ݦރ�=Y�S��-d8�Δ���O|[�%��	ϩ�:����_{\�̝
�����;��[��
�U�Bmd%W�o0�)9�U`&c>fk<Z�qL令�;D߰�#�>��E��0L�#%��Wu��il�	pԠu�g��3<b0@��7K�-#��VKA]�Ґ�H���=�`2��	Jd�\	��yd�V�WP��/#$�y!�5M9z�B�D+�r�a[Q��ĕ`���K؞�pXF5��&�RG1�j����P�Q��̛۬��8voifg�3���{S[��^Ӭ�=V���OoD��K�	�?&ZZo^�eA�`h��z�|
�T�`ԓ��D婏bڋHJ�3GskcM?4��7}�-�;rM+�%�9X���M��/�ۤÛla�\9!�}ńo��ƿU�ӌ�^=8&��cĬOi���3�I�=�bH��$�7�f�t-�c�w���|����!�'{+���V-
�:�6�ep���˺m�?i4�GM�����9��5S��K��b|Ok���~��({�=t^F�CJ��s�XS�#�E�6"�8t�=	�1T�-v��4)�Ty��o��� �"q�e
�|T>��?~��96���^{�u�t	*P��5+��$����e���:a���K�In�^����EvWi���7�I�e�w�.Y�l�0�8���3 �/#ot�1js�D�1�$l�t��e�O��	�9NfnΡ[H�xu)ݬ�z&OHoeF��̸;�yBy�������@I�F��O'�&7H;�����b�2�
���o��0���$�6���?Ȝz*���F��e3�h�juLBʻ�lm,��^��_�riXi �צ��؞�_�d�I�!d~L��y73����D�;s�7q�O~|tͤ��kRi�=�Mp7��YE��:�`/4C�D�������;+�"[���;�{P)�m���T�ϲF6�H.2q��í������Ad���g͖~*�H�y�����k���"I��0�	Kt+C�m��h;����I|�i4ͭ�)o�d�ԏ[$�Ng����n#`x��t4VÜ~7d��!!T�����?�I���y������X0�������
�/��M5�ⱻ\4BqT�� �`V��F��}TV�6�g��F�E���|���e���n�����I����-׊��։�Ȟ}�Y��@��H�r���P�M��x�hI�&*JJw;&� ]����S�6���Ԥ��8ש�(����W�]�|�S:�hHV�H8��k��p��wk$�3H����&N	-F��;�|7C��Y��*)���8�5��i�Y�X���ʀ�cE���7��-b��W��3ݣn����PVl��(	�.7`�O9~��}P``�ny�@~�����p7�6B��9��Q�l1�~�={{���ʹN� �_�XI�]�V#�B����h�@ep�G�hr��*��+���QҸ�r��G���m�n�1�����P��w�p6.?��3 �9��u�@
T7@�
~냑:Y],c��YrAF����a�M��b�WL�jڌ�IU�����<ݛ��T��&��J��l;�5�&h�l��݉��)�^�J(m+��|��I_�*�	���%�H�e�#���{$TK=f��m�L�s��������LfE��{jaK�n�Ը��0����sjR�<�7e|x����D]U�~t�)�SUiܐo�_ܑ"��bHH�bp�]ND�qG_"�U���3�ă��C�@�<����_!�� ^���_0;�����
r[�� ��{X{>˃������������\P3���nW�Eu،8��c�c�����]p�n_.b ����(�pH�x "}pS49��[����Q��_��J�%�)>�8��)�st�v���2��`H?�"o��*�Q� =��L�b׶,�
�v�g3� 	��ķ�=�½{�-9�S<`>N���`������E�Q�W�ս~���ÓԀa�0�X��\z��v�t|xUl)��L��(��ꐺ��y������X	��]f|�|�Ԛ��|&��dD��xԃ�kW���:�P'~[w#�Э:jΪ�82U8I��U?���~�f�V*���ۢҕ�G�+hM����ݬI\�f����9 "X�S��Z���îǟ6�s=�S�K������]�#�)����JG�9�y ��g�G��u T���x	+K�[r\�cVGi����vW
z6��4� A�3�����.n�ݷ eB9uVglzN�[�lne{���/���f��>R^V�f�{�g�wf�}���c��x_a�	Q�i&:��ܣ�υ�y����n|��: l���J�[ "ڀ�I�ظA�q�rFb�eP���]� �B%P�Һ��A���t�Q��$�U%A�K/�>���A�nY���H:�Ф����{���)��t�k8�u��yKN���v��_ ��\���$<�6����RHTqW%%rR��
{��پ�A�f�U��P<�IM�c�(ySC�_�}i��K[�i͎�O^��v�X���U�R~MD�j�>�g`���A����a�o<�����؆�[*f�Z�Z����h����0��z����G`��R~�%
�c�O�Sh��)C�U�SǂoV���]q�`�mI�J�n̈́D��؄H��Y����vt��!���|�QZ���o�����"�C����H��NH���k\nn��L�Ե6�b'�e�����J�s|�;��#�#��I\,�"Ӗ����<������~�%r�l��~f%�5�w3��ʎBo}���D�!���(=��
z�����g"�M��ņ �f�Q!���Me9��ct�3,����y°0��k�GL7િ�"f)�Mm	I�FÃ�~��2�jw�\�Ѩ
&���D^TN��Ngr,�h�n>����)��X��؇��K���~#���yid'*�3Y!`��uWUH�|�Ёk1TUݟ����^dȉ��3jJ�+����������l$˰*�i|˝ v%K@��D��jo8'���X攇C�݈�����1�-�{"Ƅ_�@���x��j���K\��J5c���fl�r�9vvkQ�^������h.V`ɚP	���V�~��G������S	�s|��J��K�ɝ�||�����
�#cS_�!�}R"QL�ǥ��D�!9)a����A����p�G�D=�