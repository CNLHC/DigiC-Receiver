��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ�����u��C���
ݚ�Unhi#|�4$�M���fV�R"���O��7!Ԩ�=u?�=:��}� 3�[]4O���ۻ���8�m ���=��&�X����I���{~T�}��t$ G�Qj��h�4����m���f�J�b���q  1�F% �)T;��-��!�xpC	��z>"1��!hpڤ%��EO���2Ei���Ii�N��\\�W��M=�����W��~��Р*g��MwS7|��1���:Z�LS����� ��gL��h��k��n-+ �!ub��2'���r����E5�h-K�:�e�� ��K���dP���e_`ϚVj�!�ڱg�k�%��U`��pU��,�Ҳ�?�����Z ��x:f�N��w&�.�8�fd@h�\7�V���떛��1�K��"�K�����[��ΖݣJ��Ƕ",r����EP�d~�B���'��Gv�rR�}�閞 �F����2���ej.=��ҿ⸔�9�M�h�>O#�E��� 6܀ږ�p��є��%&V�l.�����i-�f�u�z�����V�C�e�����#��F�t�,���oh�E�&�d�is�f�]vZ ep��^S��_
JF��+�m��
��ē0�2����׆� "��fU�g��\��t�(��%��S�)�<�Vؠö����w$�ə����T��Lxn�ӈ7��|Ǘb�C��1�+��3-�ZuFeO�}�$�|����E��l�)��5��4Ie�a4�f��;��7PPcb�}���P�>�[%b;f��P5r�5ؽ���k�t'�RQ�x`����z|�m�ܔ�n�Ql��h��[�(���f2圷��jsC>�����"��������,����/��*f�'IĦ��(�8�|P���e�ݦ�,�*n�9�N�GC8a7:�$-(	��8׹_џ�.���gý�ǜp��,^=b��͏,\R[�cR�pň#zJ�[��6�X?hg��>y��g��|�x�P�-S�~��&N6����)����l�z����eru������"���	�q��JE(�E$8�\� �7�Y�_}C���s/PP�%&�\��-x��S�j)�F�N:o�z��\��U\�v�&b�O�9S��5��ן#��F�b.u�u-0�Y�'a�������ɋ�@�$k�A��\�t�x�l���B������E���ݺ1�TQ˽Ő3�5w?�ܧ�9����K8���:<)�3��q!���Tz�[2��/������'��������Tg^ ��RӨ�|�^�ݑ1�C8��j�u�y�Lm8�BE"��m�#�-�P��碿Ĭ�l!n���o����}jrg��W�����/�U�lZ���3�tG�-�x"<�Ts�N�j�uQpRC��</ ��.,���c�� Z�]Pݐ�$(���E'\��ʏ�E��q��s�K �؆\}Ҏ�O�H>�~̧�Ұlv̨R��'\��6��a�d���$2�.Z��X��:X�È�1�)s��uD�ogm�ލ�#̤wPt�.�&Z�]��
w�"��S�cD�����AC��r�/�Fh+��Wv�LLU�h���&:��2Ɨ+4_���<����.daR�~-�
o5����܂��%�\}}�BWJTl�kߴ҇�9}��ii:�LW0�%�����`1֑1R�B:u�Hl�	��#ҏ�o?� s@�C��c��5�����f��ma<��O/~a�b�q�8���(u�Z�@�ص�����&�ƞ|�@�:+`w� ��oD��n�&�b�8yY^�O�,�8Մ'JSW�m�����.�"O��o��\�5��0{�8�@��I��	��W\,-�ᯡiB�e�#�_�>Y���>��	��^ȯu�W)?���'��nI	��-�ߴ��X T�Ŏש}�r�E!Пu ��=�_�a���/(g���pP�c�r.��D.�֐޻gw:� �th�WN���g	�������q��#�6���w>&�qz�c1�ri�\4E�4�Я"R����D&B��&k%��}㗣<қ6}Q��5ʊ�NU�8B�2Q}�8?ny��6E ���R��oF��?Fw�6x��肇����ŷ�����:���Ľ�¶�F>"��k�gYF�=�o\?"2	A;}��ܖMZBR�Z���J���j;�ؼA^���ߘn�T�Ǫ�'L�Dڡ�k��A+�	�r�\��ǽ�i�~mPW�)�m(�@��1�9hѰU{��-��~g<;�3Ê�9
��d��t�bD���
��x�X䭠0�p�\\K��af���n�i�}�&����)�i����N,�-)p�0}ҧl'��n�׽��B�O]����&��7��u��<q��h��ͥ� }��"} S��>�� ��)H܍�}7������A�.	c�q�u�];&�jM賓��8��Z�^;��H��4��A��O%�S���Ra���v�E_ޝ��Ugz��niW 4%�b���2��s������M���f���e�3�?�����dbҔ��8�i���x�[Ѵk)\ކ�5�l�DAM�r��˔�^%/a1V��3(�sJ"����q�m�����!;" ��?\�NEiF��ݏ�j�?hc�9�߸�.U��I���x�b?�����o�qe��Mu���Q�N@'����H[�஺<��s+j�_Z!�������z��M��I }j�X�5�矼5[CfY� ��;��C^,_5�E��)�����УI�c�2ּ*Nw�L��C�,j���o�V�o3C:��
`韘�|��^�`l�yܭxZ�g���$�}�U�d��$�P��-�^p�c�5�����%�k�s�!$����)��3>�w3���* �u�m67l�h+,���1k,p���H3�7f�L�BK)�"�z0����L�O�Մ�O�$\~���oD�H������u�1��F����T�����}093�����}�w��RP�d�(�����㶓Y��b�r+�����Q�̩��b_m���w%B혴:}s��iv��"��D��C�0��G��1��EX����B�w����N�J<�%���#r5B��r�����G,9� �:#X[�z�{�Ф�:D� ̩B�w~���'�p��4��+�ߘ��i|"�X�j| γ�uuK^ڛ۬����H�U@8\}�<�Sh~o/�'9��j���x<pp޵=�~;ej6�o㮟N��<� b��^�"����nY�ʒ $\���I�<��v�J�R��1��/}J�J���M������Y��E�H.S�r-�U�A��D�*xTeZTZ0�M����;�h/�[
*į%o٦'�>�_�}�O8����C����T��'A�k����yժ��d��h�0�l�of+����@haֳ�o�g���'�<k�`E(p� ���ndw����E��u<�Q�s3�o*' Ի��������Ǽ��w���=�o8���h����(zG��psBD��~p�\%$OJKj�4C�ѳ"�Y&����@M����s���G$���g����#�XL�G����fN�I�*O�ᜟl>�6�L�D�D�1I���**�	��B��Lwϳח�O��e���d�k���v��/�O5���a>[��~�UlƶGn��P���~]凶Uρڜ���E��%ܬ�\ӾɄGg�f���|Z��Ö���' ɢ�`M�~��>�97�7�Tw�������ڸb��~jc���dh'3�U|���'��q����܆��|qxj��%"��R)b)τ�!�uBuRW����Ƈjr��{8�)T6$�2ݝP��RfP�W��=��G�4U#Uِn��A�]�����G�?�n��=^^^����=^8E`�/��"Z��]hz8��7:DV[
��*�9���zR��R$7t���� R㯊��ZK/��81������$)�b��; �#�:��3n�w 3��*>��u��&��*�53�6(Xڠ�l�����`���]z�dK����JAy�t��T�#�qr��R)t�^F�U�?�ϯl@� Y�`{P�Sj�C��E;�.˺~ОPO���ߨ�{Z�(x�g?1�,�\Z��wCM#�z��j�M3�O���hG���3�W��Ù���K��Ȝ��v"́ZW��.	����(W3��!��͢�W|�)
��I�.m̖=9;G�`??1�@q�w�Բ�]}L��4�h&(������M�$��Q��4�*����A�)�^k�9H��/��h����ͭ�.�����T>��L+[<b��(�����#�߿yo�$X�L�b��գ��wdz�z�IJe��u$�Z�J:sd
�}�*g�=��zxF�FP��	�c��N$�j�a��LI���ҽ!�ni�����9�ο0�@���h ]�ɲc���"�>��S�(�͑��DR:Y��^Eu��~TѤ����\�#A��\Q��#Upѹ �.�4p'K� ����(8 �eގ>gx��䚏y?@�I9'g���[�6%���}f_�ż9��fp4&�:����Ë �Wm6_�L_��z�Y~�Dx��m�J��9�MN��,��H^ ���$�"�ղ�� ݤp@w��t2�i�Z�X;�52�� ��.�*���@�!�úA�����upe=��V��.}!���Gb����-KnW�H��?�(���DC�����
r�m=eq�j�Ue3 g./�Up�sI ¶��OZkq�]�-%6x�х����#Y�^���0�6�"d;����leD��_�)p908r<����EHo� ��Ҙ������qƷ��3K�ʖg�ā����v���ྲྀz�=ƽr�E����e�b� �\��s�YB[�.��j���>{-Fp+���$f�?�����ք��X�Ý��N?rA0�C疢�Z[�
�|mx'M��e!��f�j�ĺ�?��l����R<o�PJ����IWP�R�/[L6fCv��Gv

��y���8x�߯e�˩�w�;ZM�R���.R�ԘP��2�D�8C�m��U�:EAV^{���b	'CBw��iLxR�u���ٸ(IhI�P�ay8f�I�n�$O�=M�o�hJ΂D�˥Ֆ�sU�~@�]A�u��=�ͩJՔ��f��g���OX=�;��b�:�Ḋ1�Vp�}p��}ҚmrL�|��N5�OB�9I��l�{@�cʌP�%�.��&�6��A�6L�G:�������$.���/���oD^��u_� ����GЈ��+����&�b������&]�9:~g��#j��s����̪���*/��ٸ����9���^����r�����Xq�:��_{!Y����-Oz�۬�N{�~�Z��~�UȋӾ��#_
;�1MLJ�/��R�1p�����v#$,�<����xe���2'�Y�/�s0�2������6�A�A]k#��s+"�230J�H��$2��	]�\>%^L5���@�K�[$Ħ9E�}ɋ���Z����c�L�R�C�'1����y��u���y��u�|�]�D殱���g=�\yΝ�B��\�?@�\5G�r�58�CL����ɎG��v��T*�~!X:�fr�.El��p��	Qa����K|
�)q��	�I�j卯�0+���>���y��g��2w�p����4�[_\""��ٷ�'�ҷ�@�=�'F��-��;:��@�s5^V�w]K�53�������MxX&���D�e;�-x����2%�JM^7߷��G��d����q���M��3j�U�גØSo	��}�