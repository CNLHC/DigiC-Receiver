��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��.ܗ��z��3���.ŷ.>�g��p<���c_ �X`m���F)�Q�'(~�����	���Pw!�G�KP+t��(��L�p�E���l������WD�,~��D?^�I�ɱ�6`d��uSx~�}rX��Ͼ���wsx���jL���4s����	��Pz��Y���f���5���w%���C��g����G+��Щ"bJxdT Ň{p�Q���D��q�H�	�X���+ݳ:-�����YJ��=�{|�G����߼;�l^�Xf�W��h����F�p��;O�D�t�>v�!��K>>q>��.%����0g�Yg���(ph�%�yL�o�	���lJ䈒���nU$��=��QIG?�׶L}�ڷ�H�4�6k�M=��i��r���ˆ%��������oם�r����]��>0�9Ӑ���#�J��p����n���#h!�Cdn1.5�p�8C�b_�/��r�����=�b���|O��	��p���	��qC�d�����L����Vn��-_���W̰Ew�'��O��g�@緉��~y���}0a��+�?�J,�R���D8�C�� �&Oާ��v��D:dӁ=`l�l��C��-g��\*� $�y�/B�'���^��0̉Ű���d�̊�(�O�m������b6;Z���F��Չ�*"�:����p�kcY����r:��X���6'�dDڷh0�L�<��,�@a����\��:S�o��'/}�L�qm%p}z�!�/#fO⏔޽�v�.u� !p*"���=��T띗$'���%ƕ>X�RJ���a\U_�vj�s��Jce��ƨ>Ո�����E׍��;>S_l
�P��q� ���A�&&��Ƙ�,p�E8�ҋ%���h�2�H��M5���XE3f��e1Xtx͐Qj��]���W�3ጤ��ýwp���K:x6_)��m��5ܠ�%���9fj�T����Z?@�,������u�0����1r�)#IK-.c�$�)��}U�f|�A�y� *�c�����vV�q%@AV0��>t%��O`���
"�����̚G,�F����zmXm�訶�ls����J�Z̝��>�h�ȀiC�!ھ̂/1��h=���<_D,�Q/?GG*�<���Ճ ��!c��|��U"b\��x0Ԕl����a/�d�5�	[�y���ޑ-z�ԋ�J�u���+�f.y��>&8ײ�	,��L�h
$�%��C�_������ܽ7-�'��$2��r�%��s>�4o��L��8*%�z	��Bm��1k�D��w`�؏W*7����F\z��$s�1��A�w¤C��tuf�ޔ�����sp�i�fun=f9�zI�!Wk�K�@�?d�v��G�OJ��کV �@	�-�M��l.���>)�y��?� �~��K�}!R�]0OsM���;�˴ˑΗJ�MB�&�b������������=�JZ�\��Gd��Jk�,9���&�\�p�.GS�r����@"m��AN�h		���X\6k.�o� ���4�	�$|[�ؓG�b�.ۘ�I���I̤$簻��NI*�Q�y�`CY�e���Si	%)�z��p\t�1����1����� <ޑ�
��,�q�*&C,Apz�S|���(�Rr���F�_�pe�FY(J��-��(RM���j	��|��"M���=� �Y�:�#����\@�%���絻$S��a>G�xme�IDID�Gc��զ��lV��۾9�а6b�+G����ma�i=#&i���y�����\�}yy����~ '�p�ƞ�K?L�+i��p+S��y���\���Ԛ�▮U� 鵽k��>�)��s=ʎL��b��a�L#���("�] ��W�U�Y�βWa%�d��7 �0�G�ё�4.L��ѕ�)���0�E@��S�'��Cގ�B��ܕ���<r%y��sgm�KW��SZ��V� x�转�E�I��_%�i�L��|�iÒk�U}�8�=�S����@�|�F�+����r��y}�M��fYX�������`���sM�cS��_�WF���e.j�Gm����F������G�7��+8Ϯ�
��KUyD+�m�70�y�DKHb!)I``0m����;�!O���eX�'oܡ,2�S������x�{���S�ב(�'�{M��� �y^U�_���8��	M��O:��Bz�zC�ؖ2#���y��	!0������w�3:�gp�!�^0?���~���տ�Fџ����>"q�}i0�@�&��؁�{�1?��%0^V9ėt>�?�4�����,(Z�,�{+ց��� �$��aȓ�p= }X�Y #�R1�	��Ui�=ӖХp�9�[��l�r-Ijy]�&�k�e!�pJTV�����!�
 �]���1�&�����#�~�7|�xG��A�4']��(�z���N
�2ٛ�,ųU+�oE�X�݈��x��!����]��t�[�S�GU�s(��C�Z�\�W���23m)#IF��;������0����V�����!.!��\M�<r����PNשC�N׭�f�0<�R���~���9{��9}6��!��׶����"ku��9�E[��&\�i�Kϕ8p��F�m<~y�c %E*���,8=��Z����Z��gA��^FZ>{�q�LF-=k�25v=��C���MF�w��78mu|��~�M>�
����n�I_�_[��r��2!�mva5�`1��_X���43����(�-�)_��c�T3����.Z�u���r�V/��ء�2��d�#������?f[A,Г� %R����|!7-f%��q-L
 �&a�՟J�k	j(9Sͺ 1m{�C�P�9S�Mz�J��7��\�M4�X������S���!�EB��}���ʑp��j���(A3v&��=��~�	���S}��YVմ	�FUY��|��ڰʂ'a��{�F���ԍ5�U���qgQ8�bUKh�!:������[�H6blc<�b%��{$�y�*`�ǔ�8�+'ެ�A�%S�H�W���,�pR�m�wۧ�;����8�
(��ƚ��8�w@������yA �[R�yPvfQS����N}�86 ������8�5 mJz!��>���-�5=,��֠I��_n��=Q��H�H���ݝ{��l��ڥ���ȍk*#�1�{.o����G��\ '�`"g���z��p���=�BJ�&fOJ3�&��)��4�D�w^=f���0��A��vg��$���G�s޹�A�{$�	wK�9 �b��#�h|���qx	[<u������c�q�T٧��6C��� X~&�CW!�Z@�9o�++��}/Qt=�AP��J���&�f��T7 $;���I����>ݢ�,�S���UI\J��p0"��6�|W���%�����0	oM�R���l���G
<���H�k��l�q5��|z�n�3��uY�}�+yXX��+�Q�� 9�t^���8=���ݑ�N[o�-7�����������#����n����"�OR�����Zd}���s��_g�3�7d��1�~O����Kh0���hBSiɋ�
�8^�M;����B�׬�Cg�SR���%Y�{��gf@��E�-��.��s������RO����V{�8�P���Ϳs��d�;Xs*A�A�E�k����AMz!&m'l��k�9T8������ ���@`�>��#��&��m��R{����	��˳ ;p��>�sl��VQ�g�5o�����1��1�w�Ö)��P�������%,���?QA;�#����4ޜ�ǈ|nf���Y���I{�N�䶤����{�T�gq���.mD�6ɇ/�d;HQ�E�+䓯��(n��~d����V�w�d�Ҷ/aQ ���G7�3�r �؈��D9,:��?}���)M�^��'�
7|e͜�{�Sg;�L�b?����@ܲ�^i���
�j�+�AN�J���\H�\S�y����ɛ��a`II}�+t�qkg��0&���Xf�+��k�㼿� E@����$�T���w�\�U9^�����ڵ�7���w�4��J�`� �4��|j�D�ɕ�hۄcn�F¨���~D�z��9�{�K�&���K��RKW��$��Gi��~��z�^��1��������3�b@�@ò�8~	���Ȱ��ղ>F	�ONkB�qa��" �������5w�c�k8d�ǳŻR���n�t�@#��8�0{�-&*�D�d��k��A�QE�a~�J|�IP�a��,b��H��K���Ш�D߉��f�ka��u�Ƞ"�"�U"��dT���`�O*R�Г>x$R����V��gu3;�u�e#���;��|��ߤW-���:��U-1�y��Y"(���uZ܉�v�4R^kP�AOBm��s� 5�.����{�J�v�aOn8��"�=��ͧ*TjO"-ԝNY�B�X[=�������O�f&�axL Bq&�u0�q&@��{��}O\�yEt6����i��}W]Ӄ��B,WH8��~!��[*�
ࡎ%@�"&�a�Aw��T�ce{���ӂ�6l��Ǭ[��n`�{�Na_��ҹ?W��z����{���.{�M�x��Oņ�NN$/��DJ����&�X�`���[E��T�~����֬�#��'YJ6ֿ֔�9�����3��Uג��v�kU���k.�?��I2��6K��_^�cj����V���b�Z�;���O;��i��-�Qb���%\/2+NeG���u$�1�GK:U�����5��� \� ����tmಖm������)��a�mz�R���5 
��/jQ��uo4m1~F����D���])/�S5�Z{Y+���){˱փ��z��$����~��ڢW7#�}���5	����p�Ռn]f?����{Z��h=�%wq	z�^��/���3�A.��Fh���"ii"���[�>�9
�8��̟���&�-�y����>,r�Z姍h؂��z'H3y��cݘ=͸ �9����`�2��Ȫ5�e3}�4l�gڥ��4��g�/���͙�|ϠU��{71����0y��.s����*����OA�u?�����)�!���I
��#O��	�L�c/^�d$XɃ&���y��ס�?�|�|<�D�\��,��ٶ� ��)٩�GB����\=��e�1�&X��;��}�'���PM���奖 ��4 �.!�T�Zr�+�}�'���6�_t=���Ok�.�JLFLc��\{60#:J��w-X���b�lt6�q�(�h���J'�O�!�*�1k���*���!�� #Q�(ڛ��^�}�_��37`�Up�4p��uD)�C����C�"�Я��25|N+$���B�bZ����J�̙"����J�WY̓��Y���?;%�T,�R���1u����ʐ[Obis��:�7�=5�B�8y��"��yt��#n\g~�ت���5H�N#�kk� �5���/�9��ת`������Ri���N���/�S��q�3i#��R_5�7��?л���#b3޴�V�Ӯ���c��G:bsę�yV��&�ۉ�����؈Y�f���wC^����^ �]�˶qn%����)�.� �p�,���j�ɯ���h�bL�ˍ`�/]�v���Ӏ�p�/�{(�_ŧ�{{<��~�gQ)l���P�A���ی��B!�9x'��L����6V�TҺ�No_��I��q�>^J�o.y-�Oi��WP�L��Cr'N�%�D7q#����:!���Y��|�2Z�;�	㪱Sф��4bJ��~^�Xa�ȍ������o<hS�$�(���3�J�<$��Gl�0{P�/�w4�'�wz�Fx�9~�����o@�:R/,��.�-Κv��z2���Τݹ�!�Mä	�h�atBX]�L��bCM%B{�'w�Y(��eL+f��c��)@P����s{���r'ꕱ�G#�θK:,�H����ܪ>>�U�Lӌ��T��C��[�������	�hJ��
���i�<�#���a�����g�=il����h1"{u&��� ��9z?�v�Яk����8��%�*�Y���1r��(�AC�ۯ��٠�^��?L�ܛ[U[�+P�?;yc�W��aL�`
����]k,����r�Χ���;�Qi�g��c~m��|�1�O�T��.�]L����#�[vw��.��Yr�Sņ�N!:L,bq�/����iT��U"k��x O=-k��F�k�qK��z]���y����0�ɳ��:�v�@�K*~�$#���kgS����\��N}Ԃ��K�Q�g�l(!:���+o����M�;�����S�Ǹ[aci����!�܊i`�'��,��d/K��T�/X���
Ylј�n\c )��-�,��`5Iz�{= �ƥH���^�Ӓ�=�1<��\���s�n i���3]:>��{|�c���wv�^؏���]$�ިYq�M���u3N<���?do����N��?�A �.����S3��"�R�d�>]qA�p�f9
�i����h�R�`��*�hK��x�O6�������J!�[���§(���t�� >{�$P�C�y����\�?�Æ����;e�����Z��Ҕ�r���Xq�����P���$�@fU��LT�FW!v(�(�����?��W��'��vd�܏���޾���u)�&����1���b.�	�J]&�0�
ϝXy�����VEozS.!�:�oAp��nǬ�=ѷ5������\�3�^��°�s�TsY��&�6�	b:8WW�> �<�u(��Ψq]�j�7����ҳ$��k������b�w_��Ѐ�ZX��Q���+0KA�"қĩ>�[��\����ΐ�9��NK�8ND��e��O��.��望�]�z�������T�t/N����y��c�����Ct:�st��W�I�=�0�����.�1�Ǹ����iu܅��xW��d%�ޚ�u~u϶"���|��K�TDX+�[ Q-f�E���RTeq���ܛ���jT��a5�ƭN�B�A��V��de��6���b,���'�����`�*6ȅA�BM�uG,�z�w�(ri���8XCǢH��_�]&K������o�[�L���EԊ�ڒ��3��:���#N'0|^��@�#�ÇM�m���"T{���A��h�Yq�z_�&�F�Ζ�GX�6Q��L�d���Hh�������ߊ��E����3\����=��n�G)�M�@�����]+P��K���u��e���-l��C�K���RH�I�s���	|�W�y�mUj��u�������)b��rǍ7w\��DP��S������o�����7@j��ߞa��
yo��N|���j�����G�pe_�#�U��9Qh�(��e�y@$�mq�#�+�\��SӲLe�@��k>��$��I
��!;R�4�^�Q~���x�g�J ��V��M!��0"����I�Y�
M�~7���5!z#��e����)`�㵾�֒��t)��.i�J"z'�4��:�̰b�؜��{�/�t~���ҵڼ)�[�'��u{�W�qS�5��ǖ\���'.��B��WP�BLqL�3Y��"Ә>k&��r�]�E�Q�j�^)n+-q�^MJ?�ZE�����=��5D�)&����������%rC�?8��L�I#��v�J����� ����C܆��'�t\������-JryO ������z�֯�upI< �>����������t��% 0_JL��H*��5)�����a�0���(gd����;I]�3��HL�wp��#)?7.��_&>��7�i�]�D'��g.*�b�a����������<���h@��.�:D$E�?Q�o�`(8��]@I�D�����3���t�ߣg ������<��hI�1�(�ߐA��jTc�ޕ*H�b"�������ʞ�,�' ���Q��i<���4��笶\���X�D�NfZk��~ŧ��������e��E�?X�&�l5'��3oα�w����Ff#��$�"�������q6BH%d�+2צyv�86 t��{S���!����o�����ݸ��'�h>���se Qxf�dp4����pR�� Aoq�t�ђ�m } �!�r��Y�uH��o��FF6Ӷ+�`,kL��βOAb�d%�]�N�n7_�&��4�5_���m�T�+�������G2��RR�t�����n4�'��5[r�~�����c�.�[q�v~p�KU&�e�)�)�H�pNSo���l��~�?�ۥ6�<�<S@|�U�h���;���u}�NO�r��JB|1��쯏!� n�E�^/��^}��oH��hۇ�Q|0x3�<ᢑU]��`$�L��p�i��I��&1m�BA�#�q���(��_�MiLԤP{�Ԩ� ?!��)�{������cm�#�r!o��g�O\N���XzX�x':/A��'1��\��~"Y9�V�)���=g�{�L���z)�x�THP������8_�B27)5>t�Pd��؜�y�3�+d����_lڑ���_���Fc$�<F�"��p���~G��(���w��OvI��pm�*��~�=�E��W��؂(�#A$ZM>�f^z�P^�6XBTF�[2@hqyW�-���E̎�Y�7�횂Z��TׅGٞ��?�\����5�J��/�~O�T_f��0�c:��[+��4��y�LW�g2�0#�y?�;3ӝ�5���0�9�_#����Q
�Q~�%�5� �гQAY�&~��B.�D���5=�����!;Zw�I�g�s�#2g����m�~t�,K$�~22�y��9�1� 9=�3i��y �1}o����Ո�V��ꈳ������z/��wj���@ʗ�U\����$Ǘ��)��_��4���c3��kך���`2��,N�eӻ�F_�ao��� ӫ�L�ʋQ�9��g�A_���@���O$���ux�-�?�d�� i�q^@�aU{/�c?҈�ӟ�(�Lrn�Υ���R�ᨖ�wEi�����"">�+/����:Pؠ���MG���·�12>�.���1,C�'O � 
�T�2��Q����ZO�j�eLJ��ES�읋��F~S����0mPiT��R��u���������0%/���,Գ���Z�̜���d��]�B���՞�I��#v<_�3�X�]`Xw�
��XB�՟հ�*��kW܌!V��������.I�a��v��߻�R,b��PGr���σ�R-MSè"�`/�W[�#Ai�X��+������T�"�KБ��=hG3\O�5:�oU�'�|���c��`�b�&�$���/G��K��?h/U��B�~
��� S��
9���S'�a�5]� ��.����b=]���h����Zo�گk']ؽܹ6�eR���Qª  R�uc�Ŵ��ʛĴ���rơ�è	�]יh�d%9I:u���� �xyX��hG$6�D_6����98E���<{|��ű0����&�t������9,_˸������V
F�o�x�q�����N���z;�"�d[�9(`Q���@%��\��Ki���/Q�U|ҍ�)y��ƽ�c��/p�m��aJ@IY���y`[��91���n��/^ ��p�{J�' z� OKv�5uq���#�hX��h�0��ݰ�3��}Z�Y��������s�E X���=�'�_R�uc���f��F�5MЬ*���`�09�D�gX�U!˴V-u2`ZJO���xU��Z�?0��]*��x��U�W<c�o�ΧS�/����/7�^� �� �a�0�E�D��_H<���g�(�Ha�!d
���!蛁���^���P����6<�qk�6|�G~�y=�e���=��i�r�;��P�Є����Z���T0���d��H������l+҃l�me{�������W/�Z��hR�Ĉ��F��Myp�Ad���x�&9t��]���iA=[���3�͗�_�$�ceL"���|L�Y��<r%���7�)��(��{�"��/K��&�}�
:�W���N�oMVg	$P�+[(�03%ZT��;� yl3G]3u�}�+K�9^&���m����g�����x��soۃ�;�g��E*@2b_c x����dY��#ˠ��Q����ц�Z����0:�i��Q�/�i�s�$H���f��@��
�L�G�ʵ`����q<Ǥ��o�hJ�mH8�t�e\^���u��#W�>�5�\:ɞ�l�
(ܵ�\LN'�V}ѱV�OrNύ�/��kO]��ŵ�f0��	��-�� %k�d���e�{1�f��Qk�-�$���o����5@I{t�o�b�;�B῏�X&Q����WC���+ʑLe\O������H̖�T�l�)�$H���t��5�:��V��T\����k�0�E�z�E��K���_q�����SH����%W���[�ߜ)�"Ӯ��r��4�E��$s+FnBF_�@��DU�����5�R�_)VXt9���n��W�Z$��4��ZG�?�]����;�7��p �	�:��yе:{`����{����w���~2���Fxq�N�!�B5��Ԝ�TvEkIƟs%S"�6F�|M|��f�4��'�K �r�X�C*�S#ljr,���z����n�(�Ji�8��@��U.mii노'V���e����� ��vL��գ�@{`�Z������.���v�S����Ԁb��=������)�Ӛ<��P�6Bn�ѣ���S�1l����f����1�i�~.��qx�g����٤����}��^l�y����2��B�%��N�fFB7e���is]���)�m"�b>���G\21�K�.~�?�1����1���GFA������ZV(1��P�Tj#�굉�Pҏp�Lb\�|r���v"�3R�9�w�2s<E���P2kS��q��nܐ�>�tʿd P�t�cI�(��)����0r"�}b!�ac��5fo��Ôl��#L�%f�C;�B�?�O<�8�!�r_y�Yօ�ףg@ ����������{F`������ey,	M圉���H��&|��u�G+K�kĞ�(*X�j�1i�(sײcb�O��P[��");���`5"@Ѿ�7�~�!�;m��Cp'[��Q.�Z,�(���\58@L<��`O�H��űT�/@�6+����zJ������C%��m������Bebb�g͖��%���\u~��J�ǝ҇��gƫ�?��~=�C(�į��8�G�P�ܫ���3����O*H���N���5`paRY���Ҳk���g���p��k�U�ߗEcݥ��;S*v�Eֵ��qH|4����d&e��l5q����H��*�m>o10�0O1�X�Y��J����Z"�Ȗ���P��En�+ &��o�:���6,������3�]2c}�w�4�߳�a�R��}͞;M��8�xh�4���tC����bX�Y�_9v0;#u����)��k�߼�ٻh�6�% Kr_߁��dY�z��:������J��{>~,$��l;=���:�d�&��������]��j~�ё}�Mw�Ȱ!y�XB��r�T�7ZXW �,��󨶝ȧV����:$��֧�;@{zC�p��M��f� �q�o ھ�\6Y�o\�P��L�ܱ�5:��]��,8.ջa�؛(�����|���,����/#��j+A�}�t��V���!3�<�����D�5dTA��[o5*m�ӫ}�� !��sB���M�"�@���ם�_Y3Y�� Ҩ�"��$��2ٛK<��	IS$�j�Q��,�8��:�k�ٽ:۰�Yv�|?z2d=�	�_޻�c����@=��5��jO��r�G|��=4�O�߷��^_���e���O��|+��p'?s�/�:3�̲��z��=x ���:�}g���=��UVq9v��mG[��ұ8��`M^�ws�]�}�"�D
*A����O���U�k��-�*Ɯ5�8����ll��-�>�_<��+�0�c�4l��}]Z�9��T��m�)��2�`�ԡ 9�Mm?zIʂZy\��2�M��������+:��ܴ���am���B��t&��]�s�>����i*,�i��ŕU��3=���������hvr�D4(��!#,T��YXQ04C�Q�>�|���Y�!RDɖ7E����Q6)V���Z�u#�aآ�v��9�ciwgM%��3�楃��]uճ�J���<��]��iI�bk��~i�G�D�����	�ZA�7�hpml��rY���7+4��Eʽ�S�~Ƚ�Ӧ��t8��/>�l�%�HD������gߡ:b5#��@��ɰ
Ys75,�ґb�^���,�~����]6�үN�V�I�&ѐ�?�9z�������}S��fm����
{=�2Ydg	R`���$�|�5o�:�PCE硱�W�J���`���H�=�Ο�I��#]�T�6^�XŦ>
�8��>��W�"�>#���8i�T��\�߉T���2�  9���W�/׽IxV|F7��7��r�{ֵ}!���N��ž��kB��;9��4S���[ob��o_�D��Ec�SG�2��;>_Z���x�o�w.�����?_�g����Uj�f���R�,���.2n=�
�t��=�Q����-�a�p�:��H��:#��O�F9�a��gj's5VJK�7��4'�J����� =䡯#
.�ȗ�.5���z{=Ն7�5��[��%�:�;#?=�1�np�q�q��Q��!���Gb~��q*F�&���W)�"�#�aW^������&'E��� ���q�Z.fʚ#����wbg��~ӳ��fԈߜD�ġ|&�Z��xye)b�F:h:�r/K/)J�է_��줎��5=aЍ�O���a�0���t����tm(�ڭ�~�s8Mo��wA���:=�քQܵ�����D��ya�+s|*y\="gs���/-�Tе�h)�O��-��r�"{��O	�T@z��lR���Y¦�|,_m��}���|��qC�ы��K#��nW�r��A^gגԯ�PW�]��>A=!�~d�@�5q1���(���3HZG�R��3DD�N;���A��|"���g�����%�b���W��,l���1���5�Sz@"f�_�k�}ą������b׊���WX�@�B���{�Km����� �8!��]i�[��g<��=��Zs�+u��	?�g��XK���dt�:���z����b�N.f�t��ы���d%��Xi�l��W�J|M;��m.���S�Ķ�c
���w 3hd]q�8�(TB1ё��K/^ư�����
����K93>5�A��z٩�ՅN��˞MZ���~.���7�
���*H;��'{��вC����Y+�
��B�9�0~oٵf'y�u�q�O�A7��Ơ��[�W�x��3�0�hu�O~���Ý������.��Ϯ'�C�z��)�Kա�O�zU�9��ك�i�W�g�ia-��K�g{�G��_[�=��"�����������N=Ë��������0�,_��m�����8£��'�6�M��!lt��p�?d\� �2�t�B�K��G�[����-��ut�du�\�ʖ+@�V����}���� o��!Sr�L��vQ�ʳ������ܦ{����$UK! �l~ϛͧ~i�kqٟ��~Q���2Y���j<
�QU,G�^�b
?]�2Y����C߭�3vKl��N����RB�m�m+�v��"O�~�_g۰[l�_�*��$��eݤ��v��y:�]iT��h���O�a�xH���udw@blؒµ��<*ߩ�)�扮�gST֐�D��-�S��m$,��4�	�$�2��.��,�uw'��oRj�Q+I� Kw����M����� j��-We��۱jAb�:���� �:��
�%:���b����u��f�R�k'NU�J>^��Mǁ�j�#�$�����Z^X(�?���)�Yʁ��~O�gz�E��Y͸�
O`���|ㄬ�4��r��V~Զtն�@"bhR	蕀�9�> �m���w#��Z#���I�[��d�p/1��%��#��<6�w�I��m�|�U�/R2:����3gM���/T�=��:�F�g�����6O쮏�.1��8|�+�W�@��k���u�]��ұ�F��!����ǘ9�˚�gǴ8���\�w��5��2�U����ne1���H�"��2gD���I=�Qۼ�/�|KP�Xm�Zo�d�:�5%�@=�Ű��i~Ἃ����(6��Z�e���o�ߋ#S³�1E�oӵ��e�w����(�k�y@`��T��#���W�{�৵�8''���X��2����6��D6��w�΂o�7�t�n��nfF�=�RՅ�Xo��p�j;���Q�ٍ�p{��P�M�p���҅{��
Z<L��
R�@��?��e�j���@� ���{5��~�a�7�r�*�j,���ܺ����_�x���A2X���C�ǌglN���1y�e�g�R�6{#�����ҵHBvk��5�ٜ`1w�����h�T:]����:,�_���)NeD�6���[�͛�]��=m�M#U�P�!e�r+K�\ߊ5��	#t��d��W��C͈�n��vqE�g�.Ά���
P�Sq�
�u�%���D吟�2�_U�����;j�!m��pm����z�^au^V�x�UW�P@h�d�L,gy\�c�p_���Xݚ�	����"v�A��e}O�IR���V��x���'aitK�p;;�YX�Q=AW2��h����Ҡ�(�|�[=���gy,�B0��G 
g\���*�B9�;J��F�� U9�i���3U��"�.bx\�FT�b6ZA�{*�:�^�b�D���d"d��>�NmEF��H�ޚ9ApՆ^<�]f���	qe`��պ$+V�Iyë��:��#�AgbpC��,�E�k���)�C�,[�]-aJ$K�B�//	�oӾi�:��a���c�#?xj��B�𧌰�����2�5�Z=&��Q�=Xd����T�,�H����獹�ɗ7V/P�!Q�t�[*�	 ��*�U�1붐�w�ѧ�o��,�~
���柌����+ڮF�G�w�W����M_�+� ~���v�gR��9嗈֮��7wT�g��t�S��2���{~ҔS��ז�<o"=^V�q,��\�+���z*�Ϭ�Wn@�����6h���X�7ǐyC��l��z���&*�^�-Le.�J�kH��K��y|�Ũ2kd�������c>7��hd�8�OqXgX%m�|T���������Fx�+�5ؼ�+fl
�v]ԑ��uH��D��i$Q`���Q��E�#oo�7�q��EbJ%c����0$��� ?}�Z')% ɜ�U�NL����o�[�od�VB��3�q�����D-��Z��ɖG� �$Y�ٸ�}���fI|���"E�P`�,��ck�[��Ⱥ���!ߣM��_��@�����@3Ec��n��t��4V+�ҿ�W̛�R���S���&����J}tF��YYd�-�V��!؝^�j�&u����r��؂6��0�}<��I��,	ҥ*��n<�ɿ�:�u����c����% ��:Я�5����"���������^��<	w�E��ນK�˴���:��u~ Z-j����PC�ٛ)�W�P��ӟ�S�L�B�f��~
��f5��xe�֣b�FE/��1O�.�rB���nƷ;fɹ��{���34��	݅�
����R��}���J�H�;"2k4v�XyE��� �M\�5�BTG��(K1�F��F )�W�Ww<�8��|��?\VǶ�o���
�ɝș�=ʪf����4u�� 5�ԃ?}�V��ה�p��(r��,�0�������I{�m��&Z<eE�D���p��t���b����d�����"E����>m���X��K\�!�k����ًD�}��o`2@]V����JM��=�F�?������\��*�q0%��R�!�)ʃ	ő�Gͬ���`N�6Qo�۶�N,:��Ӡ�Sx&/5"CDp��ZV��҂�G8Q�=<^;�E-J��5�	�4FD��x��l��X�zn��1;�CE�0D0�1�d�I�����зr��@�j�6�M����.
�r����S��0�ly�88�����/��kEm�Z�&�`<0���s����M~�q����ŧ@�����a�e?�4BM�Ⱥ�Aİ!\�}l���M�BW��	�{N2��yO:��˱?a*�|���f�3�a'��<�t���ū��������`�b��wA��+#R!��c���2�)�4$����y��oʦMሑñ�Ŷr�����,n�ԏَ����(>v�+N��gA}�ILDj�6������>j6�`���H�����}f������f��2��~ЭY�pq�]W
�۝�O�a�YL;{�j����63�������Y�CQJ�����Q�Ţh40�Kz��Ԟ�kq�Z�#�LҌ��j3��Մ���,Nt�F��Z6��kҳP��S�<6�{cҡ���Ľ�3R�MB�*��Hb���~%w1�=I&�����٣��أ�Lh�\S�8�
���=	�k�;�}]���?�������E,��[�*���<K�������L�=��U�P�S���܊S��^&�c�Գ��QO��]@��Q8t+$�پU�7%r e��	���{��/�����"uN�K�;�&�3V『�M��d7���5�U5�a��9#�^�7`y��Lv8�H3θz��i��[+�Ob����MK^����ϐ��U�SW[�ǵ�[��_�l%F)1g�K��$<�����o��wkT����x�-K��r n0X�kO��XZzJ>)^���������AmC2eA���V�<�bު{����Q��KbhO#�\7�QO�4�j�����o��d`����'� ��+S1�w��&�&�S�SJ9���mgZ4]�\s&K��W�xJU����ӫ�:(��9�u�s��Lf9��{���*C�ʖ�đ�+&���PC��"��T�4P��5O=��L3��UL?�`K���g��l�@ZV�}~=l�8����#ld+>�ĂmZl�`�0�U�~��ׇr(�$av7�puC�����YVw���T3S4#��ĊI��~R�V?�AǦ�XamX����۞���Fnͭ��:�4qw|�Սt�R��ן�m'�n�z�DSLp�9�[��娠!�D�8`0p	�Elb� ����q7k��[�T~bȃ���;`R<�gb��I˄���Fm��tG^�t���\`���Y�4�{�.��s>�ˊ�O�e�E|���x��[�<A�R���q�!2��GΖ� ��=]L5$x����7��$yf	�������'��l�8��50b�z�ĉ�a�����f�j^Sb��e�=�{i^7� �ptS�>��'����P���fև���E��N�Y�K��E�ޮ v�tHs���͋�}"on_'����@�z^ѓ0��{p����}����h~2���؂Ɠ��;H����r.�g)l�%u8_�22
8":3�oR�ۋ�qi��v�M��to`@7�̞�&0���鮳h���$h�[+�l����#<�����^�B��Q�)�/��}�
1+uR��<��S«��_�,	G�,���35+���_��x��;��� �A2�`B��$�|g��&��w���tφ��&��׬t�����	l�pI�\D�/O�+�V�D��Ӎ�R��\��B�Q>��/���nZ�{��Zu;DJ	�r��2�\��� j�^ogG ��*.� A<�삥ͱ�V����ʣ���\���.���Y��Î�ӴO��A�F�?Rj�C��!2�����|b�s#Q��_'1�5ذ9Q k��6��!e[��[헡�o�'���/m��������X_75����T��賦�2浞�+O��S�l��
`��{�G8l�x����8�ټü3[���b
��M����
ަ�z��\.���}yQ(�k#�i�%��_ �fa�X��3�gh38%ڟg!_J6�kߊ��0���\��La��w�u��>���5v�Uv����`I����+6j��)l3��7���ȝ�X+�X�k���n$V)a�=���i7���
�`�,Y���˅�lzg��K�#�H)��*�i�ƒ.ёrv�FS��ӿ�#��;:>B�R��f[ϔ�s8]]:��8j(�m�(��Oe�I6�[
��a��{����_*hd�J��~R��C"ɼ��ac��%�xK�uJgw�jLޅ'��
��,��7q��O��"�p�ҵ��O��v/��RT��0�y!�vP�1��@�Q/TF�m�9���u������qX�Q/�JdT?Go�ρ*<�`;\�pUu�����.�,�IO���p��Sj*����iL��e�>-�j5kL�50Tkk1�Ħ^��6����V�gFs!�-�Ӓ��{�1T�Q��^��k�C�4�}���~��\�LHO��$�i>k,��#�E��n��`h�>�*��)h\���n��<�'Y�hC��%5!�B�1�j!��������"���|̇�?���վ�vR�U�X.f�Ʈ#_��"�a���w["{��E!5O����AZv�+��sA�4�lCH4D�q��`|%�]�jx\Y�(V*Ðݳ/<�~���0�����Y�_Z��j�HP�ܓ{���{H#�e�+,.s�+�������6MA�UL��pmq�Ynۓu&0�&T��.O%���ă��ڒv��=ˌ0�)�R�+���U�O�����-^�r�9�22Z�c�D`;'t��]'v��16��h1�-W@w%^b:�E8��Ǯ�]9}�Ң&�1x$��D�G��Ŀ��U��bHb�foS��/rf�dB��ｄ-���#���eg�aj����W|r�X.պ�/y�h^(C �K3\���u	FX&�� )�4�l5.�G&g	������np���^�����;j��Z��n8�wOӞ�//�ٸX��h�oF����'%�#�Ty3A:UX�����)��Hfl�;ɀlP��_²i��C����dW:yz�����Y	����dN�� ������񨰎���s����=���]�����}���e��r3��EL_�}"����V�"<��K�*�6`P6Ȃd��?�=�x6��e��[n?�\�aP��J�q�[�Q ���G"��y�%Gx(�N.�.:GK~��_p���������U�[� U��SΏ���s�����F�����ȈrbGj�e�7�X�(	3��Ou>!W����RC����kZ��Jf���T�8��)D���Z�h��K;Q��.�x�EV���f�I�O�8�z�#-��<O}"�Y�����B]����P��O�+n}�� A-��P���2���༼�`>{��Ųl�S's�����`�-[i�����,6&������$�+��Z������2�c��8�	x�[���b�es�6�@>�0����|1���VZ^Ս��f��X&��|��mO5V���\��O��އd�	�X�h�lӳa�w���R�ʉ����d]�_j�K>&��4�o���M����0��6��X:q�h�
��t��@�]_)��FԪm��T��L�P�oy���Nd!���@�(�͞X����x�͙�B��ў��K^�1hϜ����֟<[�6��󑱗'*1����G�08[���*���fV�@�cY�f<���mt�tfP�X�l{W���D�ҍ�
b�{u�+d)����6�t�3#�+pI��z�F�lD����qB���[�xXi�{Ude�q�DqG6eh��',L��!I �n�$�Q�
l$&F�*u&�h@��?X`��6��(�> �߆���������!d����#U����&x���Rz+���6�t�TkG�I���2�*M�L�����sB�����]pD)G�9ZNp��-2��,��,+R@R
�t;�>	n�	ֶ�E�n���L� Ob��:�|�m�u�&�t�OFQᑯ��A�\���K��!ڀ�c�YCA�Z�L���G-%�/����T�th�j������V٨LIq����-X7ަ"�~14�MU'�|P�Hš��+���Q�_Tm�땜aD}�,�� �N�g�9�r���<(�a[M��D� �Z��<���B��'�[Eg�bK��]�w��؎CJ3T-�/bZ� E���Ê<�l�-!�:���s�c���[�<3�k;��Q
�*�҃v �乲� G��멏���0��C���@�b>ޕ�h-ڃ�HD����ʡ�����Z��̞ z��Ce��<���@t�G_�z(�(�m��c�>j'��Q�e��O�G��r��4��*W���e���kΡw��D���9�#���Sj윣:�~; �,�Cr��l������^EI��=����plvt�-el�C]������tc/ٺ�2���g�QM kp�~�ŘKk,e�}��ߡ=��jb jc����C�1%^Fzǁa�Gؐ���`|D�|�6�b�XĦEcV4�&�6Y��CRk�����4 �5
G���J7�\Q%Ԁ��#`w�W����8N� �(��U��.4+�x���
7rq�l<ɝ�[�t]Ъ��_$�z��R8/�T�?<�����g��s7�>���.ٯ�Gخ�Z5�ΐ�nƼ&-C� d�/x�ԇێP��"��[�2L3�G��UIj!��:rG����~� ����\�/*��#@��꫶S��^�O ����� ��0��A�T��9�~�yA�Sc��������Gt@���h!��YH���T��� ��tn����7�d��~V���WXZ��B4�m(u_�V���������wW��YUmtv
��U�q�_�035ˣC��s/�<�BqB�C*�1�g��V�J��)�q))��4{]}���r4�F��LWX�ֳf����:���&9}�*(�6�Ua�@&���Ֆ���
�w�a`���q?s���?�b�s�/�Hݖ0�=T�2����Q�r�t�K'�9��`������Ǩ/[����&��O���W~�ڪ��o��۸�h���z�?Hߒ9��v������v�wC����%���l����6ʗ:{�A�v��OH)+�Ց�tqޞ ��P]ti
�}�)�Њ���a<e��v=z�\�A�����5�o�!�z�O��ž#(�"��c��PP�B�<��/-��7��-"�TӘ�,��8T�%Y��Ӧ�H0�j�(�K�T�  ��*�*��mc�tZ�/QT1S�K��������
\�{&�ik�n�;��E��{i��ݔL�	K��k�з���6���L�,jw2�)��@��X��B;��Y���'�v=!��Q�����9�#��ս���GA|X2�E�>̅?����sk5����`J�|b�$�����~enK�x��U�j�:������#������Mq�t~=�����}gA%�O
��ѝk�dj6C��䥤B��_��n1�Ӎ"S�G�͐I>C�ʗ�
��_x�?��|�a3퇈E���R�O�3y�vϴ�u���L�ʪm�X��<�S��݈�	��wX��²�_����m���Q�D"6ꨝ�E�
j�]�̴?Vq+����|K��<*e�3f�g�7]u��ؠ�Қ��U��A�����5[Li��_�}Q^���%�ºlO�Wa����f~L$�tO�[e�@s�V��Lx�cac���s��t�Z�����F:g�K}��uq����%-�N|�@Oyy�4wS��9��k#v�r�&5_������ߏB� œ�������;���#�`E���@	! ��\��U���qˢd�i���Z���I� 0����p�C������ɢ)Gl�h��B��_���h�Vp��l�l����6�d�ǫ^\aEY��q���4�$;̝�m�K�e�Z$&��hub����T	�	P! ~A`|0bJ$f>Z�M��o�e�����9|�jMߗ��. y�����i,��&���U��\�6��y+jd�u�QA���n\�$��#<��,�L��:��[W�63��B��ZP��?+k)M_hk4�89�'�󧌯�C�`�l#���C���W����M���e��KP�0�ޥ/>xJ�RF�H���,��,~�'��ʍ��,[��-�|�J҆<WF@ֺ���1t:��� $�u�@m,���/���gc���Ib�%آ����L�:����`���p��޶�r��^��D�]��_�·���2_�v8w�@�|�:	��、f|"�"���`L�k6x�� ���l���\�)���(̪�$"uDO~��r�0��:6��G���n�$�|a�郑�/O�:��C���*�U"�y׵tk�+���tL=����M%�$7���5�A,��u��&R:.��;��w��R�q�o���<Gi"�z� ����KX���E286��?d�٧r���L�U��L�@�rM�VE5�_}���4��1��U-#�?��l8� GW���`��p�N�� ��}����'ɳ��wHq��p���@���ܪB�^�L��T<�d?*$'�~�B��S�ꬺM"L}^����86
�|�2 ��`�Wf�p�k��C��S���?�4QB8���C�q'5��L�����v�|�v!p3���`Tn�<�w�h1L���}���^�U����'9%*/�?�P��r[����R
R��T�B	U4J�UU|J�>"�<��4� �5�7��>=����~���.R�x�ȹқ�\~
|��	4S~>o�T ����^q��� D�������)z�{�`0ؔ�?F��9W�ny�?�O��WS���07��?AG���â+���lۈ+��̘��@��ɵ$�c�>ߐN8d�� !�Ϙ=	U2��nY;K{�a
���Q��A�_������)���tA��G����Z����Eoxq��48J^��j��E���=���fɌm��L�k�WI0\�niəid�s���SA-	�44����?���ɀ��y�78�����ސz��X�v���>�^���?C#�+9j� ]j�w@�ɮg����}v󰦈��F�{���G*�k��p������l�k`;w<�i�5�tv{x���3�ㄈ*�������;P� wr�ZY4�U�ON�f�W�dV(EÄ�!�5�ѕI1����f�m�J�8mδ�� oaL,9�C�d���ndOƐ�3M'>ܷ���
�w��˟F(7?���G�Pv�ˏX�Yq9I@����#�:�sf��цg�$-nJ��t>o�z�R���ұ������2�V7�99a��k�2/�� 1x���A��P�/-�N��Ż[�pp�]b{I��W����:�8��.c��x��ݏ�cRq���L��"�A���˪�����K�s���%a�gO���+���Z�J2(�����9��(�$��F�댽�l�U.�X8:q&!l+f�����@J��Rԡ����]/a�V2����	e�ހ]�k�N6X��88�~��)�ܺ�7�qU������ג�O4�Nm��#���C����r`iSĭ's�oHH?��c�F�
h�������s���e�p΀T�lԍjΔ�o��^
�S�� ����G�<���I��
�V���\|��kA����vw�����v�a�cj������ײB𱶚�����K�κ�.��:�5���_5�R��+��k�n����+�vy�ݔ�I՛s��uen�g��e��Ż
e)����ش�	-᳉U#	h���{iqJ�*i\��@e���i�D֦��v5��� ;^S�n�d��h�'�˷���*OQ��өi�r�E�@z��dy]�)��!��q]�Ц�M@G�.��峒��{�;��qPYu��ݻ>���	(Gc(b�[9�k����Ы��3�jR�Jo�O`=�Qe�N�'!�E�6]��l�L.�jN�yn����F��Í����	��N�;������˺?��;�N�C4�����X��˻,�k���Ӫu�"&�Y��Lt�bO��x�6��ZB��lA1��W�Ā����/?�i���/�II��x%>k��=/Y#�d��U����U��*�v�ezV�����or�i	�F����'�O��-��ԧ��SM>Q�@< N%|Kl�zT,:a��'H�w(|T%zhW�o��*@&���Y�<!���|��t\-�8{�;�i^�2�E K�� ��&���)U;Xf�7��$�	J��Д��k;$��ə� Q�&rлo|;V(��@5�x�1���v�SE�2U��?��O�n�h����zbAғ9���TGy��Fp�:3�g���~�Lʢ~-�珦�j���5�!��ЩP������V+φo�������GQ[�����?͕�^���������p��Ց�ቹm�g���Ț.�"���??]k�7��+<� ���Ť�&�����:��lV�T��A1����dz�&���t�*��<�*9%�S"���i�2/a��l,�"	��,i��_q�9�ӈ��l��׆�ˈJ1��VA�H;��&*�U�b�a��C�,-,��B��������eJ%�!�A���=�68� 7`����ұa#�=��}��;���� �B�M�Q�����gr�� -BFܙk<���I��^����U��3��Eܱ�m_�/�7}��zZ��'/�3�l��T��*Ͷ��}��"%�SS����(E����F�ؠ����ϜV >E�7`�|��r���"�7�@< ^�7���k��Lz4鮽�CT|�t���[Uӯ�]S�r�ă�#ˇ2mS�Pq�$i����h�ɷ���>���
�C������{{t�`S���t>�%d��d�m��|:�̭�v/� �&�UC"�啠�5�,4�|1|!����`,�k$W�N�[.~�! ����W�B�b����Ovh������.��wU��j�{:M쮺�:��ŕ�c0����(U�ժC�9�d��qd�(��Y���p�R�A{N8��=�β4�-�O���W1�d�k�sn��@�3�J����dd����3�ډ.��d�;� 	�}ϙ
7k̮c�8�CoJ�!�.����=��JT�y9�����,[��tg�K0�
��$`5��F � B)�ۣ��2*nn�1E0���ΪA��  ��? �E$������H>�x{܁tK��ZB������ʅ��H�kH:[�4�"Ʒw|�]�}��&�ś#�(3���4�p�ɦ�YG���|��;����Ј%� �|v��x|��m�7�A:w��$���<P9��^]�KV5m���El�m������H���.�jKA�N�1z�fpla.��)g动OrT>;K/�(����,vg�+D�%��
�{�ui��X�m2FT���Q-+�³2�k��궿ٴ&V.ةA�Ay��r���Z�]��ar��+��d3d�ۆG�S�#��J $�Y�����o4�XOU}��l:ʉq��ժ�Xr�ۚhJ]�M��S
����Ve�Y�A�/�Pp4�S@��a1߉����I��q��9bK����7�U��	�:?Ʌ���b����I�~�<NW�S/�ΖxV	�[��� �~}���?<�~7�ց�.��7���uM��C�t�l<��/��KI�������-�B A�n{Es�|�b�4a��� �U�|��O{���.�Í*��sAύ��ٞ! ����DR����,τ[}#�S�����na�����9�}�|횲���p�?@
N�N���<-8�Z:^������\Ĵ$w(g�²�T0�����FLA��&AN�|�H�?֤��4�x���ݗ�Z��b	J�f�>����9D�MMM�p���ނ|��-��Sߛ�����.��Ƽ7��]��e��ִ�i��c�,�ꯒ�,���\�u��4�|��rM��C�X�	�Dɰ���\čM�����#w�!j�=�Td�3'�xe��L�I��c�Yj���gp�v���D_�¼�0�T�1���rp�o���Pr#LaE�<��Ӭ4��"*�h�c.}�q�􃡿���&��qEk����� ��km�ЈU`�jvR[���7�?/Əit������\�bE�RC��l�y|��(M_�z�� p��z����[/�q��vs8d�9aC���Ҷ���eV "mnt�C��õx��B�8���'w=��q(����2�	��-|���*��?�~��5�80Nx����bz��C�/s-7�Y��\��`eQ��G|�hV�1`��#�%G:��.V6"m�az�
q2�Z�}s�c|X�ڡ�W�����3�7��Y�E����`Je{+Ӧ�5/��n��9��nF�6O�t���'�49�����Ky���f���:�ٙa,̱9>=/��8c}'i��Ov~�!���;���pnGy�4��7�ߟ;2�2�<H'}s�F:j0����<����@R�(�u��ոsa�C��~�p�
��ydY��J����WpqE����tW�g��d�&S��w��XVRyov3/��)�˸Og��ZT�iK:���|�+~�![����_2D����
�BKsQ�7(��Q/��!F�r�]_�Q���Q�&��׃��
�z��6��^�W��=�/���?�:�^�A"�!��Yz�Æ]M���H�f�{�%�0<��r��5*��u�C@�t�3/�p$�tC��K�	�#���m����1u&�qQT+�mV+��q���ߓ/���:��c����j��(w}��u���2�h~k�y�b\MM=�Ho\�0��TA[}�@�g��­�t���ZUF�*A��fx�}��y�.��M�V�%M�l����=�p�n�.o��&p^��&;{a�jX�9{UeΟ��͕�o0=�������'�H��� +�FcW���K�a�ثX iTT���Zw�	��Å>�"�~8�D�&d ����j=ᄨ����A��,�KC&�6s�����δ%lB~�V5U�Ua�DĽ��mQ�]a;���oj]�L�����<�vZ�RD���b�&#x�s�����OGg��=��7����yP3�Fg�꾀Z����w�W�&��T@�B^�њ <��3�<1A�лlt�o%,�7L#!���A�s���y`NI��u��S�.ʹ��QW&�l'D��s`�����3��^C+�3H�V���١��yy���5�dWڎuF��_x:b�� l�%8�=\2���ڌ�S�����'�\� �NܙƓ���fG7/�Q�����n���-�d�@��Eg\��Ý��h��;k��yf]�����2 (?#�|.x��Q`�?9c���׉� =���kG�)X�!�8�=�.�#�wI{�ug7���J:n� <���u�oƉ���N�>����� a��gE³r�=�q��/]��vS� �J3���������.]�t�8��ܒ�Į�,ߔ}g�e��ߏ�W�o��Q9��Mp16 ���!N3������.rf���f��+���wt�K�q�F���b�5]߸�#�s��S˞p�� ���<��!/����~��".�* 7���D��,w�s�e]�'E��ż�=�V���>+��ΕQ�/���>�u�O� 檖v�k�L�Ă&�so@����3�M�=��E�QW �㎵ ���z�lO{�5�_S�=��E�<�%H�~�ΫPr�3mf����d��jS���K��� �]��"���̀�u]h�
�w"oAw����v`�b��<��?p�iuLt_7�Q}���������F�~���`?F�7��#a�[�_W�~�j�}�/g�3H9�HޒG�loL'�'s��~tWRFYwJό���}����gv�K#��T!,���A�`�D�{���|�b�ؔ��`���ʆ�o���[�Aw���ۧ����/G[3���@�H�����*xTG���g_���BHj�k�$+ܱE;�׳'��Ij/FT�cxn/�h��i�Ď�;ŉT�A�, ^Iu1��+Dj��oBE�t��!%Q�7����S�Z�RZ�����%}̦)�j��ە���06蹞o�U���,�A�M3�J��5<�EA�S���Wp׳0pM��vGכ���,���J��o�B�]*���./x!���m��H���e5=Ř��h��A!���b��]�"�]ժ�;�\�|h�p._m_-*�D�sf�:�g�'WA��db&;�-�w`b_3KĜ��x��������#P�`��-S�a*�I**��]Na�f*������j����$w��^�����}e��Q��6��+�X�V�.�B���,����\��)i���i�#�O�z�[Ɣ�"��RS������]v��c1Y��ױ��"f4�e��_�5�����U��&�ƪ�U��5�}�! �/p:���yt�c0���7E��F�`����[��$0�/L�F5++��I���2ߵ/Z���,��LZ~M`��i2J���/�����n���D0NF3��̥�$8���{�p��=}~閍"��C'���Vt2�t�?����(��௥�ֿ�L4Rrltv�n%:��S��@.�~'Oh������ ��^�����t�2���}' ��m��8㦐n<�2���Q0�:9���.�b���V�M��ZĀ�B��\�?TE-p��T2�/��I���6�_JoUuk~J5(���K�g"��@�&���$۔��d���mgի�|v���3BA�i�oB�BMȆ�X ��e��1�� ��
���^�H@�=@ɞOрJ�*	?Ü"��>��1.�}''�e�b|?��Z6�yM���0��<������w�mި���9���i�WVQ}��KY���x
D�IFt�m'2��i���攴�&{�0,��/mk�7�	�K}�KE��
���:�2B:���i�l��B�i ������"w�Ii1~����c��CL�@�]E9h��R�fQ�k����'�p��g�P\��V+A��F  �bE�|	��.��:��Ը�-ȗs"�P���!�Źo��!�0�nC����ǿLz��
��М�|�EU�����x�j��%xE���!�Aoݧ�7i����Z��y	o%�J�,�t��Dm�aeD��ʾ0h-p *"!r����S�9<���s�����my��)>�;|���,���Ve� 5"y�f���9C"fş#�L�'���8�����uGæ9� �̻Ϣ�M_ϟ���!�0���݂L�^a�/���~8nM�[/�b���!�L��E-���������8��{dX���mf%7�oۍ�#�@a��ܐ�% ըZ�R�uJ6}M�X�}��H��ӡ�
��� ����A���@6�sQ��C���˚�l g:`��N��t�
N�z���!B������|%(e���V���q��23U]3�d�Q�I:y��4��z>Pݜ���y�3!�~���))������Ǎ��eB����bs#a}��M̞��Dī�~�ֆ���UF7���=]��gz��U�,��;�.o*���=��#��M��j�h��-�+X���Qy"��W��v�X��@��j��oE	�$���IF��4Q�-:㰎�ڶ
;:��N�\��/Գ�Ł5I��/z��b����w�"0� sZQE�2t��L�۾��f�sW�a ��Z,oK�5�/��T+�Ɋ�0�6�:�x���읳"=�Ԅ�R3v���Վ��{z1�BE���\NBQ�� �K�w���ɮ�4���i�dÈ�{�!�Tc}�&�7������
A%I�� ��y��규ٽ�Z���	>�N���e�G��G�F�{!�C��Ȥn����G,4�4����#*D��zg��W�`��?�$0�.�V��	4zg���ōv�ll��ZJ�.�0e�÷fvѸ����9���6�/�����ь����ɯ�N���[� iP%o��sU�/��/�h��.�e����%y��O��'��|4����Zo:����MJ9N����Q���h ��
�,��~�#QY��.u]ڎ�:�|i
qO����Y�	���%�{}����QX}�ՃxuM��uxFXݎ��ﱇ����	U���Gҧ�jp�0�&h��n��a̉���M�+ŋ���R�0�M�4�E�QC����:��-�(z,��F{����S֧�Eh�tڙHg��i��"�����=�z��FB�9n����B
����*���S�<�"�
�ţ����\I;���t�&E^G���^�1�/���i��M�9��/,��y�j]��`��p&�=��4`|��r�O��8邟�M�/��`��^��u�@��eEC@��}�?��.B���V?q7���J
mጰ�]mߕ�sD�!9��-+f{U���f%�Ssa����I���T��=�n,�i��	cz,���@�2 ���j!��P�/w_O���9�v�]=�c�lZ�Ft���X�2�~���J�B������.~�Ut�E_}x��8�W��j{@��ႜ��IE ��C,�a�7hO�qhu�LP�d����ӗF8E�T2�jwc|%A^=&��_������^���t��L��Z�Q��ɥP�n&g�i�f=�F�������r�j� یbGsܕ�J�S���Y��OR���yLr��'�����D+;;)hh:YXTq�YH��N}g`hh��B� ���=�ŗ�Ĭ�E]�z�����s&����9c0,�o�����t�i�
����1�pKO�FZ�`�_���B�-F�/�a�M���b%Rٳ�W����0l����V���8U��3h����vw�"�+��G@���G�e����JH��7��I�vK�~���T�5���W�~ʦ�ì��R��l���� L���,����$QM��KW��f����մU��)KbfD��w3�p�3��2[[������uHVLJ�R���,��K�*�U��ܲ���`�yxHf7�|�΀ ҥ�.{f[���x=��ëVQ�7JQa����|���?W|y�*�ێkSĕ�:m�zo�^���w4�v-�ѨP�E,����%���ڿ2O�V<Zzs��eZnO�5�;+g[��P��H�E�����B*�����f��!N��v�6��~���rˬݞ��*��=�~6&�RyVf�^��t g��g�|�� ;fX���ѥ6$C[�̽���H9.0d�����鯻�0F\A{��#
(�~$�|Z"��)g���4!�4�xw[��xb��~�sDQ�'ްP�%���!_��r��B6:����)��|1=�h�*ꋵ~[|mJn܋(U�@��HꟌv��^-��֘��ޭs�i��ܾ��8�����l�Do�^��bk�gQ�ݧ"�C0���T�ʹ�K�F�a��
�∊)��U�j��G�אd˕*B�5�W�r�!+�z�0#p��ZOq��a���Fc ��ǁ"�k#�FJ��@a��:�ZF�Qh]��Us-
e�W�e�W�����N�"i�4�a�Q��f�Z/w��I]�bP��ҿ�2Q����IA�:^.ŝв�)���M8c�D
��ɾbT��J��ùIn�i�����u�����(�}4f2*9wW�/ɻ8��8%_19+��Q��#�7�ǞV��~���Ę� yę:}�i�X<�+�׮>Kjq���}H�h��ߩ�v�g�����u���U�WH+�1\y�����ŗ��J`��$��fY�" �ݾ�� P�}I�c�=�N�P�S	��U������Fk|�g4[�ɐC|<Z�ѻ�����ݴb8�s�H�./��<#������8}���Ǐ�m$������X�J;��2 �� ��RGy7$A���OF��T˲~��Q�Y�F�K��Cky��x���0�t8\)���	�x��Mb��|���r&���o��%�G��zO�O�\n�$JI��c~�����|Y�>�9�ck�ITx�5CAƫ������� ��g-�49�ZEP7_�w�vh>V�$xR��Xi�t�����F;����˽j��\���@�F\p�n�[e6�6DISӛQvM��x�Q�YͱGX�"2��O���Y��R��� 6C�	���9Ŕ��|G���SKͬN�)$�M䛨�ڕHUM<�K�����Ɨ�n�Ug=5���P?&0��X�+-�b�FpM�7��<>Z� ���2�-^�I�����X܃z�^�W���&С�6;��j�&])��KB̲������pJ=�
P�~� ���M4���t��s���3Ol�?�U�ջh��v�����2`Cn�f���V,,�"	4�Wg�\B
y�?M~���ne��U��בi�L�=�
�O���$΂9�lM���������{$�σ`�Y���Ϯ����_c��(J űL<�Q�۩<[Y��V#��9����L���C�����M���`�m*p�/�R�68L�m�NY�)? 9�l����M�!� s~��i�T!垯�J�v`~7��:��'}��{����Ju:��CO���-#K�$�YƩ�Z-�*q�$��vN7�;~���$�����13��Q2o�����4#s�l}�]U���
Ԡ>����#�^��/�J�
�y���-z�X-�oԓ2�e��5�Vp^����p���rIrN#z��#ه&A%վ�����ُk�+]J��AgJ�{\oA�&.A�ֵgM/��d��Tٚ�kQ�$�j�+%3�Xõ���i�G��SL���r����V@��4�͎Ѷn(��
J/�~����t.���U[�pXĤ�Y�뷷��2ݛ�(��j9�gu�ǸN�_gB� �� �;��yݬ	�H��2�2�
��d�>�:��y�m�d��k�=�jd�v�V�������X8$��'F�&���{*��']>/8��l *�ZRr$�#ȣ/�����&��<�W��A�Ld�v�P8��mg�W���Y��L+�^�Wf� �%'�} �s�����m���%�M&�3�{��ED�Ey�W��y#p�c��l[���G�/�\<���D2���<�oo��a��J`d�T&=ݠ����ź1��e�=9�߶�4ᱎ$QA�>ʂ.�K��½��PL:"!��~�S�T&���IB���:<��c�p��ސ��j�����\��V�jЄn�8��e�:t�m�[�p��x>V ���є����LǦ���ֽk,�f�w`��M��>�%��ӹX�}nLˁ�)�RFM[��4�$~>WaPH���g�n��s�K�6����&�G���3�.{�E(�Wͣ	��0�AN�l}kOyX��������:�s�b-�`i��<�b�-�-�W��L�5_�ʩw &�&����yq�\��O{ I�)������/0��1g-�W�6r�mL����N]B� Ǖ����{����d�����t��<;�V'��\��!%� �h�.gӂx�I<4�+���R@gs�{�)�[�MUk��`�%?<?סBuA8�z�'�P]�G��m��\��"��!y��~�[Կ�`�?B�@E)t $���x�'��E�z�k-|�-N"PNBtK%#
�!��T�>�`~�5Up9���s�I��ya��)VG�����У�Hq�/�}}¡���V'6d��-~FVv�1�@,� ��A�(��G�Y�jjx����U����N��kWU������InVŚ3p�I�|���ϋ�
�H Dvm�� �Jx:��ȼ&�C�v���1�a����t�S&1�:PTu�vJ\U�p?<�X�:�j
�;�Ȃ�r�|��˴�:��&��'L�(5�j�~b "%kqi+<A�^D���B�x����Ɋ�2��l������(ho�Z2��Ι�(ߐ��d���L�X�.��"L�CaO��VhV��lT!o�� ����9~kba6�犔1uԭq�C"�e5�Tz�VUj;�%�ї�x��6P�ܞ�S�eN�����+��YuyÝy8]�B�}K�V%F�Δ�r)f��wS�1�&CtY�1� ������{T�E��X&����bnø�)���(��u���P�d�3�	�c!���Ad�#�0�������I��;4�^~P��9.��13_���U�d�4!rI^)p㟌�hJc�s��K�v�~2�ꫡtșv)�m?b�s�!&hVN�۬�!��&���TN�<3Ur�%/���+���7��F�@{��\��5$ǳ	�p,v7�-Ԑ�R�͐Sa�y4�?cg���Ib��@y�C�W'�ȭ�׈K>��-�>�6~��![�kj3ܾܸp��E��N��K�� �N�3Df"Ҭ��W�*�6��_Zlڀd��A�Aټ:��W�$Yw>I�@������He� �зd���,��L�z����������;嵟V�"�I��ʧ}yє
Vw�j�у	�b���+�վA̯�-:$IX�јb5c�X�$��$SAM)j�vZ�@5E�Gp�[��Ťj���~���q��BQ���D�A(���4�Q�d	W�GyƑ�0�:���P�����L(�i�)7mtNU+9;�e��3���Z�N��ύ���eE�	
}@��NR��KG!Y `|A��w���$����<�lHx"��(�rF��7������-!+��_|�K-�����
35�K�[5��G�°�����H�Z4mOV��Ⱦ>��T⫔���q����C��|A�Nb�?���dgt%[G�|`?��}O��.�ך+&f��T+@��{Ž�Q%��`COTfٚ�"����b��X��Gwuczg�{TF�*�H��yV����<{��Qo��֪G�&��\y`�����N��:��Q_d!4D��m�����idh_`�y�.�eħ=��Z?헷���XԪ��v��)�������?���HIL���3_��h5�vGn���Fp�V�'lg?��+F�_�w
�\�ӫo���b���h�Wj�=Dє��u8S0l%m�L�V8Ȳ��4G'c*xp4�h��;ݭ͚G5ʤ&x|d�@1ԳYb��&o�ua�����'Kz��h�-+�(��~�_Amc��mB�����b��2�k]�?�K��D!�T�d()v�\��vHXtIC'(�MH?�2L5�J	�g��:�zk����`�0�vYpO_w�]�\瀕�mb{��l~�m���%��H���z�
j�h���#���
��!K�DdB��/6&���OBAʼX؜�3>x�)?D`�n�h���~�;Cб�W��<�Q����r�ϋq��[�!D�xD��&~�mV�n<�=��ک���I�_`�H����F��,�����BL�Ji�R_�����T{�!��&axUPp-�ﴓU��R�u֠`"���<
/�Ҕ�����& �N���hFE	!�nn�����9m��6��Ep/F��l�o�E_g�z �;=D, q����ڑ�I˽��GgCp�
���p��5�q�n�刓�J�鎜>m4�7��6�P��4�4�~q�0E�O�*Ng�ܹ�Jz���/���DC�)��R�e��b�����
2֑��'��f^��`��ۏ��:B����*Å�y&;P>��zl��M8'�y����]K�*VtF�	q.�m�o�g���oJ[ܮ>��fG4�:�E+�O�<��A�[�S��RҎ�ie��t���x��B8�f7-�֘����V��DGK�W�����t��-kb뗣�?��P�H�Ch)Pn���N��ۈ�e�C�ṃ*|(���k<C,Z:� �G���O����	��6~[2r��ʮ����@ܙΠ�^d?S{u����a�&�S�R�ixe���+_1CI	�	�K��~.:�&��($�#�~�oh�����(�]1`ҼVR^������!�k�j��nRa�e�L�����Nv�pH�);���� o=�a�iK��MA���0����h�Ѿ���Y `�mGA��i�t��6<viH�w�P:4W�UzV��d�Ee��)q2���'I���.����+�xy2{��K\�+���a�Ip��(�0�!�ڊ Z=@��R�ׯM��( ǵ锴>|�� ^j�f�4�w�UZ���t��ސ�r��j��Q#�Ĳu�6��ڏ�L��j�JE�*C�tz��hȜv����ۜ�WW8`��#I��2#}�?Ic�Z�Pξ���A'�l�U𚿰�G�(=
�z��+§��@_6��Oy��.���(0"HE=����2���=����<.�`v�Y��d�0{�.|�oӖ� Nr����K�#�����)���~L���Z��_�,��k���b���RT�c�vg=@���&��̯>�o�����IG��OM� q����+W�`��k�ڬu�x�O����4c O�Z�LlG��Σ��͇��8E��������O�mA .�
)�X���h��C�pG��K�FTV�C��/�kND��5e����q�L?\g@S.�^����f� �q��x43/�Bzj��.f��}�*^Dq:b��VUi;��Fچ���I��u��2}<�F~"�!|dv^�bڎ�{�#`&�C���`Ī�*��zp�fƋO^#9dO��}/5x��q��*�L�ө�b8�8�kNNl1ļ�Uɺ�cH����r�˶Il6NJm�W����+��V�U����95Tuw�ꑖ�vX�ԧ�aGj����א��t'O[���^�?�����"�<�r}.�Fg�c�� �Y��_������îUfpc�E"N���-�v��F[V����/�+��(ɐ���`cӈ4�v�(4��f=�f�,�lؙ���"J��-�!�u���R�$<�J�'��$Sy��=8�P�����O���b)h�Ks��mHC�ϼ(����Lw�o`�U���ߝ�t��/]��~�슄*���Pف1�6T}��𯂷�����&�����Ou������i��(I��Ov��)`��{̠�x�ѱ�MB��#*z���~���H�^գ3Kʿ]A�/��_V���hǧ��PjdM��1+��Z���*�옫w�:yƻ�7�������
cٻ�f��fBMM��*m��Ű"��x���s"`���]�X�}����A�-�(�Q����Ʊ��&�F�`�1��W���o4=���&�q��J�#o�H��� ����i��+���N�4%��l�3c����8�̞��Rf[�k�����ؘ �t\C-�2���[��UYͨ-����"�U'H��+��B�ޓ����2>����Z�%i��e��%N���b*��uF���p�����J��]e=� J� �����q����A:�_���+�F�ͪd�vGg4+���f  f>L�[FIo��R�Y��%3���[*��R �E���2ǉ��DYN��� �D!�	����ʙ��,t+�H1�y>����l_�x�YI�D��e�y����u�'U���~���|����S"���M�+_�<���ʛ^�)�Xn���_������;����fA˲$��h��S��o+�۬*�t,x�h�A6j�Y��F��,j�����/
�>>i�K�ҁ��9&� {;��?�)�/]��M��+�f?K#�����ﺨ���+3���:���h��T�S���YB�`�� ��G����|�N����R��a����bo���Q�	�zN��Q*�X9ۧ�<��A1�#�;�˟���x��}Y)e)Q�Ł9�a�k���~�c�օ��ǆ��ů�ET��b.}�y_{���4��zA�ߎ˵��-<�?�J��<�_�J���
E��I�
�E�oot�4	`34X��[�Pr�H�8~�!����2:cv|�5�+��`a�|<�z�$c�����p�;�o��*���ϣ���_X���e�GZ��q"s�T�*K�PcxJ��}�,^M� "ʷQ�E�=\}d���|ضvO��|���f��D�S�&�W� ��)��Є ��/��T�ZaGwaW�~�7��$7����%��� Zj�s��B��e}ë+[A�����|>F���oD�3�Qi�Ы~&W#G���T��ԯS����ͳ"e��> �Oğ����%�D�Ү�+�4�M�A�*�Ra%լV�r���Q�Wt�G[��zVb��dh����0��F158%��z"��G���T�ֆlWsƍ��Wx��Hmއ,=y#�����^60��{$ٶ��I �Wg��������ו�{�N.�H�J�a,��k��m��ka>�7��q�5Xݺz��lp����J�\w���U�O�mpg�:`gc%���7�b�M�u񻹟q��+��;W�M���,B��P4%�'^�SH���0zb���_ד$�tq�~Uv�&*w.�D��Ҡq���N#E{WH]����5q	����Ƽ�<"���T=��2�H�_:,��C����v�e}bR�F	�ٸ�]�0v�;��'����f��ad�<��{��DI|V���A|3��v�ϴ�{Њ/偋�&HL��{�����*���{�tV���֠�=���գJ�i$Q��a�<�
������O�$^��K���%��D]�x=��A�<=O0߫�w��hcrX�<h�k<�$w���&�V�Gz��꿌�7��'����yְpsv�߃L��Rv�����xu��aI��d�=���T���\Z���9��̳z΁���>��ߓ0�J2D#�2�'m`���l��ɢj�Y�3A���|�cpL��d3�Q����a`c�`�xN�p�_��;��萂9�P ��4���r�K��;�u��wV�.�<��x}�"�������"�Q��+�r��;��(�qHA��gxv-���AiMY��N��x�%��p>�L����z*%Cx;m,�ʢ4�)/�^�a���_���Z�@ި~O1������=����@J[6Qsl�7::���4�����.�Bn�|A
��;�3hl�ܿK9��� =��s�)���E���f�H�g��;���w�ʦ��IWP����bEU��5ʙ�'�)
@wy!�����{1͜6m�$ec|�� Sw�x>4?�P1�����D˨����n��I��"��r�>��ļ��s;����A",����V�l�ג��z�UL=)b_�qbh�.�t� 6g������B�e� "����h�O�*ϐC��򠳭�>M�mt���U]� No)R���Ͽ\Z�ƒZ^!����,A�["R��N��R[K�������y���	mg�"j� 溽���/J��0�m�B�e��!,� Γ:��C�R4X�4'��s���C����Ѻ����K~(�ȱ';n�6\�U�������yTu&5�J�v�@&��w�-4�K�~��<�/4�ϴ۪�e�R4�/��,��	�k������Z�2r�B.HN����t:�@z�ҋ9��?���W�yu�����o��7�ƎetI��/��ܱ���Z7���_k�5P1�U���#RL�m�?���V�^*I��%Q�So5f���ސ=�����Y�t��|e��G�����$!Ҧ��qtj����:�D��G�� �Q�!#�1%�*n#u?�` }t�uR$,�BR�폀��'�8�tR,�4�%���e��� ����|~Gg󴅾������yi[�m���yJ�+i�R8��D'�Y�ǰ�N�H/]��͟�����}���a+���l=�.'f��o��Ρ�*������P��RMI�Y�������AY,�Y��ݥ#\�g{=���]��v�6Z!��g�D��ܢ}i(�<�9��h�]��z��r�|�]r>b�ͣ��{�~(���'�G�C��sfS)�j�.Z���#0d_�d}/ю�"����+qp��	/��q�Ek(��(D�*� R`�/�����~2Y���W.\�LjU��a�)�N#�B��#���`p^����"�ߘ0�\�t1I@�e�Xک�(!���y9���[��e���/	�:A��&[W6��\<\zo��S�&��@m����4}]�p�� oMm���}L�=�mN�*I#�S��#������h߇uN?^{{�ؕ���=�y>Uu�h�2~���8t%�c��~�M9ݖ?��D u!�D��m�Ѹ�(���� Ȯ�9 eg9V�����7�^�`;�҉A���}0w,[z�n��Gӊa���#C7���z8|$U'H!cA��0�����a�i7Xܼ:�V#L1�����kT�Q���o=�Xx��J%���F��7#Yx���.d���6~�*$�G6�8N�W+_9:yә)S����B�t��2�	�M�	����j�J�/ls�@qA��&BM�87+�����8�w2�N�h�ǴT�рY��s{�}Z��5G�R��Z
�$���C�%r�=$"�V��A���WO�����`i��"T�7�D�9�9���r�Q�� JM�H��=���e,1+��W��L;q����G.�ݙk����7�.$k���G��qX੶O���o��9j|�y59D��сIQ^��E�Ĺ~��O�t����ݑ�x��7Ī+ES�)�ݼPȵ����YN�Έbuj�����ai}o�e����З�qq����! z��T��z�f̈�#�S�=8T��������8xVs����۬���ߒ�엕j�O��A)�y��e�J�*��`Q=��\���g^�t��H_��(�_�ZK��2�'�X����R���5�/q�\Gk��x5qE.�� �����mU��D�о����D��䬠0���C���UCR�lo�*NF<?J�Tv9Ѐ����Mj��noi!��������a@:|j��$6�� ���<�\h���t �0�&L�a'�=N�o�os����s���[D���K�T0�`�\6�	"L����Kl��&/����Y�����?�YIŪ�w�̙���N���� B7���1��	���gݑ�Nh���e�6-)�'U�O����9�=�b��ԥa��K�F8\T~o_LO���sFz�0$@V���^�g��Wz��H2��.��?�dO����3yM~m���tal�ko��2&/�)��d`�<���σ�2K����/2�ǒ�0X+T)�C�>l�*���&u4Hƿ:� ���3$���t���1*� ��y�eUؾ�XR���p�⽖Z��{�3@��@&��n�A��o2�ɴ�Nz�Q��o���<�[����n���`F�/h�k#���Ej�#+΀�r��\�"���Uz�`�ExDm�7=Ld��9����U]d��8�  A9�TkfE0>|����E��c���A��/�豙��,{{O����w��bז���T��v\E��D�8̭]NW���y��9Q�Q�"�~�����Q�m5�<6;�G
�ȔH�L	���%�5n#�~�@r���|@:>v\Xw����0=�q�38��4��/��!i� A���|��<,���7�5����O�n��k��1�j�=#6����:�.iC�}�%��G�t�`�F.%8.��!�0��i&n�/	��	׊�� ��u
�'Si���$T�V_V�?��V�����ܦܪ�����%���b���q��?�4�K�@�*�@�
�h�Pg��ֳs�m�H*c������_�j_��JJV��<0�lc�O�#�RUt��ȡKc���E�*r%d�1���JE����=Mm����/@X_h������$ly��˵�@:���)(��`-�q\�%���x���D�/�q���B����9X ����W�\{�v�˸0�Kz}l�`�7�}�'�t��)'��0��*󡒾O�%�f�?x��׃"1"C :#d��� ݩ>q�/pK^H��'���Q�`;9�G�����_�9y,��:U�o���Z���dY�] ;�X;�\��gu��^�ܲ*qܔ��1��K%�\X�+��"�� S�r��NC�0�V91W���5ť�a�U�;~�h`@�����7��:��]����ʦ�{��a�n���!O�Ӌ��P;�<ɖ�U�Wd_1��Ѐ�}�)d�Z��o�h��(+h���8����2Y!)4�M_�t�:��"5]-�*���H�g,X��ܥ%��K�CB�M�*��� ;Bv0w��	���0u(S�����G��.�QO�h���<���ƺ��]ߍ]D_ڦj>)���R��7����Mm7�E�+�E��u %l��1fJ�9����Zj_'�:��A!c�����=F0$l=6���{W�SF#�� 	&�|�i����x�%O�EQ�C��w��F9��D+��Z�zp�;P��a�p:��h���Jyk,���@*�7i�C0��%l����sC��z������������ו	&�U�L�b���93t���~Z�5���$��=o`/��1b��k��|�� �\Xs>�ғ�l��~݆K�P���
Z�!g1�f���QbaS���"�L5P�e�+o]�("o��ͧ%�Yo�5�l�@���J��aP�8瓺F%d%�G��=�:��Z�(�WQ�j� �),��|'8qN��������E8K1���t���6%���r��	�C�?k�*4;�Iߐ��֩�j���:��#u"�c�<�R�mջ�������g�Y2���o@)�<�c�=Ӂi�v/�b��J�~�O��º����<�j����/;D{�nc$ԃ�Y�{�!Ƹ�"f�n�G��u����"8����N֧H��d�6 �m,�&;:ߢ״���$�ڮ[z����ʡ%}���5C��]��z�Rr����G-ќ�ۗ'���OOa�S�0�|-�X���������Ez�:2 �{��1Y��h���%nHw
fFZ ���7Q�{���R[콡iC��ͮ���f��kt�|��J́t�H|�d�ik���.������W6@k��a�����TKTj2y�(,52��& 4h�Z{��ew`�5�s��^�XP�Mf5�זj�S�����������[��^��X?�D����haDiH���%0�EvP��tBC�r�%��^_4�%Vj��������{�m=
&l5q��_��R̆��M��Nh31;��f�zO+>��r��s��]����m�_O�-��Hh��)�&�����ʉRY�
�`H�h}O�������ޢ���M&�y�'_��c�蹮N�T�K��$#U(�����8�?���*�y���I˳�������r���ҵl*���$�U��Q��^v�$�tM�����Y�끏#��ZP��Tb��:H�c��C���f��6yk�b!]P�LW�H�D�a�X���G�	�z�]�&Vf~�H�ܲ��kZp�����kR$m� r��$-�c����lz�.�wBJr3'�:Iy���p�D���S�߷F$	l巨�p��k�J3+�s5��2���g�E�tMq^�-����i�`�y{�>�.��+۹x�;��k
c�]N�lղ��i�]��p��޿��z�v�f/Yf��8Z1�n�5BG/����yf��Af��<�\; r2��ag�d?�w+��Z��^� ԃha=3%�į��i�u�8��RA�Y���-��w��z;	�b{t��d��"����:B���|��
"H$��eZ:Ls�Ա���ٳ�2�Mp���Gĉ�*%�d�^/ҠE-��}ӎ����WL6�N$Q�3� 0�ı �H1�7嫩eJ�Y�!�i+�׉>�T����Z��f>^2��R��=Hm�i�vPR��,^��Np]��U��o|o�&����ƪ����{d�h�GT��]������R_Nq��wa��xl�Aj�Z�	y�,iW��새�*�a��3���N�BFC��l��vM�hJރ3�:��~���h,M5�M�I���2�vz�S�b�@���w��"_�A��մ`������YR�^,G/D5{v�?e5a��}�k����]�u�YmZǕ���$%-3L��S�7��0�4��n�-4Շ�����:��K1e+l^%��TH�d4�u*���N�r�A=���g2�A넬*��[3-�-��j���ƃ�K��u[���P��\4+ CA1D��X�#�,"�ZJ
�٥	Lʆ��W���.��n>��;�(���p{j4�ӣ��%����ЁL�l+O�Bk�k��2$DG����a�D�v�'���T:��i�"�3��&@"�I��p__;�X�h�0|��5���&���d�cVe>���ȢKqB�-��ҽ�܅���K��F�� ꊙ?�:S��8��0��&�(�kt˭�	W�@ AR���~�p�C�$jͳ�Ex�C�߭L��^�����a�B$��9�l*��X��L˺]H��)�E�ݙ2��ɪ�lm�)�m$l�p��~��һ�΍��+�Q�|(��~��~I�ܤG�e#d�ku�u�n������PS���Ȋ<d�0|＝c ��C�_�������ܮ��7�^6���s���]�K����⪍G���t1������Х����W�"x�������{�E,�ͻ�h �Ҷ����`P�ܥ��l-���&������B=]z#�������3˿���� 7�!��+���2�U4κʊ��a_Z�ųQ:-ˑV�3�x<��C�����v��T-�S	d�v;1U�ٕw
�*�`�Fs�(��ɵ��聧�h0�@�;�ݘ^��|~�W(�^)�^��d�䐄�2h��d/�hX��]&��r�s*���T�����:̙��;�s>�N}v B!�38�)����9�-�O������xsy�}] :�1 �Ї�c����[KN�{�)Iهmx5�/���h�� ��y�NϽ�L%�Q�1��<ri��6�>�c���5K�r�	�A�d�;6�1#y�mi�c	�|'��=�E��Y?6�#æ�bNb��^�`Fu��؂&�$���7 �+R���2p]��:�$T�y�}�l`E��A����֢����ѓs��?>�bvM��"�j�#�ض��MV�"4yF�̴j'��u3�kU��6S�'�<�n�t�����Ǡn�<�J`qpK's��gE��As���;e�MB�V%D
�}eG��+��!�����i�~�C��ζo��:?d� ��ŋ��8���/W3������#mD�IM X����M��W�u�Q77+	�zS�AHi  �G��y+����
�b:�� e�%���TW*��a�E9R[LqSjyW�&ux����}��e�V47`��;��7�� ��O*NZY_�x\8��i�D}�E�ϓ�}��|���D漒�V���l�xp^ߪ�ܹ<Q��X�E�������;X��q��I�{�A��N�5�*K��hog�	[�!�7�O|nNs=�Mܛh���K�+�.�+�@nq�gP}��]��̡�U"�:�r�E%Y0Z#�k�;V'�����ȮX�O��lF-��Z+w!N�����GX�b��M�Z��i���>0˓��O�A�a�x`�`"ˋ���m�U:�&IZ���1���y��[U:/S0�l����W ������F�*h��,Ne�#�1��4�G�jm�����~��_��]K�� g_[�P�Uh��¹?K��U
�<&�ί��������vܑ����ǻ�Ti��xP����U`T(nJꙝ����M+.�m��"���e�
q���̂�o�wSk�rK���#���B5�2������F�~��<tyn�R-HD���^�*�����T!�l�@7���TOG�G�>yxd�<�W�.q�/M�~��b�۫�>�_m=�pu����L������%�[�C?�8<Y�D�%w�3(Q��wx݂ Q�
��V,�Pj�f�*._}/9�]a�3%x5�G.sCHW8I?i�,�N��/�.�67���}�u�V��y�ʦ��b�2Gs�6���r�n:E�����Y����6��hsr��[Qs���R�l����N�쥫�h����*���
�3��O�?YL�/m����܁9�xI�s#�Ź�.KPګs���ⶮ��'fMs}_�ÐE�Y�h���1�>��C��#�P��2�*ڛ��{���l�':�_oi�'R���4i�Ɩ����6ŏ�T�{��3�.0�I(	Ѡ2z7���{��^l?=�(l�Z ����X��Z[t̹����mU#��W�Q����U_��/���������A��gB��
��.��r2�;Ǌ�]��Qw6���\�nŌu�:�nY��J~f9��C$At�q���+�l��E�"�~W��lC��V~�!���c�!4Y�T�����ΛeUz'𗿩{�p,�[px�/eh��'@�l ���L�a�Y�@�i�@�H�a������OB�P[�]�L��'Z�n�������Z�8�b6�Uu��OubL�f�x�XӉt1I}��_��ʽ(�������9w{���	�r���/
���p~���b�=�f�@Ȑ_lvcU�i�C$�G�F��������k��x��ψު�X&;tF�;�!-K�\�u%w������� ��C�b����J���]�7�����
�	��	 ��������'��T�)��Z�ҡ)��i�S�S<��)�1��AI+u�VuY�m�J5����i��z�r�+6�K�ky�������� ��~M�e �C�E���
��-��	��0�)c�}��׉�X�w��íE?	�H��*�n*g��'����L\4U��{H�Gm~=EX��e
�Mlȏ�����K����-���T��`�
V�k/"��|��{�0��u�f0]��'�]��S��N�B�'IL<=K�Q��#�p�������>�@��D�g��|�X,�%$f$�\><�}�?P`Ϥ�6u+P�~�O^����d�$�����}|Qة�sY���Xk��3�}�)���#�S�H�T��lN�%F`��qa����]����M$�{�-�o�(fp-�#t/D�t$�ѯ�)w>*��u���Sݟ��)�,�&=�o򞡶�E2�׆�V�!F��1�D9u�j�vu8��������N¾�! ��hH�a`�)��u�$Q_P��k2B1��:[R��F �o��ʫ��Vhc;U��͌_Wt�e�,�^�����b�1������ᭊ�R������y��2R?���
$!y �ڗ�i@� ֢�f>���Єb� ~��*`2�{�E<M�B�%"Y��}�2 ��2ۖY��~�i��VND���&4�C�������oF]��6� �<� � $���4>D(��2-:�e���x���mv��/DݿPٗ��X��`E����GOm��>���~"KԖ��suQG�@���K*���ɫ�p�?�iU~'Ode0�s�@�c�F��j=��`"�x��c�� �v��� �����~�S��6�ʀ_��Ɖ<Q=x�� �e脰Ȣ��מ&r1[q��ʧ�����(C�h�//�h�=�� ��fI$ƺ���o�$�msvƼ�D�:���� ��%{M���z��/~�Ɏ�R��5��d��7������ ������K�L�2k��L��g�����$�xo�଻��5���$/K�d6�^p�?��D���'���� 6��y�o7*&��ˬ��U?����a�7�ڄ��%wŐ�)�i�+[b��Lq"�P0d�Uz�����ĩP����6J��ҷ�KW6E�T�K����|e��}]k�����N%$f����	�-�l���!��z�X���^�h�
�3���yf2a�|VZ>Җ0$󲽺����?..��%q�.]έ�.U��{&Z( �<���n�������_ǟ%�jXF��x�bJc��*ȏ�@����C��oW{�	G��	�ׄ�B��f�\�5V��*%���M���e�4S0&1�[��o]����v��'�ӧz�T��5w�1J�Xȏ��-��u՚��;� �8�_ƃ�Sqgھߺ��_h�+�fn_g�s\d<�"� ��6�k�s����Ȯ��Z�nS\�iU�4�#sL$nUآ�ʽY����Mq�f���6�ь���~69|��L��6�wu~c��BZ+�������XB����v�iFtS�D,�G�*�s��mC�=�8	[��L^�g�n���0ٿW��v�/�/���\�!��؈``�#q��*�v���~?�V]�$ζ[[�44U��hH���"����S���
r�E81�J؃��ui�B�����F2�Ro�	.�,+�&�[�� �V�0�z�s_�Ox�
��q�bmҜ�/��&��-B�G	���e��H�"� �n��Q�+����X<D�L��S������5�@�h��i��W�İŐ���κ��n��>L�=!L%�������G���\�����u�֏����].D0t�B\��h��9�VC,&�|Z��o�5N�!w�!��V��5��wx,�t�ť��ve(��6?�&�PC��!ۿP���~�
��X�R�G��+{P]�~�.�E&N����i)��{ ��+�/P�Fo��������<��	d2�d�a��=���0L��������0��2�z����p(L��ݳ�կ<:��3 ���/���`���ꮐ�S�Y"����ȟ
�ut�[%�VE4��M��k�H?���ӫBl��^�73[����4�ag#R�p:Q:ʖ{u��(��7���۸�tÈg�}�#�ϗږ�&���dXp)�QaVo��\S� �	5O��0�)v,�ó�Q��8���l.�f�&����0����,��&J�<.���P0�ͱ��#���<U��$��VEA2	�#��!2���K�����{K��9 4�䬥���]�}5a���#��
rIVK��a�p��#j�wiZ�&���Eǿx�R�լ�ڳ&���F0��ph`�#�a��	2��J����M#.���^Z�`�s�O�۶�'�z�F.,T��f��'N1JU_���O�D�L22B�{�^�`�mw�b �����Y��|�5k6�xCś�B�
�<xK��ƗR���_��䈔�Ar@�:͙2�f�c!q�C�E�:Bf��a��	w��ۓ�muJ��b�9a�]U���S_bN��*Dߦ�t�x���C��70E� ��ZBG���ΔB/����󺭑�u�1o�z]q��?��1��rO�<�d�v��!<`!k���4�)�-�Q%����sb��/.�1�Պ��B�⵰+����{B��%�b��;I�}��˶.�U'�쯒��l*���e�v-���X����y0Ep�*t�JuiH�RX��`��j��:OFʍ:��4�y����>�搥vk�|�������:v�l6�����|�Y�$��J���{@�%(��1�������h*|��q��|!�g��Ɂ�����b_����U�ogr.��5�*\�
�R[�vf��H|[U_qbW�50!��0c��pʫ��B�y���5�<���a*; ���	���!�P����S�=�ͯ�(v)�c"�~�Z�t��&~��\Γ� X8v.��Q�e�	7�d�=���O���Q�{�/,7��ُ>q+��!��w��c���"��U
2�?il!
��w���~���Q�=*J�b��>�'XOd��;sl��e�F���7ԭe���zHH�H?x��B�3<���$Iz��Cw�>x��FW /��.��>���6�'E�A?/:F*�C�=A�q���l�$Y�3%۫�Sv�"Okrӄ}���X���
,��n�Z���*���z㏆�"ŷf�}HER ^�M4�o��Hl|Z�3
ֆ������,<��7���iL}^�q��N��u���� �Nꇍ��X��Ί�2u`lt�v�E
� �� ����^�Y�r���7c/>�k�A�Ƶ�����*c�,WT�\�W��狋�ұEBh��H�t>�����K�����-U�M+� ��#�R9�6������b2Z��B��G(��ۯ|��U���ۈn��+:+�T'�׻�n3��`����f�啣w��TWR���YI��`��΁���9�}��y;����x���΃%oQ�Pd|�e��w����G������+�'"f*U��Q���w�q8��f��f��!���xuQnǎI��:�X"����Z�W�9kZmE�6�JEv��Ho'V���M�:	�.hq��S�ӻ��;�f��W�%B���f�l*;�,<�P� ��S��4u8zX��Jw6��g"��Ǥ�����O)�ģ��k/�<K�'I�&ЭW瀋;�{L=�3݂眪������A�mh$&_���Y% �|���	���R�O.�`�Gӟ�:Ñ��X=�����F�kW�F??�xt�o�,�T�T����I3|�
�ԯ*����aʅ.	$?Z2�cX:��|�w\>N�}��w�������0�ZQ�V(��RBm�N{��ն*"*���}����\嗢fF����
���㬖��䒍���ep�Z�h6��V��M3�=���-��1Ao�5p�����I���_�<�h��y#�_���z��]���_� �;�焮��8j%�e��)����L�̈́o��
����ш�|�,��H/�87b3�TOz?��V&���ᓋ6���Ej����܉�$��ai�����F�dуg`�W���2�A�cW�χDv�ȵ<��]ŞC2�Ư=vqao+�$�B��AQ8đ�a����o3#s���̂�ar'j&��Dx���-pV���2�襒9��w�*��&��E%n���ތ���y��+c��_悳��K'.[N�zhT��v���=��e�ŏ�����Əٯ����׭:@��m��뮳Yd�x�2+��"���a�&+�Ta����`�>U xG�b�\+}Ũw�U'�%ٜ4�HRc�è�w/�
��{@�J���	2�Kŭ��n3 Om`2��&K��~�c���n�~��N�=��HX����Ѐ��#���H�~�i�6���{�%�`�����搳?N'��=��X��[QQŽ^tfr���4��oڐ���+���ǧ��&I�Vx�aX�!�ol��3�o��'�7��7֔1_we��/�����I���&���_�W}39�}�a���Έ�T���-pc!xL�l�")X����L�d���}�)�Ĩ�r���H�U6��XY�dK>�͇�w�$Aޚ<R6� p[ܮ���p���S�.���O������Ky���f�j���)���u>[J?-m}�?�G�|5����N	�`)������@�:���N\i͑(Ft�kj��/Y�Q�ݐ��j�v�)�p�% vA9I��t�)�(Vk���Dҩ�f��km,\�����k�
�}C��5 ����ׁ�>��H�7�\7�hSɈ	y����$��ݙ�N����+���Ux́S��&P�޴Dڴf��/�-��ģ�*5���ar5$�m����[#�������_�`��[�ǻn��=N���4p���Q��ᔽ��\f������_�l�g�+�a�hws����Y=�f�"w8����_#fV�t�G�-w|�~�M}`ʉ���*���7&�jF~K�赩��I�Ê� J�<�9y#(�d&�x���ƌ�Ac����:�N�*p�=��q�Z5��"��#g����� �1œ�^�NOo���cR����
7�vq�x�c(�����i�2�����y�F�g,"�?�R�"�!�Ft6��ko^6�m�������o��T��Af�C�o䀤�H�j��o��I�ï�,r{�ȟw��}8֋&�j�����;R�m���SWO�D��q����eg�����rA?k������.�%��V�"k���а�?'%�����'�Zl5h�d;�;��)�&�1ذ�#H<�Hle��mbus��#�����"4J �r?��_�n�����Zx�m�&�z�ez]}���`,��˦& �i�,R�1��NT'��1����К#<X�oHJ��#2eU�ቦ��
d�D��{���hZ�F�n���vs0�J���	fS����DK^"�����͠VޗXK��Um_��o�e�J��-�!Z���|rM�ɎU��36I�wm��S ���{f�!fBJ�ՠ9��ude��=�ꆌ�;�OLlcM���C�����!����T7���#�DWx-��|���'$�'8k[���I}��s\�ՙ�~�ͨ���ug�r�{j`��n�50���q�:�[�@�)�8=EvM��;��7�Rn���I�=h˒ �I�p���b�')��vҡ5(�� kf��RG�NFm��,�������s�b�<�1����h�����C�p�X�;�0)�MQ���6����-��<�8q"g��2��3��?�3�B�jd�9�� ��S )Gxa(`'��R�=�� ���L�Ii�㔩��3�!�\+�u)\$��닍�K��ׇR�����娨�Yŵ4��c�⎺g�&Җ"��KxC�;/�@#3v��@���}�p�O����Q[�@ ��V��WV�T�+,YVL���t|J{�~2�ȟ��Y �X�K��j�^)O�ߓP�%���~�'�P�m�M;���*ώ�b9 ��W��Nn{�O��%D���:�l_� ��r ��4V��[Om���Xf�}#+�xW� /BoŌl��� }Bhw���@���tY����WC�Kj�x(��i�n��a?n6��[������z݉jL�޹�WZr�'OC&�L6�RD����)!��uC��i�A��ZOo�������l-6C�&vȓ*_�G�D�v1�@͙k���i��S���C{�yO�w�W��~B� ��V��v��Q����*������K˗"�"g��~��6ء��񋚼dE<`MQ<�h=Rl`��S]��Y�g-�� ��p�b����ʏm��D������)"|j������J #�s��VG>1�?�A}gjt��r`�D���Fގ��' U�,&�i�:���su�ruY4#}�d5H�~%�_�N��4��}�V�h��@9û��+8�|t哨�xt�4���X���֞���V��x���c@e��D�V�^röv�z&�39K��c3�-�@�[����MO���\�(��-R���\�8Lir ͚t�*		M��`M�: ����/�U�L�r�H:T�|`��������W](�v0NK#�c�h�g�WZ����i6���Kp���K�yjf*�2���t�X'������^�2��pl�J�LX7}S� ̟�<"w�����P�Dƒ��B̺��BEJ=�2̵Bz����}`^k98��d�8 �GQEe���&{gwA��ZA�l؄��s�����%��$��%,����A�O�-���E�t%����L������WñmDDhCg�r����5��G$ݧ�I�o���d�d��_a��ǝ�F?�����u���������<���{_�l>����އ�Y<����֖T��o��r�ܧ���T+��CܨM/}�OOťKs�H@���5�l8�?j����UywHλ��{�]�;%		c��9�A�C��(��k�P<��D(�.��W�fˋK����x~8��	�7Q�cf��%�ֲ��
X�8�h!$��YT�+�Yi����T�"���ț����,?gW`G�PMd#�	����^5�Q����+���zA�p� �k�2~����,�9%u?:G�#y�-dE-$���,\ ��X{0��Oԭ[C@W�#�a���UFH���t���D+e��w�{��.s��9,l��>����k���sj,hq����6}��M:V�Ek�HM�f�!CƐx�yw�"e�3���WɄ!�B���S�bq>c*B�p6�7�}�q;i���A��KG�=5Sh��ܭU�2W8�1%����B;w؃�6"�ە���b��*�~R,��n�j��Ä.˙�9,1��D�9,G�����E}����\A�p�(r���
�Ô�g?��/��	lU���{��&�ZW 8�3C�=�������gfL��^���YnS[����oN�Cyb�K��*�=贒T�+?F�� ��f��q���v&y��z�L�W���k����n��mC�.�h�uC�C�>Ӝ~'/�zԎP$B�T��@[n�@�6RrY�`��]AU$*R�=�K���O�q�naԽf�/M�����"�xK��D������{{z�D�O*�[r���ԧ|.�e�2�����^�.6D~H	z�6 �.�6Gs�
G��
H��<Uv�ƙ� �:����I�؀H�-��2�}����U����b�a��	bh��nOx5�������Q$�]�����Yv���
#b?>5����e�cfT��s��t�s��B^�S�%yo�8)���O�jP��L�^��U�q��j�@�e�l�L�:-&���,�%g�F�X\��麡 �O{#��W(s�"5C$����U!��u�fx"`�������T	��WhAB�����a�5/�njm�Σ���z?�u��t����^M�Y�������)�����՚-MB'�T^|T�]�ݬ�R�!	T��.x
���6�p������E����*4�� l�=P]S���� d4t�7W���ĆmX����d��^�F��˳�f��U�^w�>�2�/'=e�ڙ82}��ǆ���j�����w=��x��#�{Cݨ/�����������yrP�w;r>Ԑ�+�A��}t�H�@T2Ј�<�Qf~P�o��/��w7
B�K]�簳�[��b�/��U��)	r��PkCe\ծ���/_[��~.=����z@���	����%LTB����.,�A	�Ft��2��L8�R2�i��7?��u��W�ۯ��Z$��q����+E5��#�p��1�E��h0�p�O�&��\u�!@)X��έ�&�?8��p�h�ρ/O�� yn��&��cqq��y���W�ck�c'����Q��(���L"Ha����tA�F��8�A���F�U^�}�����C�M]�s6����,FT�L총�)crƦ�/�G(kIc�z� z���ܳ�K���F���!VFTa��&�NSi�� '��t��?^�V: �B٠ă�TrL���h�3��p�qM��b�g�yU�pb����[�Ӗ�p��tߗ�!�R�!_�oi���Ν�V�Y��ފ�^�<�\��f�s���jOꢙ�d�8���׻J*�`"����,DHK4Q�DE�\�p�q�?ސZn����Rt����9A����vR�伺�|C�J�E&�3����#a}9��:�;�HXe=�}e�����ȵh5s?^Zf���Y@��b���Tb��´�Gc�1��QK&�i%x�:�����zi[�����[���f��p�b=��Ibw���mX���֯tφ��t��F��~n¼�K��Q
v>+����,�Z��C�HC�+&���+}":��6B�+��b0R��c��@��/1������b��`�,����uch�V�1F�)%��^��r�ދf��&��uLk�m������e�H>�Xn��"2��nK~:�Js��wr�>+B��հ��	ٝ)�&���U}@�*}_hI�_��U5�,屛b�b���Jv��ݐ�W�7����4Ж1��{�;H 	�vv���Qb%�ԉ^��f�hߊ �5�~�rb�r���vH�8<���ّ��w�9,򼻃O�o��2=EkΥMz,�;=� �#[�wJb4�#R���ii׶w���hf}ٺ�UF[[���WX�'ŕ�i \
u��&gx_-"Rl7�U+�Qor��9��E�S?~�ş]�%�xC4�,xչg������������ť�ӱ�<JT�L�.����*�(�`!\L��d���T��*S���/o�%���y{io��[~בA�.�$J[?��`�$�cG���*�L�e��b<L��h�����b���S>��0U��i�`;&�	�3�KMyB�b ����c�P�(_��ú����FtR-i��MU!���J�&���0�(X� -OnW��.�[���.�c�Ĭ!Ra:m|G�o�b��J���I�+����8���B��d���i��=���ܧ``NR���Q/^VW�r�i@aS��O�~qX!���M��f~����]�9��6��SI�r��kz?�o�B!,� �v�px%�G��x��k=d�ivʮ�)��ݛ��Gu�<Q��I�ǔƀ@�A��<��^F��ŸN���n��'�a�Z�S�-!5�$�ƿ縲ǿj8F8�Y���I66�|�뼄8��	fӏJ��	�qْ�AnS�^|f$�ثA4>*�A�Uۄpj#��u���d)�/��^o��ob�;=o�8��Tl,YCN�h������V���;���ɗ�=cŕ{*i�$ik�����) ��$}���8s��R����q !��m!�QE_�#H�B�q�fu�2N��_%'���1+�fn~IJ��?^��u,똄����?���m�@�ҿ<0�F��.o����;<�3��4Rl������
��d�H��pֆM���D�NzKQv�=@k�.jDD���|�d��3 X$Ӥ�����ie�"-�w����?�Y(�:{¿�|
I�6x���Ųa�����4��kBk�y+0L!�6�����:k}�f�fy�~��s�ga��+8"`T�;�"�$6}��Mgb��K�f��t�G��<�X�br�*�t��U3���D��s�6Y�|�L�DbL��>�]n�'�@���J/�%�R
	\3U�oi�Uo����ܻF�ʒF��!eB�z恌P��C���>ѻ6af<�zk�k�vq� �I��1u�7�������d�������jʹ�����Cc�o}or���n�&�|U'�W���z��q�,:�5����v���G�+���)���;�}e��Բ�uXu��q��lW-Z'o%��e�ç%Q_�KFO��p>Ѭ��.C��-��I5�u���w�:�����S��>`�f=�P?�?��f�#!O�-Y�X�י����3�������.n��qЌ@���6�z�}]�c�6EǿO�<r{fNyi�����+�b�X�Of)�k206����=!1D6f�&ޒ��0��/��mƿ�>L4\���G�w�wd����(�$��[�~��9�F��*�j�ñ^^����!��85 �we'x�}y2R�%8�T��q(�q����[����k�ǔ���b�T�N�3B$0ã�Z��?�F{���.p�Zޓ�6��JQ@& �P�W�3�p�N!��/܇���������1f�b���� (�PB�Tf�kԮ�p���@��"��̰n�>�C���ԍ,�+oC^���t�{�����a�D�wѢv��ǎ~�5�D�ܶ�Cb!�81pZ���NX��<C:��ʨm@C��=E�r]no���7A1/�tpg�չ6�h�֘�a���S��e1���R�1��ζ��BF5�.���F�z�Ԉ��k��+Qd�N�F�:J�G�õ��pX�?�t}@���{@F���YQWWEJuc����]J+V�~�������BzZqN�]v�J��/�_Y{�e<�q+s�ܻ��R���_,���#]��]�e�����	Ka��x'5�j)|150��ן-h���� n�OyX�RD�$|_.R(�0]���X@P�:zA���QU���y���e���v3���:�H� L?���`=;�3�MG��Z���4hF��,��&���*���C,߭��+�R�\e"�\�5�i��#=��'�]%�0�"�LH0Ò:���!�
T��}�E/Μ����>�M�SR������O Æ����:�/5Mi_�Y�����^���`�1Z"#�J9˒��ݍ���|:]m��_̧�Qk6�?,��������������tߐ�.�8��Ol��?�I��I��ѧr$E&#�rWa&�7���f?+�4������,e�(��ţ25[���i��BlM���c+2�=���M��Ӷ0{9���d(Dl`M�d�7�!�Y����\nK	�����xDq{;GY���t��T����?5��:s
�ue�j)�a���:����c�D8~J^�Gp��R�]��no�\�z.F���⭸'HB�4?Ef."�B�0�>��:�}Y4�{���H�/1�kc�l�^^@:t��Y�̇��pvO5nۅӲ8;��FnmY�V"�X�)>���~��&��K���j4��X�gbC�K�#�MV�n����Z[��s����N�)a	_��p<��K�vp˙��-<��)�b�~�2A�឴�e}v���U,�}��+,(V]')����ᛓQ��K��N�����b�.B�dR���Yrٜ%3C�߃p��9�/ �o �N\����M�����$�����: ��s�{A��Zh״ �0���:p\{rrݒ�zj/���K��.��NX-��Ԟ��.���(b��m]�i��ނ�a	�s٦��,�u�"��L�J/pjiC����ד�����֧_q3��E/�ޤ�IR_!kZ��5jk�0G���Y�N2�n��9 4ly���Q����8}!��X�X��r$*Ѽ�{��t����f���w�Z�/�;]ͭ���'S:�����h��1���8�$�*D��g�i��?^�Lo�(i9��ڻ��!�3�u`a���lPD��5|��:�^wN�,z	ܶW� O�,�ʘ�6``��Գ6U��aI���wO�	��X��a)�}i̎Z1��!Œ����]�Umxq�1�E����Ҹ쵬���b�KޘI��%0}Ӭt�o1����:��K�)]me��~ ���Rq%F��֯�S��>���ySM$`$$��X9�1Ja���� ����{�"�4�]��V����O��K����Rb�4�bJ�ڧ%��j�\%|�I̧w��m���#	��d���7]Y���K�d6�\�r�gay�eO_����%��U���9�,��e�� ����	f_si<��0�x1�['���7�6�מ,[&��ZeȠ|�Le�Y�[X��e1���KMT ����S1b��m|��$�_�1�u[��c������L���w��>�l����C36�ƍ�&�5��Xݩ2�4�M ��q�g!���X�8��>f��߅k���҃[�|���HUI-��_�t�Q��50I��SQ<�?�p�nGN5�^I69'��V�!s�����ŏ�6N}k�ʫ�]��q_s��z�"f��m�^�ō�I���7��q�tA,S@�6��5���U�Ow�:�׳.���M�ȋ��`Y�@lZ+�5w�(���[�������'m4�ex�6#<z�^eЅ�:�"qX��4.�h��Ii>h��h��e�C��Q�� rn�����r�Թ){��r�W���i��z�w%N���[�ю�%�mU=S܆1�����3���_��N��J�S�O����d���7^�\?�=$��g��H�����6���@�dv���m,��{��.y�SbyJ���^S)�)#��_�sQ���u�Z0:8eeB�o�Uם���N�Z��P@�Q�*�1n�-��$�����u�>�)� �6�c��hJ扞1ޝ�ܰ��=�m'*A��a�r@��mPj��^�a�l���㵻?�/G�㐓��ް��0'��q��y��p ~3�	�j�xMm���B��b<h!�Ӷ�v�y�rI��Q�����^�DL�����@.�|�SD8�IT6�YM���� Tq�x��kM���_��Xah���Ҩ^_��Cۓ�Ӭ{��O#S�lf[�o���k�{����/�+(t�e�FOTe`�}k�R��if|�Ǟ�rTtg?�ō������`S�+�[�+��(D?����ٍ<0'����Oҍa�X��+�����~�!{�
q =Y���t�oc���VԶ����,mFO��G�%=�"�^`��Ф� ��cd�C��Ƹ��_<Y�K�z	83� f����ڤ#�|��A	X'�  ��5�ڕw�Lf��ra8�f;r��#y3 9mw1�37&�QI�/��B3���TG�]��pf�'C=���U����L�R����"�9%2�[0p��cO#��
gyjR*��pO��-�x�~L3N�D��)�@��Y񽎟	�Q�
���J?� �t��T�?�4��͂nR��$��/hJ��ثfO.
�B���8�F��I�0����h��.����/C�̖��#Ҕ�aa����T��Fә}J������"��������'n~����͘}oX�y4+beUG��1�2	WKj=x�
#�.#��\�=ؿl�3�H�C��`��E�{R���T�����@�y[��1Yz7��y!	.f�D_;���V��������-;Z�O���-I��r��e�����A�i0�0���m��#��>"����k���־�0��S���J]�ď�7ٲ�5�����Eb��$���_r�t"Md�S)��V΂��LE�����<���j��.���x�Ew���;��|6Y~lX�n� �������sQ� XTB`yK4B�(�R�^r�>�_|"z�zڗ?��%J,��l��L�0hUM'�
�P���}�F�C�B����A�˛F�1�.7�����{�u��7�5���ax��Gg�Q��M��'�����L;�Ą��+�Y:��n=�cy��2N�����4�2L<�{�m;�ݹ耰��~|�Ma���d��7������X�ܝt�$���膲�h�w'r��@ ��܉��.yC�I��y!�n£C�0ez`��o��
L��;�ցH����(m�0�����w�4�@9?�/���9����W�I����F7K��>�e�5>e�������?H���q7�c}"0L�x����hJ��v3�;%�A�U��2U-i�fٙ&�L꩙��%�Y��̠ZH���>Ӻ:1#�w����'���j�L�5��m�s�œh�`[aa*���
��^-��fm�f6|yʎQܳ����dL�Ah$�:�Mf;?υ�z@pZj18[��`}%s$�B��֥z33�N�!c���p��O�z1�m��9���FX�ɶ +�M��*/��?f�T��'���b�5@_&ߘ�<�����/~��D�#[�5Y��ȁ�K��_^��t����S�:p4_���[w�lC��Ꜹ���)7��]�sC:EϢ-�� 28���cE31�(�3h���eě����H���4�<9���9w9P�J��e�_�]7���˴��drzq��E�Ǔb���ӳ�DI4,Խ���!R��q�N�c/�䒑���&3�޹c$�P2��EI)o�- d=e�N���_Ƽ3a�����9
m8/f5��zu��1w �,���"�4�>�f���̝�`٠�����|#� �;<�]3� #,�! �`��/ۇ16��4��Ǌ*���@�o����'����/�E+����;w����1���:�t��_]F�A"_��1Zj)�]�
�DIF*��5�Y��x̲vt.��G��Hv`���n��4y��}R��Ӥ&+e�9��A�H㣕�,����]Zk�"��%P8��|�{���av�?e���S���Is �s��q���
���b�_��32��SY;��1y��q�8����c���7��O]Y��͂�0��U�G���T21xֹ!���7�]��{G�S@��N���턹V'E.B#�zUĵ�
�^�����W���̉[d�3��?� �{p؁#Ԗ��7z�2�Xê8�Nσ�R�T��̵�f�g�F\20Y��D���>�w�����cQ��{��Kf��?�Ǝ����m���ӽK�C��4�Ơ�	�nhZD~�52��7Ө�)���p�N5�ڸ�j�}~��d7`&��gw�+D+��d�b����b�j�Fg~�V?*@6k��x����{_�<��2#ў�#T_����Y�O����tD��z�dR�����3K��6�1�PN�56�k�/�4v&�%�VZ��	� ��-:K�/�>,�O�S�\V�UE2�-�>�f�į�z��������|�>�XX?+`e.�=
\��$w�u�qb��&��מ�"7�ҹ���q&�W�.R���1�
��<��J��=��|%���w�
����,�{���fT@�<�F�o�j3Oy �V�Rt��gw�����~�>[/��yW~J����B)\9��gt��}I�������._�j����
v܆S��q�U���C��R�����]�������i�lt���E�Ay'̓�}*���¹2�m�ӓ��2k���@e�>�\�����������9jL��n�ѓs����������w��LP�Y OM�lr�!��3�e��/��cj��	^3�������Rؐ� 	�̬$�����ȷ8r�&0�8@�n��@�/��a�׹�6��}��p�CG�ZM2W�j��ϕ7�.� 0h
�ۋ��T�d�q4�[��ʏ�xb�dݾ��8X�S��9�:���pE�΂hg*~��$���{��l�5t�ί��Οmk�k�^��Mk�9
���.A�Q�рu3���
�7�(}�˸k���?]lJ�Ǟ�����TH��	���E�+f%��E�ދ{.���f�ڊaAa�:������O�#<�X�PN���ϴw�^~5�����22l,ږ��63�yՍ��V�-v4��r���}�RmV��+]�;�˯��X�%te(��b�\��v��5czl,*�W�t��
t�Ԕ��2�qUq�� ��A�Ԛ������omT�����6�	���1Z�8����e�qet�l
a�­pR_~�.��36I7���k	+��`�(���#F����k���:s��6đ��Φ��5�j1�p&�4};)'q��f�� ���G*��4ю��Z߯��X��^Ź���9C�03%Ċ�=Շ�Hw>7��Z�n �ў�#��I�=�q�Y@�P�C��J�w$'}]׍����%Ą����n����"rf��L��'���!�~�w�	���b����>Wܻ�ƕ�`H��*[60|�a(*��n�/�E�T�e�vם?Lk���&��,}D*�n,J�y.Ƶ�=����
��?��S��q7�6�Bn�Q���+V���*�����p��I��6�R����gT�z�����B0s�0�e;�L�T��)�a��ޒ«�ݲs�l�Lٵ�z�z��RN�����j6�HF�Y�"�����V�+'�!7\p����#�{�&��L��(¤�Ř���Y�^zX�k5 m�mԲ��.�
����Z
��@׫'<��"�T���P0+Thc�紉�k�.|�K��,=z�t��S�I��P��G�����AE�3��T-���&���k�����%-O{��w��v׎1)� �QYm�5�Lb'@b!�se��̏:9lM�U}XqI�!d���S�<�Jܰ�<m��_L���N�N��e�;�����#�N���֬�m�O�tn�j�(F�I���A�pV���8->n��%t�C��B~�;:;�k�l�)��c�L�i�⭺�PU��I�O���Hؔ�{>�l�t[��)��jL�����o��7>2�zGFn(����f�K�����:��>���+���,�LHF(�'h��3,�i`�������z�s�9��Fk�,= �wg�{Ɉ*.
bG|י�d�< 0�Q�n~:�A�ʈ#����Ic����|x�r�P�t�� O/���CgaL�hN
>�YF-����&)�aʻ�u��B}lz�vJ$�n`�v͸�~�J�w��^����(��'$K�{�P��v�5��	�`0|���n� ����{�N�I�Wjl���K��ؠ��&�K*UH�X�6����B�ha�Q����j-�b��� ���r+2���l�X�L��/�lbႢ��M��E~�tz.�������.l����{��W� %�@z�2���@t��t�i0�E3�4X38(|�v'��S;�@H����i{9m��e�}�*+�q�n.x�{A4G-�(�X
X������ 
"��!�dѪH���Ii��W/ݲ���h1@ٓ�h�fr��?�e&?��RlU��T~��-[_x&��4o��ԇ7��J�2*$�7�8+s�TVX�F���Z�����&�[h�I[oP�O��������&o�)����G$S`�8ޮe~����IU5t��b�~��B;��θ��c�Iڷ^U���Rm	)��f��s9rⶑ�H����u8�g��h�e�����㚿؎<�@� \�����F=����<��ۢ�.c.��ߨ��iM�7���B^ �#�_|H��3�q�&dר�m�ˀ/=�1m��à�k<?��x.�و���v<n`X���> �}�󁻀t@���Z@4�D�*��u��~��C�bT�:Aq��umH���^�� fV���'w[�5�?��9�ZB5�i(G7eP��%T��ڞ�H�|�4�EB���Yp�}�[��/p�}������4��]��F�d�ӞKԚ�J�&�l���{�kQ�T�74�K�m����\����Ͳ�<�ϒa齷���F��;}�j���HO�m�%�!�)��1%�~�ڙ�zd4�B�b��:$x�%0:�+�&�;�(��j5��Ew�4M�R����� Z5�1E�	7jzQ閑ou)O@���xdwfI�B=W�쎡�A�Tmݒ���7�耠����\�jof�G�%KI��n����q'8ʈ[ܽŗ@���m��1�|�a��ɧ �'��>����AD?}8�ŖIw��Z����ah�M{γm�j��὘y�1l^ǧ�ckW���6?-�tQ��6������O��ʔ��Ҍ�X��e��v�>�S�8���x�ȎU~����oj���)�����5O� 
��,;� ҈�<��]�@v&S��R�9���;��~�y�[t{��y"��,��q�}��QV����z�x�q��+~�6����_m�����vB��T�̌�NJ�:f&��t�E��ٿ��>9r�4d>G��*��m����K�4c�l�۳hux��������'�)BWh��t@p�aJo��:���`�\?��2�Zu[���{�|WF�]u�M�!If��9�������Z�׃u��J,v\�d�U�+�!�c78�Q�|z>|�}�;�7�/@��Ŏ�;�O��_F�}����4^kj�K>/���~2�&�b���ɝaV��|-�}�W��v7��^�s^���x;�d��"e(�4%w��H%��ԛ�v�! �紼�P�]n�8j�yf�
E�)�~hN��鱜�=��ۀB�ɩ��P�A�8��"��3�9�;&)���up�br�9��ܭ��-v�r�����jF֋X����Q��^�y��>Ä ���aOoaWe@�d�;��]s*���f��Tk���)V% ��|"�Uz�I��؊�j1^,�c_x���@U��+�:���)<��i���hCYz��|��2�����j��?��d�'�U��N?!����+Mo��x���p����
^#�dr��*����Z}����x*��&m9���m�eT8�.u���!�y�P�=����!$ଛ��l���d���L!��@��*^��7Z0�k'~��xc�x��=a"+4�^^���s֣'o��i"���W�h1������=ּ<[:h��ҊF�k�A,���&ө"@&����/�U�U��Mt� I��'�*-A����Ԩ?bd<�P���8f�^��Q��L.P�>9W+�ʉf�y�xH�3j�jf��iW��况.F���$s#����[d7`�J��8�"�?b�؅Eu����W�L�DX�c[�Zwi~ o8�b{�?ˮ0��J��7�zy�	�l2��C�<�� :�U��0+�G��x��Q�P^��[V��q�jv	��>e�O1�8Ԑd�^�jJ�E����<8b���A��=	��R�n�3�TK}W����l�f� ��9����{B���?�8��p%{Kv��M6mF<�6�~ޯ"�A���%���"^c��ߐA�p�~���I��f�o����,Q\�1�|�G=VYĎ?�'�/���<��};"�\j���ذQ+�$���c4��<2`��5v���)/�����ά���@��$WWE�֣F(�QB��r"�Z�Q�0Fbv���}�O-_�k�G�W��Y9g�:��vI��֗JG��b���P���8��Vt.��f�a�ixa�샛�Տv��*�WG"����'u�[ɽ�����Z��N���b|ۀ��դ���9UZ�ꓐY����DV����W*o����hI�����}<��tJ-�WL�wܣ�hk��s�
�gi!�cMm<w��	.@Ђ�/Ā�JL	@�O���1NU�āB�lyw�j���@N���y�x8 �b�з�oͽ�rV�̘��&�ך ���f*���	x��l��K�lD~�J�^�ql,�E����D�~x��U6��������*����:Z�9�۩>l��h,���	
�f�K�!�3Y��Q�3�p
�u��ϵ���c�T��)�/:��*I��f�)y6\2=���G��Z,�)vΜ m��S��Y0���_�D�6�@�kB�;���]9���U���Wp^�eBO����ю��?X�)-�9{D���W�9fnZ���)�VXq�����b���ϒr�`:ԚU��:$�v����,$-��3<T��9~ش8YH01�j�9��t���"��Y�Q�p��U-�D�pT�� fz/�3��y͝��ma�Y��Yt���T�`r>��M���n���f���̭��q��ȬT;B�1�� Ui�ޓ��J\�����K!�0�]�zk��ͪ�
�7t��~����f��^��%�,�ｮ�3� Z���<��y-�"��m8��Ȧ���E�����G\�=�9Z����ش^c���:�d��M��M�Xfg*��ʫSQ�k5���������c�}��� ��nX����RY*m!���~���[����L�nks��g]�� :Ya���4ᳱB�`E���T*���"��w���eT ���g�R��G��y-20���F�r{�\.���1.�b��� ހ!����=��<���˸q�N�2yb��b�J����=G�-�����E�x���~�¹�zZ��Q�̛�WⲐÇpKD��&Lv������ܰ!�C@wt�GXO8�o�	_YZ55p�(r�+5w�Ƽ�?��<����Z�\�����L��x\�xa��;)���N�߰�n)�U�W�-&˧:b���tT����9�UDZ��eZq��g�3��p�Z���g�}�W�{��}���d;��|)O���M������o֓y̖�@*��}M*������V*�Ge�A�����U;b��
�;�����*`�q!��)TjB����+���U�»��� {%�D�x�$� ���Vʉ4�$d�Kz��LWa������A7g&2I�Tp�:��4n|9����Nܱ�.�q�'U����g�(]	X) ��c�[z�ԗ[��L���F���Iy��q��ž)"�y�d!ha}`X�ǒ8�g�@L��X- ,���B�Pj�mX��=-�*�l�[
P"�HC�3�D�U�����7�g�#��E�c�F2��2яa� "�*�J�Ɩ.��"t��*c�p?Qs$�F�W��S��y��!N�5�d|*�& i�  ��H�Kq��`��K���5Dpd۹jH�+d}��*�[bD,ܻ�WE�{�S]t���St#8��i��C� H�<�z��bZ^���e9��o)��U����FeG��;=�����~��BA��A*{�Fc�>�L������S����`�	� B��dF��o�`���S�����п�2�|��}/���Dg-nV�,��|��eP2^�`"$��j`�� <j31�:(�����L�;�p�"!�E|�}��oqo�aH=��	i�8wۭ�M���M#�
'��iةIS��g�H�����٩�Q�kY[��N:AH�M�?�N{)oL���$���l�)�P�}cgx��j�Kl�)힫cM��xv�$S8}S'��b��^1�L }�Tn}�
�nR2ݕ�?ˆY �pF
���.�I���o�k�m&�:���H�
,�Lt�P�5X|��$�/Z}�v�U��uUO�Ui:�����ᵴ��¦�3|�b�N]"+���}O�������"� ��̯K�c#ͥ�ZcSg��m���Tf5A�U�2E�A�a��텘L�1��E����dE'^&���*$�,��.c���*�$��t=Z0GĿK���7.%A�.rh��	ݢW(PX�K���*mC9�ٙ�f�p���2��G.���g���T5Df'��_:�	�c*p�m���f�"���"�������S���ܓ�v��<ŉ��w��t���(i����+t�m)0)�CG��d9B�P=U֚-jjV2z��2�'�2�J�4��֐<U��8cn�g�ǅ#�K�ס�- �JU��z�M���T@��h�e��w�W�3I=Z�X_�t������F
�����R���k�RT_r���mc|��p	O�g�w�
�!��Lm�����1�H���G(Ì���謘>�-�Sc��-�m�K�Ɇ�s_�kϛK�y��P�}bp�tSPdC@�2]�Mtb{v��8e��e?�7T>�������]:v�._5r8�WaG]�����7}"�W�Ծ��Fɵ���ˮ�g|:?���v;��6c���t��P]5��{�q1��G�q�Yf�e��o���I�w�ʹ#C�m���-9��'p�������f�eF���Op��~ ���<���A>$����4DSJD��F�DqA�<.;o'V�Ն@
:�-
dK\�oK����S��� $�Q�9@�<+}e�Aȫf��7��?�QH��r��v4r�5�@B��,tԗ�&�X������e'��O��?�aʘ�B�~uJD��rSK {���iK�����VbAm��Df��?�'T@ϿpX����uT�\��?����i�?���D�D�9"��f:ޱ-.a�`Ƥ(*{Uݘ���N�#NH?�hr�@F@�A����㜤^��|z�#쭭3`�x>�C� ϵ�݀؀Ԍ�XL��H�ۛ���7(z��n`�.�)��S�k �	���w��6�q3X�s���NIo�=S�+x:��Q��<��E�W�Ii��F��0�l5�V�M�l��"���k�7&���沙p)�Q�?`(��kH������6�|�N�9�4 e�*�$�k���'��I�9�"&_��z�����n����.��5����	�u3��N�����^F,&<�A_|~IS^��N�N�I�{"?' a�D�����U0��t��(�SnL���{>��q�-��"K۫�8�ߵ��I�)�d����N��	������h+XL��I,\�˚�b��2�����Pq�T&���z4֯�6�'�B�"UƷ�IP"ꞣw��w%�e�f�Ω�� Qo�P�nݧ�6�~:$s��B)~o�Z��]��d
+�7��O%���[-8�̧�ش�������W��"�_�C%�h�������[�ځ�:�ŉ������<9�"|gތ����攑�5Pt�E�pr�.��Q�'Hwx�&is�E�qW:b#��עXR4
��2��O�¶L�V�R�3v%G���Pw�G���&O��N>u7͎�߿?�Kak�K��ö��	�U�Zxq	���PsQ���A��ju�k��ũ���8�^�I����P`/?ʮXvJ��
�L!Hm�M<4"�uzwiB<��&�k��.��gu��1���P�Xf�Wr{zu�_D(������p���	j�䐀?�c��k¿��ҬHB��J��U_�Ƀ���+��=���nE�����w��1���cu�ܖUN}e���2���y� ��żx�\xR"�š]��۰E��\D�aE�4[H���������:�%kH�W��5�!��p�޳?u��D�r2�#q��&�]�TA���o'�Z�-m��~����0b�08ݽw�:>�4�L��� +\吐{$�ƽ�6����J���r�c݂q�n9C@~_!or�I��I����
<g�r)��#���G���з_�eF�M}qV���>��5s��bmM��%��$�' ��ܨ�Z�WvPS�<�2H�঩�Bc�W�o��zx���6�b0�_�Qo;�?��-�5#��fsP��
�cf��T�|g��3�L�J/<]�e �5�<�N������B������z�Q�&Ok�뵽����hoWt�\G�	8�2�$��9���-=���ŋ�('/U�;��Ts�(ԑ1NJ����}2�[J���({���%'1�k!Pl�����H0n��z2!�n_3+�BB��3�b�� ��]�յ��w�n��Mck��	�G��1R/�
�͐ e��a�.���H�ǚ	��نX��<]���)lL�B�(�JIњSR^-`j�lUe;��*�����pҌB�DFu�o�̪C���b���R\��&	W��`v
��d�7���*�Vc�D�O"�>���뽾���i.R��Iz������a�����A������:ߧ>n���K��x��w������f�tÆ�0�LzK3����@G��w�8���������Y���R�� ��FS�Z1jd̄�֫�a����z�&���H�j7M%"�HzB��%A�E�
>S��DOrg��Z|:8�5���d��3
;&�gD�� �R�h���W)��ӼW�[�2����z�y+c�T�|Ӓ���
��tJ(��7u�;$b�	�U�5���u��
Nl?<ϐ1��bE]��"Tc/�����J��}��Nl��VGgoF鎯�L��}���Y#>�J�)����_;��r;�'�ʄd��l�H5���7ɈJp37�ǀ�?�k�ӭ�+A�ݓ5߹G�&*Bթw�/A�9�Ȯ�����:3ce햔I�U �x(kW��#9�:L��o̲�鏋'�vU��iv�a�u�>��JCh�pD�H�*�ݝ�P�3Jr�GCJ���9ށ���xT1y�x�c�}����\)Iy�g�a�6(�nN�_i��J[g�þ}�N +jo�z���D�>�=����9!V8J3��>���Ձ0����l�=���U��r��X������$M�E+y*� �,?U�wv"��UsG����*�͉��?�zu6.C�������B�1�V���[@8���wF󐽗�K�tGtP���ƚ��1@��\��>4(�a~��Y�g��x��w�!4����6�b,j����1"pN6�������5��EQ9#.?h���	-g���'� ��^[c:�Ӎ��5>���Ϫ{��������WnJ×I<*�*��(���%v��yz@F=[�5���:��L����8+�"�&�x��~�bas�6�Sβڧ�/�1���3�{�P�� ���i9�Z��YS��d3J��&q.�~<[�wƹ�˷C �ӆô�Z(^g:RAj�g@��<M�V�*��ϯ���V޴�/�a �x�qԾ���Q��:�����&���G؂[���W�����,�?�zʴAҲU3O����Նn�d��1Kg�lэQ���X�k��)-t���eE�ܶ�u�w�nh�i��cD	߷[�|����N��~����`��|�K����l�o��F�ی�_8Z#b2<�3t���)�����Q5�R�;A한�S�X�D1�6���7�-�^�.�.���KH��B��E�>Tm}����0MR�ه��R��4
D� @�B��x��h?X�#� Y���#�]0C�m��8�AV�����[#�cAѰ��n�mB�2B}LAg���&�ߖ��D h�����I)��|V:j�����=+J)�mKM���!���)*�i����r��q��O��д��0�fS`������I{P��$쭁d?��>�%�-��G-�X��8v!S��B�fؖ�BU�m����Ba�Z2%�dh�@e�� n�N���D��$���G;0q��=���^8`�x��g�����#�К�B�J�0�Y�/V\����}��ϥx{�W�U�/aI0����fܴ�IoO�~=�D*Uv����ǒ`�㙐Lf�bi���"|K�6������Fi,��	~�����|�!�&R�p�\�a�;x�y���ϣ�%����[&�,�Gd�m+·�5T�x�!��:UJ>�� �T:�JI����'�]nAc��<E�׸��4�4�TZb�n�`���8�;�,�Bh^��zԪ�t����1+��]���;��k�E���D:��z�/���@�?3�8�����~%b;�����%B�5J�I�X}����/s��"���Z@%n)�"�+������z>��d�0��qdo�K��N���?�
�H��!�^r�n�'�I7�dd��>}�K�S�UD�9^5�3�d��Jb�����ZAM_
`4�"�<b�"������ҼHŔ��<!"��gːLoAo��j�@6��~̠di7��[L��GS'be/(��|]�w���'�!����S(������yC�V��J��~$6u��o�P��Ǒ^�32fk�n>Xn��r�iC�_���m�oo�JF`�D=Lm:��=���R� ěyQ��֭�:/о�6Ƞ{<������)�L��>�YV����K��N�r�F�oX��L7���B���"��=���.����Px�;��!��\��J- <�r/S���MZ�B܋QԘɰN�^�� m��y�Ͳ�����	�q�-C"y��R� �رG���h	"ۓ����X��Q!�F�W'�[ǨR�0��mI�n�bͫ���!�j�_�������̩��;P�let�s�1���Xji�	T6+C雟����w�-��Fm{�\ATb��N�q�GS�ϲcn�<y>Ha\ș+�Ը��W�V�I���'{�_ùCK1/{��MT����hjK���s�T�� �=Fl���f�`�,�"��
�h�N�6��J��e�9L��	��<C�7ܙ
[���/do�H�<�_2{�~dCU�ËEf\3L�~`����A(S����r�~�r@=�d��.�<��WZ��l�Mg�x����k�������qlk]#F,N�+-$�*ғ%�^	f�!>oeMw�8����޼@�ħ�z?j��>O���,���$׉�[�!��q#�n�L�1��a�^�kt�6� p�Zuvï���֩	�`��Z�h��z�ե�	(�q��Wp�M���x����Fga�X��[���b�W�3|�I}�F#�!`�Ȇ�8�.��5�E��%X������]����ei/ЅM=��g�I�$�xwn[�P+�Jk�h��p�N���SL$mr*�����X#�$
;"��V>?��u��Vl�5�$���\�FDHA�α�22��>�7(�(Q:�A��gx^m���'������!AW6�Q���8=5�]�K-��&�psR�'L�2��T���D|�B�ױlj�X�A�<��5�������sJ�dry ��޻z�ğ����g���mR���Ñ�fBT��h2�]x�F�TÔ�1��_��;�'�y���2*�	Ĥ�������:�S����.2�6<��Pm���Vr���F�A)��lF����_��mL��)=(�"��
'`�Xc<[S;�g��dyJ�m�܃ E���P��}��Ϯ�s5��@�az�i;w�+�.��G7���3p�丙�V��V���v �������:D��N�X�oi���vW�8�]Q,���w6�,;u���؄\��h@�>�������ٺA�i���p�!��F��S�eCK�oZ��[�I�>�#Й=�kL��i!�<U[1�V,�(�V��?h:$2�)CH߷�x댔��|V��늚��)��*�n�Z�A��5ӥ��: y����Q?��Wv���f�C[5A"򲫸0�#��5�F�o:��E�y>K>_M&�J5CD�&�u��H�~�{���i3N�2���C3y:�E��G+>�hB�g��(?ly�i>�9\754NN�G�^���.ol�������� ��m�a(y���d�@�@�Bˮ�-�����-r�R��R9l�?��C���n!"
��Qcx�TGٷY�?���*�T�e�0B��xш�C��a�FN�T��J��[�B��B3R�<z���Cwz�K]�La�׎?O7���؜T0��N���1������Jc���UA6��$,�xy}!�-���n<�JS�!��3g[�Q�5��8�d/DJa��|�p|V�F"�HE���)�|� 4&�Hp7��	��/�� �eh�w�3�hq!�C�=N@|�
���XU���p��H��0}��4m��,/bG�$�p�gj�a�>��<9�n�X���!5�|�?'�˟�y�EЌ�52H���b|��0!F����+��Dʝ��sR5�Y�˽5a!�)�q�?r������31Xc�uya%]Lb�������q���
�Ì_����(������"� ��*��k;\�����L��o�TE���3���� �Y%�+������p�,B����M�z��JV�Z��,�ބ�����`>~fR+M���U��)���?�n�3Ȃk�h*Ns-�k+�}�[{6�A�����7ʗے�C)80�`��"�K٣ȯ|�����CB���,��q<-�x.��eυ�u?J�(L"��8Kf��)��:7��*lMNg�l�4r�RT0�̙�����\G:�i7�!)���+)�p���8�Wb��<�.]��P{�k��9�
�U���.�߀��P�+��.y& Q��ɛ�������XM=ჾ?R�'��Xk��EeBok=[����	���cJ��:�ܰ�)�������4�iyK��=1��43�&L��s1x嚿���B��
�����7�[���T]k�x"����Gͥ�{�|��!���T� �E�\g_4Ρ�]���^�@\��mP�w���T�]���
���4ʂ�v��h�U�Fک���7C�M��� �D}�B�Y�p��1�me�@Bt64��EL�T�M���q�ǭ5�w��B�z���i@�=�����Jں�t�9�����_��"�D���>
�.�VR�wN�ƕ��/��ܬH��;��ov�s)��	�����"6�"�s��`8W��$ M�"����I�l��>�#�_1���}�����XAY�\y��y0h�׎@6��Ȭ���H����D?m_��f�N���@�2�}�ކ@xAG���.�B���V\[ڹ9H�֣�l�?�3���ʳ�Ѳ���v��4��=J�-�ozD$?+�eֽL��降��E����l�T1�GM��[s�sH�+��0��^J�k-���W���nL�A�����{��kN�~�A��\}��-B!�)t��!�)r�M���o�T���C��mV�G�g�l?u�z=��chĚ�+��$mi5�:�~�� ��* @�	P���B�Ñb0F��{Nw������C@��Fz��73o��xFn��L��_��BOY�4��?�F���h.%F4��"CI�ζn��E��k[�s�}���ol�l˓�I^�YR��#;��d�qg�@1��H��7�9�B��\��o�@G��f�������p�4G0Tpq��<1��w���	��d�g�O����� 5_ܒ�1g��$���Ƈ�_�[�����f�X:8},?���:�`녓+R���0��K�0�=ޓ����Ÿ���:������߬�`d:\H![�L8d�+�Z`��4�o͵|.�Yt0hR�lЖ�m����i?��أ���k��R�d-�����U��Q�2��vr$��܄���W+�C$sN��B���n����+�u1a/\�ܸ!���
S���!e_$V�U�� ��Τh�׫��=?�r&�j��v9��J��:7nV`�,sN0�[�u0��
s>j� ;%ګ8�H�W��t�P�
��	�ŠC*�m�*0qD=��|�^��Q����n۫"@��i�����՚?��3�!�!���Ue��n�Ƌ��(;t$Yݛ�
�:�*�I��ݫJh���HH:m�L�3T'+�BA���'s?���m΃(i+=�$u�_�X d"f�>��2`rt:�	�N*='rZM�+��4���H���� �w�1&IVWXҷ��+c�&�_f={й�x��i�E��-�_d<sv%Y�B��Q
�h"��H��M��R��t���IX���m���Ǿq���z�`�E�P����a�[B�Թ��ukK9�/a�+P��~�ġ�5�WRVv��h��f�_9�Q�0��Q�* ���r���h�Ru����c�-"	�YlQL��aa�R	�y�NX��n/�y���f�eC���u�z���`�X�/����?䑚2=�9=@aNJ�).Ii��T�1tkd����QL���&T��_"7Y9�}0�,<��wO>�,��a�^R��iGd�D��b�cqe}��"��g��,�gv��(7��	3���-��6���]5ClB^&^��ZiD:���m˭ȚY��x�A���Ɩ���j�����l.B�:!>9A��s��z���JqJ�����\39ޡ�0m�ݳAp��~@>x������E"�/\�%����u�7(�^}�ER.��-���/z0h�@������X
��Sw�"e��[ ?vA��n�f�u3��U�}pZ�e�K����gAɨ��>T�#Oi��j�h��b}�L,P�@�'���c(��͖d���]t�sh�a8]j.?���j�q�k��F��w|�9�N#Hh"�yd���T�;��%#:{�f�j��'���i�=�z�*�ǫ�v�{�(/ݡr#n��fT���`��s�����_�K�QVSAG�|��~���X������)i\�T��Ί_]r'��d�&,�B2�i}���@�CýIkx�'����xj%�Ƭ`�`qO�A��7���i�u��U;��=Xʛ2jHe7�}�{X�wLe'�9�m^q��X����0��.v��)д��D�1�qj6�i��R�$E��O,y)s�'G��L�c���� ��������t��f�zRP��s���n��45Bb�U$p�P��_-�GP�|��Svt�5�%_. ���Q7�>�4(%�^A��6��x�U��d�����(��3�M���0$�N�8 씻)!�Q��?6�t����`�� �n��]S��t�Ø2z�-����잍��2 ��� nl0N�%Z�㮢�ZL�_y�*���d������o:� �M�)�\��9c�v3�J�����%WS��;Cev"��In�01΍�hA��	���k��ޝsX���$��t���U4�?3�Y:��7s�ر� k����Ҥ*��ځ�X;#�,_B�"��~�g'�6r���������g/z�����ӯ2�L�z`9� ��.߆�@Nm��B��%pOϞ5y���;�v�<�%���%����G��L+_8:�Oƚ���(S�r��*�.΂$Qϫ�͒4�����&KV{HS[��n`^�lnS��zx�O�<!����e{�4�����TBy������2j9��1mjMn��gP�gC�AZbo���y2�>���9��È�5��E+�h�&�(��ü�A���]ī����כ�5 ������z������*
a�h���'�O�_�8!z�Y�B�ͽj��L������2�t���+h�����ڕ��5Eѽ�X�����Q�Q�����_�l����� ���;4���]j2(�W��o���J�-���G�ʃ_�^c%��.�t�8�s�W����q�kѱl����|�hG-�(;y�S�	�pO�Dx�R,H�ė���x�_U���kW���'�x�sh�>G!;�0."+O�@-��v��)�m˪פ3Ϟ^�EΈI�XK��+�����������V}l>/�r�x���|�G���V��Gʐ�\���I�������!6 4��Kd�hh5��"�Cګ ��QJH�<���#;y�^)�MuI^f �۰�5W@�?rTu"�׉�M�?�<�Q&l����ǝ�[�-
a��� ��@��	��~F�`���}mzS~�"�
���?7lQ�?�mJZO*Q)Ceħ���Bh	����G�!�)��r6$�>�F)ې�7!�AQ�6u��H����E��2���U��=~S{B5��K~��9l�&���6:���+l:AI�UW�����G*�e��bnW��t��OƑm)�\�^�f'�P�В=1��!�d�L�H�וH/m@�5�3K� 鑟8�7A�ȳ����F��f��	q��ɞ�iH'M5l����(<CB���^(���D�����>;�DZcڢ�M��Y�^갟ݏ	��0��K��q�Ɏ�A�����UK��S��^ST����K���P�ƵGmk��"�z�8��m��EQA�\t �Zߐ������1z;7�3P���	� ����j��*��V�k�9�	yoz��E�]_��M!P,I��`��5p�3n�A�����V�s�c
���fV��$���( �j˘��?���ȝ��n^PSA���c��⧜`B�a�$��*�����4��j���u6QSu	P�g��X�V��� ��b��&�֕�:�~��Ng�ԝ����#o֭���z6����)2���3|�U��b���LY����3�I$E�ܟ�a?Jض8zH��w��{8���e_�F�z�-�K���h�j�f;�R�N���Qyc0�2���Tܫ�"���>����f�����Ɨ$������`�a�4ë�"���ޡ�CY�R���>�vWE?�!��Fkv�F�YD=�ŭ�1̆�h�����#b(�@��ٌ(w��C^0��kT��p�c�yʷ�'-:��'�i�('�;��	�Pb����\�<"�f��47�>X[R���R*x�`3f�Hb��4x�S��;�>k�Q�b���g�AA�0��V+mI�!j��o;>��>�j�f�~�.�c��㊳�7�yWL���F��775y���b�'��slÐN�b0�6
Ė5H�ȘA>$7!^��|���ҝ�R*rVX�*Ѯ�x��ܠ�,���G9��.m��B�����%�9bW���ܵ�:7&K3irJL��Hw�`?�;᧻��_��S�[�2`�F��B[W� �|������m|^Ʊ�a�"RH�6�U-R#OJ��w�={(�X�ٚ�B5r)�h��P�[9���[�7�K;��
0+ٿ/����LK�FY�m�δt3J�����/j�����ͨc��,�P�{��Ϊ2�=��yo9|� ��`��5t���/X��5���8W
����c�ٸ}���#>Ɖ+#$���gj��E��T������ig^H�X�q0����{�_����{u�<Ω������0B%ڇ,;��'���jB���縈.@NК#R���dI�����34#��4�>�u3xr�h)�v�k�R�>&�q뺾#,Ϯ���8����T�c���<�-S��N��톨���M��ʃp�F�b����`����+J�,i��n�Bg��D�'�~r�^=ۮ�=�'�a�=������#Xo*Plm��/��
��v���
L֡9WM/����|���(�&h�V������ϓn�+�
��b�9b��oa��L? <G" y�0�l�6C�{�&�"L���u+)2�����h����r�k��ٷԎQ�c�R�5N��7����Ö���\b:&V�U��r���{Dpś��S(VψՎ�|�6�(�/J��3��n����pF3��� Oυ�%xr��b%.������/tJ�� 5�9�
:Ͻ=���(�9�|}�����|P�i���I�J~�h�Nȷ�@�Agq��SC�:(=��{Zp3�mЄ�?'/8(����b��5 ]q��(�]�2:�o�n�ي���Fqk~rq�5�̛�iăfYU� �9�����f!��Ե��>|����/v��<{��y{�p��b͊��!���<e,�t����xԯi�o���7����ګ�eW���/ܵ�DX����'.m-������7���aor�������Bs�$��T�vd�{�.p3�,sFÏ�n� St�����ߙ�"��2-`bcM܁���G* �K=��	�>t�NJ7��p���nP��I�~�؃���Qƈ��%��hQ�ݟ�#8Y�K\��N�-����Phk9nl�����|�3^zﱕ������C\�$І���БΓs��iY+����ޔ�0�n`)Ɵr�J����"��bIT
؆��@��J=<+UϖTz��R=��a�8��n��I��q��KU
�����̹���6e�*���C(آ���,�I:�	����� %̅t6�e��*;Kg���f��FE�[a"�"�y��|.ջ,�JZ၉ac`Z�'�0�0xc[Y��{g����h.l%4
��ܿ�4SL5���kMNM�Z��r���0��n��P]F�
��×���1�p����Bk�GM�n=#�MW��=��k�P_`�N�~�~h��!����~ڥ��Ds��\	�P��p�>_��'k�)M��X��GI���WL����Z"�m�d)/��d��쉩JY'���%�׷,�E �������g�8%�>�0|��n��D�.�+���j?*��hDK������"�� <�Ŏk����-7�����$��{�%4�ݘ���e�����H���O��"�<g���A�C��K�IS�V��tӠVC�[L/e�hO��+GK���:(/]\ʓ��5����!�n+�c{{B�o%�}����'���Dr��\�UO��(��*2��_�ʻ��8I���{���;�4��m���)5f�����I���IK"[Y�Zvwz���s��.ʛ��a�wI5[�Sa��Tl��V4�v����{�?���%����
�5�Ų��@�_�Q�:��e��`�mT���h��1|��Yt�L?��"<��7��l��)o���D3Õ�Co��̙�r� !���!|A"��ß�=̏�T��l����y�*Rb��J��-�K�LS�*8b-ľ���>=�d?��b�Z��H�����V��6���.�Iy�\y�G�<eN�"�x,f����/5Sa�2��ބ�P�u�Q6�eo� �_:��=��/����95��/�o��6=K�S#Z>(��ۧ��lM�V�$���U�M9Z�����^R+���Ƽ>K;��b�\�"p�$L�DSxȡGYM�gk�2�d��������Q��\��AvE���A�h��Y�ck˺�g������υ�%i���]�6��t�Jq����.|Ɓ�����@0��hP�V0;%�ٟa�q���u]���B�����l���/�y�V#�8D"�7������{A�iA�s����w�N	��� Q�����,��T�,G�������m	Q
���v�K����F�8��hk�	��t�r�1�F"� �w{�~����Ml����s��3ˡȄG���&�rgD	^K��P�Y��k��<�u�"�F�4����YtK����U�+ܳ�S���Le^��П�ۮr��ƕ��Ð6����y�bEB��B�h�`�A�!�˞�B������|,F���	�`��UP+c��,�m'�c,���'R����I~��--�����`�u*M�Us�X�wLGu��A�v��\
s�m>0'����])�މ*O�j|S���nB�4NC��!Û�ֻ:Xv��9~y�.cuwe�<u;��^���1�ki��aD4�j����/��v����O8�U�r2��������t������崩��j@��X�X:�Ք�;�Ÿ.�M	�^�[J���2#ȅHs�P�l�y>E�ʉ|$��[IzF�'M"��sv]˴��*й)tN?/�[F����/��rn�|�3�����K��N��"N�i���o�`�~�Ŝ+�90�:t��_�3�7�Kіrt�P����`gO�Ȯ�p;O���2�t�6�/�.�K���g%�f���e�y��v��φ$�化r6`�ꘔ[M"M����+�FcW"��q���y�ɑ�����s���P�(�����|��XvCh�%H����&L�i`2"I��Þ]Y"5�-����
w���O15���']v��^�������<�O�³�Ɣ���>��N�/��J�������]���;�
v��f�Gɖ_^61�uK3���u��(��Ҵ�p7�&~����܊r�f���˶�}H'��*���rZn��k�ZlD<5׌��s�%k��l�}_�-	mu�
&ن���<.��Ft]��$=c���6�o.a6�����T��"?nf�%JY{�~�2�)�呭�D9S|��+ڸd��n�NgҺB�>�F���YE����~��8g��:�~�z��}�i�p�a=�I�β$�[�q�2՜fe���g �e��o�ۺ|��<��%"H�F�p�������ЙV���:� �-��n��N*+8_�N��ko�>{<�;���5����B6	����B��
�鷲o�B�p1��nǻt�.�������[Ɯ�cRZ�����

�k�k�Qοb�!�O��w}FQ�����^Z9I�J�e�`�y*��6fcC���t)!7+�/7DX�Ĭ�7\�7�DjtbR[ȶY;�up��d����*�Ͻ��N\���/��v �'���nK�K���L?�;�~E�����Xa�]�{һֺ|��Y=�`]v�Uu�+F�������Z"p�d�:0]��-S��g&)�Qz1��r�}6�)H�i���|Ӟ��W��MXT�}�0�^�}���Z wP�/YN$ɋ����V8�]l�\ʧ�� ��ݖ�����֛�)�Z�O?{�ꋜE��A<)R�KzGk�JKg����'y���~�g��n(�ۢc"��SN@Y�:i>zƝ&c��﬐_��(�� �%��^�z[$B��o@_d>�(�+�х���r[�A}2C1c���qQmZ�dZ��VH(��hb�œ4-�� f4�������3F�(��?]yO��x4h~p��)���)��[$'�1S�<N�'�lP%p #��$N|<C=B�)���u@�]��
�m�VU'�T��� K>�m�E����}İ�鋥��xCkE����y,.�Dc�i���˸�0�M�����W��D(H_����Bsc/�К6�l���{�m��
��>L�Q�Y,w�Aɮc���v��ͮ��/v����j<��ik�.a\����Y�����5��p�~:���H=d����Vy���'F���� ��Nʧ�3��q̤����uھ�Zͦ��T��{>;�)�i�%�������?>'~����s�C�c �{WB��,�%��!N��xn�i�D8��v�\ޡ�u���V��i�8j����F~��i��%3�x*z�I+J�KV������_�� H�[��Y�)�.6M�c e����;��|f��c2��->'�"��enө��6�\�cw��{���8��J���O2J�X?*K���V1��rc��.��l9�ɣ!�;��B�T���[�1Y�UQ|J1�*��l.�+�!���K���F]9\�T�=}�S���R�f�D�N�=�/ C�Z<��s9�,e I�	�}� ��NR��3����KUap����R:���b��<Q��u:�`�\�a�6��x��,g6V;7R$��2�/�U���$)�J�֮Y/��2�d��ߙ�.�.���)#<Ƚ�������DU�D!�Jt ��iӠc?V����R;�ط�U�������,=��J����s���[7x$��V�FϽ���:0��2>��"ۗvp��#��*qvj��K�<<��Ҥ���<���p<��z[ʩ}�P��K��v�My�#Z�D>��@�C�sk��c+\�x��iX(�:Zb:�d�h���n��O���Ǭ��.�-�;F$�y��
_�Mo���t�����Sbp*x?��~��F3���^-�6��t�0_�ԃ=�!�����e߉o�r���-z6�L6��a�B��^0AV��f�����C��IzZ���O�ֻ�1�Ϛ⊱
�F�?�����kk�j�ӣ㳌�;����7r�5벿����Ç�y5�qE�*N��Ҍ~����%6��U~��҄��VIM�jW����%�^�����Ё7��u��\�y��"���=FY�A��G'����U��9��S�����(۴y2��pˡ��}p�zନ{��NA��	4񞌛���d����a�[�ʃ��5P4��K\��|[1K����Mկ�C���jX��P�C#�"4moW�w�*2����� |�<�K�U��`Z~��2^`�{�x[s	��9�8LǕ�ڡ��ϝ�7��	�&#��$ j.�AY�{ȵ���ܱ�x���-�@@u�?���UMؑl�gg䴤ƌ��1����)�=痄@+p_� VM-�Ji.�ІW����O�%�(ϴ��A��K
���Hir�`m� N��y.�\�y�K��l��G.��ZŁ~T�e�R�-M��v�bXZ���}T���>�
#A#��ۼ�G3`^�!��߁Rd��ݙY�'`O�(����t�E���i>Eʁ����ݞcf���5@���
}�D}E�.��h��G�z:]ݲ��7%&ЅA�p��\�1��"BS�i��E��J�k��e���n��g�wfN^ҮB�s�9�� N��iBU�(����#�8��L��z���/tp�'�/�싖����v@hI���d�i����s9}���E`	���Y�uHh�y`�Oé,�@N���N�R�_��=W*���?�C����h��&b��ͭ�43����i:(/I����Z�~J��`��Y�ˀ�蹂Ê����Ew�<N`,�՚�n(���p��;��C�_o�*Y4x#gS���G�񥦷�Z��zei��g}M�b�����%��(7k��t�HR�3�3s�Qcz�Ԑ/��ٓBo�����*& 7�į�Z�p�ư�lX�aoP� ~@N��ɩ��V=�fo�+|��R�b����[���޼lJ��#��� �7^S��>�G�m�31�$���hKV&�o ��@"Lk��#�̩�Ff]2$A���/n��K"C	sd� �����;��M�Āi�)��fUtW�@Uz���X��c�C�cxv��o�A`oV��kk���S�8��Ā{Nl�ѭ�g<�'u5?�H$���6>�MWjVNv|�Sx�,W* �r��>ˀ�ʎ^�e���VY�9��+6U�A�.Nܣ��ML�Ͼ��>����啎���/�!͕�ë�v���3f^6��'�3O��m��T�Ah1u\]�p\vk��GD����������C��TP,}a"�%��� )� ��\����q���g������� wmQ�2�zlgh���Q�>X�@��퀷~���x�����c1�������ӆ��&3�	�ݹ��*ټ4�.qXQc�Y��i���ډ�P���*�1���:�h��{�ƃ���}�r5���#���ˁ���,�D��Y�H�(��,E���;���J�F�u3�ܴ�%Ң ���{���=UE.�Sՠ�Ai8�x� �U�b��k���:�lq��Q�a�K�z@�{�TXƘ�F�I�I��m)�MWD+���'	+8
=dM���f\[�pVX1�(�gkCUbgX��#`�����>-0�\)��ə���]P�-12}��`��$����꣠���.�"J��QS(��f"�c��u췣m�%�N
��H&5���㾌�NAk]?��v.������,�6�(K��I�KL�D!��q�iG��gj�Rf��>p���=ъ�5l�9�ƫ�X��8�s �~��S���-ZݗK�E���C�I@e:��r��t��	�-�O[����������:M6�� ��TD3 l_JOD�h>��]�hN��[�?���泿	К�l�q*��\���ˣ���@I b�1cg�9� (/L���A��)�
��=]^(�}'�u񶑅œp���OB�S.r<����%߇2	�'�'�"����n&�

�p�j���U`��WL	꼧���L���|(Kb�]���f$ �����9�1Vk�=���L�QV��H�<i3����3�3���
�_Q��6_�X�Ȧ>���,�v�(2qN����� ���ٹ8�N��~GǍk3��l��x��qk�|�H�M�d��ic�pr���y�¸�)�C��j�	��WzTr�� �U�Y��r�L��x�3�J�!��{�bg�x�Aye �_��5E��9/��Q`�r��U^M#��X�x{·�V�J��W �C�S}T��M��F�<�h�9������9���WP{��c���yWc���M�s��hR��-Fw���N�� �7Rqk̯��_�^z��a�[Ѓec��^rXu@�Ϙ���bE����Hσ娠���2q���CЋ��x��lY��$��l��<+�Jc�B�A`��%��.�/�/L�| ضp'_Ê�==��9U$q������֦�Ѫ17o`���"�K�԰����^�hj����o^K�G ����0	s'&�=��"�֍cG\��;��!��	jd��SlS�㋉�2IUE<P�
C�_�T<*�D��}�A�k��si�Ѣ�в$�1�Fo���!�ʪRr��B^�ьA�̊Pd��� ���ڳ�����9Q%i�+����Q�5uq�����Ou���qԒֹ�����m�͛�C�����yf�^�I��Ol^�a�v��$J�*��n̩5Ei������Ey���(x�Jv��3EP�R���f޼3=vQ�`X�Q۱�����y�|�HF��1�S_��|&��B�4V��Ӧn	�2Y�@��A
?r�	�+�����Hf����n���!h�d!�-h5�:�O�2$ T�7��Jp��E� S	q��f9%M�q�p�4ʃbMV6 �Z7���փ���o��r��ױZKCjg�9���ÃVq�׮�c2m�ty½��$��${՗g�����^�iB�$vΠ�왌�sw��w*���*��)^ݳ3���>g�c">�t!��pY*��ww��0�Ǉ"]��h7`���+E��&�2Ӣ�9o1�9�}��՟��>�=7qE�2�ϠPYCR�;��?�l@�3.w��g�B�"�5�/��>�B��=~��ݓ��bǭ�"j�`U��z3��]$N)fW�b��y�J�i��i��q�B,[� ��ߪ�L^����$+q�R��eګ�R���d��S �Q�{�2�W�j;�����v��b��A�<��d�m�LSLn�8T}�md��D�$��Cd���c/w�p��?���(���PH�!4���=��S�u�ݥ>�-I��XʨZ JWێ�	��B5����i�S�%0���،z���Bz"iǀ����0��I��:�W΃��!�Sf�G����+�^�򖻴Պ�f��6{���2yn�A���GӜ����i�6g�\b�w�.3J��Ȓ�(#0��o�L��)� �	�����釟va�9����C� �uv��Z�X41zZg_�>]ܪ]u��":�t�� ����,H���F���)��O��h�O���'
��| {���3mH��qm�ex�o����P4�0(D���;����7��$8>�_�5�����+s�/���w�Y�a�xaK��|�T^���0u����3/ *�l��廵٥�Ν�\����d��@�p�7dPԹ��Qm��.H"�����d�p�*��w�A��F�����{k�����&'�$r �0fQG�i
N��]�B��ǣ�������K�	�ʵH��0�l'fη������e�E�e�5�Z/U�"�v�mY]��N��,5\�+*qd�p'��2�J?�M�_�!z��Z}c}���U��4h���Y��߱y
�~@�JܞZn0���/UMs���/˛y�z�c��+5!t�@��V�կv�8,����U�#:�>q�¹�"�}�Dw`� /"�MN�s���~7��v2J��)��`����&%��^±��{��ؓ���q���kk�^vB� jϭs�Z��е^Rq%�2� �J$��P6��t�|���:.����?/;���|�ӝ�y�C�p��ڤ�s�p�*�����eK�&'59EgӬr���
@�b����m��4%_t5.4�A�6��γ�`�s�K�Fo۠��$�#D+�-�� �l��=؝#h���B�L�"�����o���y�O��;W=z%RfC�qv��\ *p*^�Q�j6��1QnMhR�/C|׼@[����U����?�I�ŝ�I'$�۶��z��@ܱ�GT#��hˁ����ω\KC�
�7u
%�WBLf��+�9�v�}��=s�Ř��*��w�y�@쫍Ć��%��cU�6|K���k(��n�(����{���1QT������М��C����kvUJ�����g�774]�����#�r��y�44)f�NU�ME���ܲxS3���&��-�[m��w�No@s�H��uۑ>��-�UN�{ Ԋ{;�� ��3��;���&M	�Ltl,�����w���U��|��t+���3ڃW�9<��_�u�e�E+Gۧ����d$����Lr76�������M��H���.Hj������0����u3�]����W�2�OXTp�C��IQ���k}F���D����jX��<�H��z"�8�,�Z�6�H��z;�\g;y2������͵`�g�W�Q�\5�!Ejel0�`��)2.(Z�$@�~��>�jg@����<�MJU�F
�a~�K�8`��r'��R�L/�zc����Z�t6�<Ǻ4ؾ%�$̱p���%����eW���M��aj�VV`��Rٌ�\6�2�Į&���.��n�z���+�TT����e�B$��|���"#n�39�`������]��D�M^����Xta���10�' ��V��A�t`CO[���j���ҍKl�0�5Ҫxk	 ʸ�|��&0�l(��d�SV������NH	�s���|>yӯ3���]|�Ps�ݨ:@�Ū�창j�|>ǅ�0�j�}r;�B H��F���Y� �$��uںp�x}?� ^��c��8�y��4TH��k�H�]�g��#T�	)�}��|��Z�t��v��_��Sp����N.����a�/ Sr���SN����e7��I���/�f��uE��U&����I���m��M�?��J�`/hݡ�Q��j=���- ��UӋ��QUK�%{���4����l�qc�A�B♙�D�+�ǓdO���BX{b4��Ы::.�ͻ�,��q��):H���F���
Q��o�)������(uQB��X�0��a?)f�[�v�	S�u��:��n��T7��
hM1'F  �*����� �*`>~$C����DM �90���E�:�3��k��E�X�:n4HC�8�~X�~�:e`3+��03(��&K�\9����?�������s+��^I�h�~]�ddAq�Y��/�d|���|v!D^/;A*8t�1�>΅*�c]5c���(�2��-�ʵ��˺0�)���2P��NU�j��>L0v��F�#��S�8�8��EO�w'��^�KX?��6Ȭm�$t�%�o}V!vbj�ɺcI�bc9��ptۉ\	��"Wb��"9���#q7�;$��[�\�7"0���*�IoZ������9�I������2^��.��3��dh���v}��ʰ�%�n�|�Bv2��������gT�.��t�79Z2� �����N�:�}oz5�Ԇ�!�"�n����=��X�7����%���ϐ�E.�yJZ-X[C(w�4��x�k[�N�;P��u\M"�i ~kZ��}K�'|�u!6JL
���]�t_NO����	zn�ѹ�z�n�"U���BR5el�a�"7�<��ࠀ�C�g^���Q�Iګ����h�=��{�9��W��L��L�i/-�g5B�K������;{Ӊ�/
��Ԧ	��$qe�ƃMq5Q�ϡe���M���;ѻ-P�)��j��?���l:����D�BW�L�<a���p�/��J��J3���;$��F�F�UfQ͎4?�����N�L��@�� �H���@�\��	��Ƿb���_����׳R"��B�\+�_���n0��s!�
}ux��A�K��V��N�~�ppG0^�/����Y� /H#�Q	��u���kwy���3����10h�$�I<#����A��,:bm��*�.~��X�A��F�F�AӐyjjgF�c����}�+������A�z��5ե��l�`�»I9��:]#@7nN~7QĔx�ۊ��+�x��^2�Otė��9�"E����5Z?��zI$h����"�6�ȍB)��w�l�c�L3v��`�>ħ�[��8���e��GU1/�N%&h�bZo��:wÇI,>$[ljk����Q�
����P����{�2=ݕ�3�M��{8L�y�Qq��R���թ�C�w�V��F@H%�.������;�t@����(+�Ҵ1s����Ezϒ�p"�E+�z:O?O�4�G�όi\�.V�q�rMp�dd�("|�C9t����@�|���J�cK�:�U�3�o��~������j�i��piVIr��s&M)�D�v�́�tEWvT��L��J�j~~ū|��Z0�������(B�ވ�;$�@N�э9b�R�I"W�%)T�K�*)��@d+ ��F�����,�~����d�m��4+־�@r+�`i��.	��e���tÇi� �6T��a�G�;d���r�T�\�+2W��/`/* ���UT�����ګm�V��&���RP�)S�0��ٞ+��ˑOʷ�)���W��n��_y�n��Q�R�ul�lF����e�(f�sZ���8e���R�v�+����.���@{�qG
�5�U��.׮}��� Cx���(V�:�u�`>��<���R�9���BvA,��(DA��Q�hP�s;�?7)�V��Ck@�H��`��O���M݅¥���m Xl��TNJ�Hn+�xG);���R�u��(���Ye9��wv�b�k�}
}�$������n�:R���]E��m����l��q�blU7�3b�ؖ��+��zT��3�ĝ�;�2Q*����qDUp�'UإKj�6X�����Ś-mT�9�$�E@�z���a�ôp�𞟆[�q����ß%���7\�(�i>�T^]��h<�x��}���,p��Y�����|���v�)��&�w����z��8ˋ��-�Jw�6P�"� ,	����xɦ�ҵp�y�("�$%y#9Qy��J����{��nf�����m�k��s�F�Q�ݘ�<W��}:3�=�0���\�51V��<(X�/�dy~5�vJw��`ښTe�s�NJ��
�1qg�+�TՋ�F#=^(�u�U~����\C���j#�@<̧✇J	h���O�����᧜V
qM��}t4��L[p�':gܨ�nb��E�A�D�9�B+��4r��`�o��ۨGi\߆�ּ�;�F�f��Oƙ�B���-��?+Bǫ�h����
�NZE�X���.f9�Z{��1Y��vq�F�\l}f�W�'js��7�[^+���:�>���N�'��<�#��T���6V^�$_��@J�<���D/�UD�ݪt����`�!�t�+�y+*���fA���N���¼yXI��l��o,@b�9+1�W�hp�rS9��:#����W�Kb��I����|+5�w:�x
j�w)������:�񛵐�p@q*�(���Q&Ft��g�OTi�D���`V�rÚo��y�/X�z��y�����2g�%���r-�_π��L�[���W��'4|o!������F��Y�O��������~ tiH6#2�a� $�Is$�\@�~���5!��&#G�%�:5ޟ��݄�&>Č���3���N���e'�_p0127Y���7���gܧTn�B��YN�������2r����G�����5 �e�(�[�˧�v�Es��p�����)4�`��*�?)�ը��(r�<V�KV�XL/(���_��:�s�uzy�����a�O���_.�\� t�yB�:.\Ar[A˜���S��p�)*�ZTLtZ;p�O7j;p�Qɠf��~/g�(��)�6^�x 9���^�!R���V�<��H�N��K����t�����q�<_ULtP��;v�=H����d���涚K�a7^��ћ�M>]�/?�̗M���hȭ�m�9b��l	ycv7����WL��c�p��T8?3B�9�^�I��nɯp^�d!F�<��!|ȡD�c�`���7�W�A����ɚMZ�3W��j2/�+ڢ�^��Km[��^va{�??O�:�~��v
Z��8�j�	��|�F�P�cfmbz0��`��N�o���5�V=D{8��0;��L���6؍��3�N}�8��_�)o���1�1y�hfs�>v���X�,�^:���<FD/Y�.}BW�1�ab����x�8*O)Zl*�X{nW�W8���#�9�����|�1����Z������Ww�ɷtA,�6��-߂ݓ[6%A�oɜ}�D��U�Љ���>������q�ټ���R�A4�%�ƘY�|EQ;����]!TE�m�q�f�ˇ���6�($uVEel��F�1M)e=����{�>PbvMo(-F��� 4T[;��u��1�ݳᒖ�c���ƙbDx�:�5��j's(���_#m���k�{�M��sd2XO��y��R0��4aH���{x)�U�&o,W���}d�����Y;r�+ҩ�~`g��O�ȼ�t�W��
�E�ƹ:^��+���=�G���k�Vj�E��M:�*F�P�\T��	�Vs�~�6H7/a���9n�#��(/�諌n�&��hr�c:?���z����m���o�n�,4��h��Ƞ���XDd��.�vPS�M$K_8� �6D�fq9x_��q���4?�h�MME֍���{���Ǩw�n[(p�`η:_+�|��9bp.\)��7 4Z���9x�|��d��)͠u�;����Q�?aG1�zr�ʷ61,[�'[���*Ҋ�tBo���	]�w_q�~>���#7�EȔɷ�O��$i+*�J�Csm@��f �S���,1.��~�q�|Mb$6`�%��͵��,�9_2>`�eܵf���@:�i� 9X7�IV��O/��7���33T�~T�')�p5��Dt`-����4�6h?S�܍*C@��=l����R��=�o�&�2��&#WI�W�A�����(è{=�-
�W�K�u/�@J�39�Z8p%�-R�Ç�:��c�.C6�Y$J�'��'CZo����W~@��a����7��>U��\�EPo�dp+�E�.�O%���c[�|���;}�\������9.�LFȗ�_���da�.�`�3�eAmI,�I@:u*%��b/�dkE;1�ݬ��UG�e� �����捀��.{�[=���h˽��_BK���o肋"X3�ߥ�����I+��\�qm� `�܊=5�c��%���������E�G���v��7�1U�b��p����2�m:�+���4Z m�7ċ�-��ٙ	���"�C/hs�� �_�hz���&�!pIhǦEWR/ɼ�e��l�ڭ{銒2x�>�����������۱-��2� �`��	;���D|% ͉z��t(78��uEYs`[Y��]�J��d�/n�>��Xa�?x6"Q�,�6;8q�3��\��Ը�60�9#<Z�}Oy25􎷊�95� y��8q��RQ�f���c�0g{�H/�ݎG�5���/�/���MC8�b�9��9>#�h��bV��5ImH�v�>�$��mnӼ�&�(<k�f �t	�eqBp :���a�~ ���)x�Y?�'��rզv��%�����?m�?`f����o�b��b#�K�CF�0N���Bۘ�\���D1�h'��yqH��XlO���kq�K����7�ԑ6��W��<9i��8k�WN�m��al����J��T瓓��zx��>�,>�ZXx�Y�wܽ��T`�ٗFD����v�z�%q�X�]/�s�h��~H���?�Q��"�n���nUyn��:fc�4H��5DB��r^TZ�ә>A�3��ڜ�R��L�����S��+z+�2�ё�J=r�Kc�K*P��B �,�+3 q�rX� ޜ�X�����k6�'՜������j������g��M6�~<Q��x��F���f��z;��(Q����j�'V���	N�tj�K{>v^���̯�ȵ����o�2�Z֜$k���Xe�����[T���K��*����>���=��<��׹�Y�Q�qC?�_�bТ���fkW_%�}x�����j���t�$��Q�� ^��]��0$�)�_$�ԩ��_��1e�Gj�O�D�HQ��f{tY��%r�`h�1/1ت�,�#�����U`����|2ܸ�%'Y���D`|���2Af3�#�7n�1��(��x2Qw�2w&n�a��;S���h\�*�9/D{��u���f����	�B��Jwq=�
����^t',s���|�NF�O;�-���+����s�N\c ���qė��0		�:� ���`S��>k:Ņ,�O���+vÄ8J�@�O#X��` 劁#�W�n�$^M������z3�
�	�(Է%v�7�*2���Ya���xˑڥ��Xĩ�H�bD	c�1���Ǩ�΋K����*�J��b��?�J	\�vAm�g�KG(w�:�f닧h����3k?4�r�d���_�"n�~ ��BF�/���0�5�p��o����Y��nU�$bR�Ul @���=�X�F��E�������cox��p&��o��p���F�=Sʁ͟�.Z��i~���(���\xk-LQ|Zʟ����W�,�B^�(R��Xcd	s��mS�m&i��
+��H ���L�R�{1s��<�|T3Y�ݥ��t�!a�|�]��D�.ʗAS?��}\�:[6�ڃx0S2V�Ɯ��|&��6
�R� �x}}�'Ѡ�7�T�|֊9��OVW%��n$�M�Ԟq�� �U��b�/:�H
��+���h��������ӣ=�[y�R�N�5�Ȗ�%#������'P~r6v�E�$�T>/{�����˜b�,�h؞���R�ҭQ \{�7�p�AwF��gZ��?��ם���bU�?u�X0���9�	5���h+�%~�P��$���uo ���:����ϑ^�iF:J��TY2�{�×���|*��*��,n^f���k+X�,�1�7q?�I3�����'���� S�ń��|���B��-���d�T�̧A�.}��o<^r��,��.v�-p�Q�n���nR5����
R#�9����3��K�o�o������5���e��r j�`���v���ͷ�O2�z(�up��#�&�!sÌN�`���l8Y@ ��AW�;��u�����Wxm::�~���|�&{�4x��$���W�m����5 �$xe�Ncǒ���=�R�Nv�3��K���~���>f�/�r���{)����3�E����w��Y��U	s{������s5�PF�� �D�
��?,6�݊8���"9D�����w0�[#aEȥ꽚�үf	���¾չ-��r������TRYE0������,8u]k���
�Ŝ�1s��x�ퟂ=�-%��#c	�vù��F'����-L���{0������8�ܔŜ	Y�7Lc �O_y#W��6�e��#"�k��r���eC��I[*������;���h'9��_^��t%]�ל���d�YQYR�ț��\83�9��,���B��l_i?�;5����PW��y����*�E���oq�q���_��aE�P�T`��ݐ�>Cjc����������h�4��!�"�]�����٠�0�╝ߣ^�k'�(1p~|����}
�\�_'Թb4/���B��>�5ڗ�/��KXd�8L��	JaC�P���-����k�j���AF��/6`�6�.��xVh�o� �������w�h(������x�PI�#Vfnn�m��4'��,� �����R��"l��A�;�$�<�~���6z%)sÊ��p������Jm���aqt-	�s�2'wTQU�-̪[�φᗏ���o�WO�4���~�6��\