��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���1���"ء�����$�iZ���@a\wT��?�ُ.�B�-����8�î���u~��Lb"���y+����(��4-�Z]�ݭO�^���$�{\s�!�W\���]4�
�>	��#/Q&��'lM)�|2э�=�6w15�)�נ ����X����
�X��$͸w|lT܀g������MD@�*[gn��"|�Ϫ��_a�޾+QAu�6�M ~��Ĉ�&��N@!���^���vL%ql���*����S��	�΀.��
��e���/eG4�V܎ն����$��u�M�r:�	$	���GQ̣�qz��m�5S{�p&���u�)�չ:�_,���mU����3V}?��K	U��+U��6��,��94�!r�f�zw������������#*���� ����O�w'f�E�[�ysos4|>��߄9� Y0#!.����=4�<����-�m����y�VS�f��pԁˉ��:��:��@�'�mU��Y�5���k#���c�R�UE�*j�lf<��6��XZ��^c�~v�l�~�d�n�g���{ ��Ĭ��v!��һ*p��n\�TB���}J��A��������1��	�m�/lP��n���_�r�N%~�����
�Y�����{W�B�^Ԓ�z�X����>�/༫��n�J��i� oe�����,K`]�ua@�.o����oއAkP���p�3��r"0B�W�q�ۃT8&E���A:�s����LN���l���)����mzB)��_]��p��{zru�@��{k6��o*y��t+��w����]�"|r]�3���������2���CAtX��bd�0��o�R4?MF2�}9.K�2�hn%�M�@y�SJ��@�QG��l��+c�3a�Z�cMH�(y:�6Ob�u�1O(݃�����j8��?|��t4���N}�D'�B��}�ՎRyB�/��j�T�r��,�߀�%Zy��3���g�)cͮ��)Ӧ��m��4߯Ї���X�s��+|��a��ژyAE��FG=�{�X�NC�Y�d�����N��e^k�N+��9�~�c�q�C��ɾ�doi�[,j�>j�	�V�L�{�@=�5�=9��HTI�^Ԉ;�X��L,�z���m�b�B��e$aU~�]$� �ZGUՑ}��]v�#ES�4.$��"�0Eeg����`lH������z�{ ����ܻ�u�ݝ]�t�s��$y�&��1sX��JlF�W�Q�\
w
��LG��#�ߍL\�U��<L�����⫀�T�I��M@HVa�(ɿou?��[�?\!���h��B\�"��=7��3��^D!7a���^l����.�R[��]�
��v�F�O���ge���8�gT�%[M�A�q'���?ּ��@��r��ǰL��/q����Q�~�K[���-�|�*A5�C(TM=b�l�F�