��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��AU��iuɱa�]�=��w�,s�J��I���\c�bQ���lf���H}���Y�RCv-r:�)$�u�z�@��f�4[�">�7�����Ar�o'�tWLc��P��ϭ��ܑ6,h(�
\@��ԼF/IF���l�%��}-P���f&�~r��YY�����1����L'�d���f��>��l�^0�s��J��]�ߕ��;�u���/��������*Ռl�K��c�\İἫ�L,ˤ��3�����믽I8Dd��ƕ�_��
�t�:xtf��$�,����� H���\�[�O�����t'ɱBM�/'��-���\#W[��A��"�x;^�̀���A�K(�Ѧ���O	�D��5�bN��O��z�� W�Lu��9�r��U*�؛�V�, ��v5ezi��P�����_�@1x�(�;	�ب��z?d�C�z066�䜗3�>���0�˖·2�ʎ?c�@+z�ƏtYv��2�MS/<ն*��]��t�Y�1k�`
�g۲�a��I�v��wRY�V�5]-�,�GP���&2��d?$�/����݉�`� �-�у�mد��:��2Yu�i�R�������_L���M*F��j  𭢌��J��?e`ԍ1��Ol�E���?��mȗ/5��E���6�ܧ�Bm+%T/n\��9�<�f|�'�}k��#�ψ5L��I*���.�>���A����]����|�NW�+lo'3E]#b��Yɯ��/~>�%���T�y�� ����r�_��Ir�-2�,ˉͽ����Q���8�;ۓh���r&n�y�R��Ɖ��#	���00�X󴆛��s)<��ا^���GQ8
�t��PI}���%W��h���{�C�T��*7vh���%k�c2苖����]h�6���.������L>�FHo 1l8۠�E$�Z�Pk�HM��wIeU�s��j.������i�L%�z���\J�5z���YN�@j�l��w��>��H�Q����N��4Tz	���Fp#��n�~1w�`k�E�MuzX^�X�u���p9�m��ؔ�K�`��v�'5	0�0��X��c����J';NU� ϞG�;.���+8\������	DΥ6kama3���hu���N�Yr��B{p�߯�į1�#��/Z�Ă�k,�h���1����:��	K3R���;߰�����-Z��N�;���t)�#���0�ϮY�c�	�uP��IPe%�KF�b�x[�@pt��=j�l�����<U��(�}2��������6����F�\v�gs��,[��ϳ|��u�|�O����s��D
ʢg������5��4܂81Y|'�/�|;ߤ|�EŢ��hT�N(�ڃ���&��S�IŲ_U�Tz�R������ǿڣ��6ւ�
ׅ���h��P��HU���5RF�P���ّY~*�M���IIC��7?��.�F}��e��P��fsPÝ��bB8��*i�	Ro���t��dg�Ou��l�:����mNbUb�DD�Y����V�I.,Au��"��2~:�KWfٔ����c��0��,��a=?�q��z�`>�^�o?�v�K"�ؘ˩��~X�}�(����l�w-��4��}B��Yp)�j�V���K`ehĺ�=��z�n+\�`:ht��{$���^ ?���v������B�=7�Jzvj����)�a�猕�(��� ������� �;�!x5��>�"���:
5b%I�}T�<r�^A������ʳ����28�[�N�e��mߘ�p�Ix8�ք�j���9w���ρwO������NK�5ren�����k���R�x��hv�:���V��d�S��G)�q������s� � �(�S�Q���ۣ�ʻez�߆��s�A����w��񼋙�/n�TĶF�;��F-��Zݯ}����=P�m5� �Ȇ_�`�2e��j�IS	�#|����g$���E����PG.��򽂋-n��+,ݿ�g\�+�B�����?";�0��q�b=3-�H�-5\G�Re"%W����e�Bޘ����	��#�Q�q�$��IPd���R;(zu��h�A
F�?\*��]Bv�W@"����P���1C�*���v9P���G��������/T���	�=����ْ����Ź�r�VnE���R$ɟ���%I�'��)�����5�b��p��Zod���i���{8�!�.T��t��;=�
$f�]�����L�n���u�-���y^P�u�Tl�*<��6b��Q��M�6A�1����ߛ`�����@�1�n���٠*�gY5�S��|���;&��|�:�G�����E�`)��8�z�N|H%[�]��;���4�����:����SVX���~�c;[�f���;8�_��-�d��=^:�u��ǿ��]�Ilo'��n���1/#�q��8eT�Qbo�Y� ���ָ��N��t��]�ٽ�0�Ni�$�sЧr^����6x�EФ�p�9!�t����-�b}\09�KM�sTPf%i�q�&��T%��
I�D�E���%�Yy�-NؽuC�*w��~���{{C�Q�~�'�C����¡w݋�%'Gl~�k���6r�Cxb��j��v.2r���Nd���m]�kU���]�,�w��K��SW���'����\�B���¥��)}�#�Ƭ[�.3O	��g����.��7|����ޥnY=
�]>=lG��D�"�uX��k,ț\��Y牊����/3yCnۄ08����!�}G��u����,:�k�y ��vN/L�m�V�}�۹,a��'��rҔ�d
���s+�"�_���%ƈ�Nt�yE��8ߘ5վ��svBZ�ٿ�{x^�U&��u�:�0��
�wj�����RY�����T/��8)��������������O6�瀹�O�F㎺y��!�w����F�����4�f�M ���ls�2�垹Ϧ��wh)8uv�Lk�N��6���<�LS�wE��b���*2d}��u�䗇�M?HgFDWd1<G�v!\���!v� �p�~Et3k�+�ڗ�{��c��tDGAT����~��Ăƈ���J.��z�g��~g7�0@I<�:�D����x��J�m+,�������h*=�3� ��e�[5!Zm�n����+�2��������̿������q$���y�:�`��ع+�F�(��?�2�p}_�dAٝ�j�f����T��s�nNDv����mw�g&��w��B��FZ���X�ST�w�x��7�y�'3�./,zE�u�I�<ՠU�Fm`�D����Q
�����F��5�Ҟp�0*[R$�~Qg	�8a�u󼁴�����&�2�G�#����o�s�V�I�a2��%ę3N��)�)\��]�M�;-�ɏ�O]@r6O��ܠ�˪�IJb���\H+;�
݋sK>'�г��F
WS�'�r0�� `w�<E��d��r9bhG_zI��+�ʠ�����|��t�9���/!��|g�sz�*�7�=�J�S�Y���V<�8��:dw��E��5T�%�R�~�b7�����q��|Sia�Ea��^yGԺ��8�%!�<����0Ƚ�Be߅K��$�c�<I�SP�:�\ޒp~�����Ԕ"<a�q.�g��V�
��D�R�{6�Ĭi�{>����'wCR�>�6N3�,��?L�Nգ��O�"�6su�j�o�>���qpG����eƆ���t �A�G�3Z�Ż��"��g��v���!Ԃm_�O�˚��G�С��(���9R����Ǽ�ڀ�Gsy>��K2i�M�V�E �n"4�np��=!>�6�@�кx^U�p,ӹ=�H�;zE���4Ũ:o���׊P{���t�L֗�#��"�~7HMW2�F��	�
r.������6P���1h����j)�x1���3���咺i~�,ΔH�t��YsNXc�����x�fՓ�D���$�m7�i8�U~~������ƙ�=-2��7W�#^i��]�A����nt��^(M4��`'�g2� s�E脀fC�E�V��n��]�I�\#:� ��8��/��(��k9�yE��"�iZ3�Y��.,*.�.}��i��o��aV����N���=Jn�j�� �ck����0$�4u���k�ru�2�U�s&�Q a��t��5(<���q6����\�V��dDyy�(���Kt��k5�R睲+z"�WL�*[���^�|W�lO)	���@�O�i�=���EF��w~{�E���%����x�� ����	()�X/��7z�~T�,s�a�ؽ��{���HD����g��#�R����HTg׻�P�{s#A:b�h@�R����%p4Y�w��Xi�%�oe�1�s�q����[ _�,Ì�bN7��y��np�1yM?�8O���%��#���ت���-!����;�.@G,�Hv�gqN��&�9�"8�rF�$��
�p�Q�Nnw�	��H�]T��pM�y#O`�K�!Y@o���V3�Ϛ����$��.��[���V�,��6�9RMեw+�9�4��Q��t��.������T��2|< �>��'� �u�Ѝ�@�V���y��H��N1�?}6w7�_xS�ۙ������B�d��g4��O�B���^E�9�ol��$d�,X��n���kb�~��������ޏ"�J���u���h�v,��O���D�яJ�����C��),Fİ���.Qr�u��Irf��jxp6㋻�簳q}�fH7*%%�i�z*u����)�B�{#%R�RF�]Q> #a'��$��/�&�'j��&ʦZk��;��`1�H��TX��QO}��s��~f1(���yyhV���~�W�c����ݚ7�T��J0���Bz����h��p����3��W�͓�&���ma`�1���� �T � @Tv������R�4�������|�LRT�L ƨ�k�E�u{i����h�O�u�ӗHq�{�8����ڻX��Y���t=�v�|���:�����A�m\^�j��[�,=�9�^a� Nb�͋��=�j٧Y�g+���A��41l�7�ޡ5�Ů=��9C�����&��g�8�D�U�(Wq�&y��@YKW]�Z�4�d�6�=�b��W�3F��8�'�uTX)���ൽX��9� �R�<�ث�_T<Õ)a�=<r
,�yWw*�}]�������I�|bfR�7:yB'��1���iC�X��Y��YE����>�= W����z���Kn֝_�n`̸�Ϝ��V��pc��Dܵ��ycQ������1͑+g���d�^P˖����M7�9yn=셦�X9(��#�0����S��]6�i��%�9х���r����Jt���F��]M�ܞ��7k�'���X��QO>%r�>�TS#�;�.e8�o8�*ڬ:3�9�O�q�}�/:�;w�Έ./u=�$��ꃿ �6&�T����I�u�//�G���=U����*`�#��fn�h/vu(WY�ka���O<"߰�m����W��%v=,b'�p��N����i�Ts��Z�H���f>�ݸx�f����q�.7SOtl	:*�f��(u��1����4��v�����wwNR�"���2�Z�RK�}�Z�����!���`>��
ب�N��SۃU[�h?�ku2WV0�\��ʡ���z�i�b��/�z��wNSD�Ҙ)����l]���fk*��q>r@����e�����9�HzGSv:̠(��N��I���Y���1��A.q�!�gn8�-H��|�����?���y�t� {Ј���x�Pi��₃�/�ҫ��?��h6m����;]�4�)D�,Rzo��:���t�v�y�b��6搛0��F��@)kA�ќY"Sx�7к�/a��W�)�uZ�D�]�35�I��ƦZ$�o-ч|�.��$��M;�'̈́�N���k(���	� �Su*�k E����$9[F,j�s���^�o {������ﵞ�房�\����xz�`��p&EVcM� [�7��%`�zm#�h4X/ܩ�׎���w��ݠO1
.�ц����aỹY�U�6�;�%�<Y8���(+����ջ+�A8�Ijw�.g���Y5������v������yvV�N�W�X@--Bß>I:�N���tvA`��-)����/_`�x���p�Y?�_�x7�ԇٲ(E����Ȥ�p���tF����/���C�:����c�)9&��5��)�~����D\��IC���+yK�.���Q��I�M�ab��Z����J椎>�"�߽�|#雘��"��"�����f��"��Y^|��*���QdJ�'�vq�"�����+z���WZ�|�ي�=W��n�0
5S��꺚氏�\��`��V����dt7�,h�^Bͻ�צ�FH�Q�K��(�.�
�#GB����4��]�Ϛ�P�6��@���ج� Cq��(�`�7>��~cȋ���?q���$㯤T�;X�
�Ay7W{��݋�!>b�g%�0��솀᷐���,ڜ	_8�	�w����Z�1�'�(u��`9'U2[|o	�ytt'{��z������O�4���X���~Df3!.c�>#�f�3�I���f��(�vR|���%L����R7�]�~��jg�f$^7�H�̕u�y�5�$A}����{��1}�w��َ�#��X�
�4����[�� �,�5�(�W�V"=��0�v��
Ü������1�H�S���o5�{-	�2�R���'�K��x�ځ�7�p�q
�t�z�wQ?Q���29�,�G\�W�\��ⷜ,���1��'�#]Eh�r�q.3��i���%�Kb@�Z�t�#(���Dz�<)Z�;�����?�?^����#�כ����X$\�I�w�����՟�\MS�0��w,�v)���:M�u��0�h\�$J�_'QwJ<��0T��_ҝcM> ��9��r�_M� �m��J߯5ѵS��E�X�Qܴz���&J˙��[�~ZHJI��D}�s�h��vI�m�z���P~��TCj��av�z��=
������w��ɯU���l��+I�,�Rt�ꡋ��#��m��!�"|{�s��W� Hs�`�ף9����+�����q�k�W	iMG�� �Ô
��K�_���! ��-����lT�n;��$���f~��f���§Q��ϋ�ǂ2.�iĄQ����x�He�.Z��S��?��rC���߶���7%i�0����(�s~���]�`���=��e�py57.�U��ghh�Ap��G%�ͬb�q��S�{�# :�s\��T��>��.>ā��5�+�n�McA>�5�1�6��9�{]����G�5*;�(��=��������+p2�Fh}<���"*��)��?�9�5XAlCM<t /i�F������룐o�M����BJq��a_�P�_9|f�'q��r���`g�jF�����di���̲��ua3��25q��c�k�At������M!��nio�c7Z�cmd��:|�ER��t�ó�p�I:���9ɇ��[�\[5�j߃>��<�P�-����ח��/���m�H/<э��!��䞥jl��+�!B��c���szWUs��L
����t����Zw���Q�'��($���#���!�9�I����e��t��T��)h����VpP;ska�\����7jz84�}���Ӿ<N8��7��q�
��?@�t�/�����&��I�J�2�����i=[�p\�?��CT���_����U��" ��dN���X's���r�&������}#�7wU.��ne������t%u�8WZ���{��������i(����g	���gx��d҈�[M��\b�2���XX	��@�Z�rɻ? 4��d�w�#Z{&UC�}����X�q��W���K����AGV�'%��ݙ����
NΞ�̔��%m'8���ЄB��<��zb\w=�D�9C�x��bQ��q"]d:��z@�zN�]~�����ZZ����eyLK�7���\|�/���+]GVxωEgg�|���*f��%B�4��Go�'����ܣ���������&�S���|�f��/�7�F� _����a;x��0�9V\ u�m��
̛��*ٻ�'?��V���
�� �mT�کa��GM��7O�	n�$���X�
�=Ў����H@���52�<{2�!�9�2�.�H�����2��ٷ�s�!>}��>�����T+%P����&����d�+/�=J~��<]�`�K�N�.�����@;4����δˇ�Ut�%?�mJ�D�7`�:�t�M�Γ5��S�+�L�#f������^w����-$t|^Z>>����)���".{"�{�E���uERź.R��@�5h	��I	O�}m�
��wm�̝ca"ڜ!�#
�k�3���:�O�b
>8sM��>�jwֱ���
)O@&��2C���
���~Ga�E��ZQN<v��n��b�j.�:^C�J���
�������G���(�Vo�L�f8Jx{?�X�4)�~��i,Ms���Gd��C!2&���z)
�����?��G��M�IYf�@�9���
�q8%�BT�F��� x��f���W�U��z��%��Sx�YG))8���f-�Y�`h��ݹX��S�y��n�d�w��Iuao�"IEI�V�@cD�_���mˠh�OJ�q��$�:���7�s܉��2�^C�crF���<���{��ӧ�\0��Aɛ}��v�G̱~|�c!YdK�{�`z��2�(�-�1s��62�tN�UM�+*�0A��
�1 ��|X�x�Jqf�s+�WA�e�5h�l�?��iiDV�{=yyL/J��U�^�w⸄��>�� ����#s����I�>�|���l���:�$2նۂ�Nj�}L�S>��\g��S�Q��-�x�tRg?�^Hcg�qs���x�b�]�L��<�+kQR�+�e;��LB7�4�%^4ݓ�n ��eJ�[�vz�VY��0"J��ώ-�o�����ާ���\bSkZQ]P��ß�Z{�m(�N�]��kV�oΏ��k:m��)��R���yTM�5us�3�C �F���i��̂8�l_Pmӛ=�-ա4�mY���R-5v
3�9�]A�6�-k�5�ga=˖%�51>8zW����DI:|�	ߜW�D��#� oaΡzD.�y���y֛J���^���wa�O+ �H1���+pʅ�P���:�v1A�0[�2�� �662���$|���W��/�-��?ߐ��^��Q`ܧ�C�Ѻ��m�T��8�=��.��r�?$�D�fS $����7���&�I|+o�6���A9g�В4��}���F�<��#�<)�Al��5�7�ߋV�d�AB,���oz�֝?�O?$c~R?�4F��CQ7�G(z��q!���Q�L�&�ac���b&n������������	��C�	�ņ���֫�"��r���$���	��.##��fS��:~,���p�p�'��ㄙZ M#1j�h��KA����C9*�9p��.�7�(F�r1��@�7�T���4⡂�Q���������+q��r�6�X.�Y[�WV�J��^��>2+2�SVK��w�
���0!. �����fĥ`8�E-��cj�K�.c��J�,�/F2f;���R�|&À1Kǣv��<>*?1mܣ@��Be�� �t�c�bC7�7�9�V��p�sglC��;']f���28���O�&�39�ݯk�*t�+P�\ �L��b����\�y�򆀅��8�ן���g]������?��f�����,qŅ�$LQ\��1WQ���Pg˭wi F�ē��i����������+ُh_U����s���\#�b�\���=�_���#v6[=&a��٥�H�g�l�c�1&C7�0^Q�В+��k��u"$���X�M�h�`7
E�؋n��-�(��ݦ���0�M�E�-?~�ڝ���j�;s������o�޴5�'e_�V���甆P"�-�/˄��#c�>vA�]���b1�U�7��#�SԃT��lQ�������%����A���xd�k��e/ ���8D�UX}��Q�P�N����F(���4a4�<��<�չ����^B��z/�	X�E���&�]����!����(��8 �t���0o�4߇�l:H둯��+����\;c��H��ǩ!��r��c�}��ٚWۊo�ΐ�9;�]��CC9s?R�^1ƙ
�@�I�
��P�	������(�ܻ�H����;�bk,Ԁ��	�=�nT9w���0Η�kp��k���!km�>خ�wQm ,��ޅe���,q���ʛ���;��L���Fj��	�h�}�������9��:��i��m�_ӧ���E(�[�����C��R�����kƷ��1�A��a&/k�R:Է?�ЦN �E���hFU�����^�lqVKO�zWP��Ob�o�ѵ��/T;؝㷠t_��R��&���y��{��*��RH'�~͔oyG8���3�p�i�������Ⱦ=e�j�=����h�v���d񮹽0�?Ҵ~�������5)Uz���W���`2
#�_f���dU߬|�K9d���0h�[��f-P� �S��Uz��ٯ=V� .v<�1�`|7X�p��ut
V\�L�T`ؠW�[~�ݒ+PZy���ؗ��U��%k��YS�Vw���w�#a(���S�S��Z��NB?��������(����}�h��b>9�j�����I	l�Qxٞ�Cn��gN��)*�筕YT& `��质^�|M������j��%�t;]��ʔxp��}'7�o�)%��t|��^D�d����{^G�Y��������Qv���X����mcf��)�d�5j�罗��p�U�mӰ'l��=3�	�*�^Q5D#�jy*��G��ѫ���y�8��z�kOVa�ѐ
�<��(ȣ ����T���!xw�P�I�UY��U�� S��Jf����rj�0_����_e3��H���c%���0`|���.��ޜu~�H��e ��F�Z`�F=6�>]P[k�#8�o��Z����|����F7�٭Eq�s2�FK;D�y��>���u��"�VN�>�V��{!�H�*�Ue1)�ϙ�w��z�q��ÂB eq�ϸ�<AV��?ۖ��� d�g�}C���jw�i2��J�ޔ��Rw,�U��uCґ��S-��7H�Y��EHx_�,�UY�!L���|�?�����>�,	�^xep�#��S�hp������'�G|3���Pw�$�O��*�s�X�����f����p����Gz��`�J.M�M����pJ�Z��WW�/�2�.�R�1��]�A��Y%#'<��n�Op9Hnd��$KN�pR��:��5���7��ކh��iz�{�Z?��&�t⒢���%�UJ#�NAS���)/D9��I'�`��mVo�ؕ���V���Hw�f��U_��u��և�>��:a ��0#�u�&t+�4�a��n�
����U�x\K�*��T|�^I��%,GqC��,w�ﾻ�=���Y�f�5<��[����d/�Yn�V#M"�,�yJ�K+oIO�C���%p�N���C�)&�c��T��=ρ7F��F8�x]���y��w ʟ7*b\e5��[���#b/�A	T8Wo��Upe���?M��Ca��W��=!�����U.������3&�[���\1�L��ԣ�^B�6չM,����������N��Jr��)�W]\��G����|����^�D���T�3��*��|��g�"܆,fb�Ȥ$��� +��7	��T�3��wO���&���Z���^/�C��ǔ���u<S$? �����g��s�G����d��	����B�Ŀ�i���a>�]�@]̣P�}�\43����Q�T	,�a�c��:�;�ȩ��C��!�;�B�>�����O��_�����V���$Fӆ�P�q��آ���.�r��D�J��	����C�Q���\E�od���3h*G�^hN�`�`���ad�l�
�%Ar<\bYD��a�MK�F���+�����Q�)S�S�\�rs�奠��q/�Z�EBW��R� ł��`����H|��n�т__$�_}f)R(��T��AG�Pv:��ps�ՠ�������m0�2X��=��y?����Ѕ.�}z)���xKu/��w��X�y��%��nf�@դ����A�k���"�h��EWuG�gRde���Ƅ�R{�Q����.����6$��3<_�����.E�Y�x�Y�$��(�}�;��Hv�2`�o��33�u?)����(+>Q5�Z��{�hd�7y���eU���� ԧ��>a�����[�?ƧN�g+8���0�eO���o!��p�߁��Ԩ6=�k��z��f�z(����$|,��!�I� ���������0
���=����P�x�A�^���F�~ī�w1pA��lp�J�����q���=�b��0�Y`��9�÷����|����g~�W*評y�#qq(����B7,�Yy�.o-q8慴>�=�����2*͏qYO]���t��\v�3��\ș\���	�y��A��n���~s��8���ᙕ�I��F+����~8�V�|b]��.�;*��+�Պ�� b��v÷\^U�f{6����.�m�$8fX~��f�j�/˻�A��g!|�2T���ցn�9�� I��H9�}�G�<'��Hȁ��l�m+^E�Z}�^������H����HY�]���ڴ�4����ԞM�\qsI��8�2�2ӡ��i���K�7���6k3�IJ{%͞O]B�"��<�� �F��㑠���In�V�y?����}�-<Q�҆��xԘ�%��o�̦�TE�pe�����a�25��OJ�L�2����NSA��]�[��v��ǫA2��DQ�8(�cMQR�:���"�gZ��$�������<����\�e\��>g���>W^4-�6�G�ٿ��u�e ��fF��~ޣy�T#U&[��'��2E�S�z��<K�8�R��u7s�Yc�ٽ܍T�+h(��QF-ۻ����
��Gs2l�R]Ro��z��Hk�^�H��C�,Q��E��,�ܭ�|ԁ-Wɬi�M��:�&O�OzԎ���_TW4���{.��_��)��G����螷^h�U?L]^�(�?���d��T�E�%M	^,�Tc���u\n36�.�8YEv�i�jO��Y�b�� S�̕�7�}���/���T�d��WIh����� ���b�K*j�ιTM၆�(��ɶH�QDF�u��P��L4���Z]�6|�4J]/���s}4�{�˾8�9ǑK|�����#���"X�}MJ��A�bo�.��vdM���������Îp���获�9w׮43<���Iu�m���r{4�y�]�ENZ����㣖i�]?���f�,6�~�z��T��@V����O �D�K��0�yn��M����9�ɺ(���\���9}82]|c��Bʍ>�5m�lwr��x�VF���D"?�O�����n�n�5�[�P�����$��������) y��!%n��m2��JȅR��'Ƀ!�M̔)�t�O;|C�#��/4�΁5v|h7�l�Uq��(x� �m�߫Z�-�<i"�(ug�1���б�T�ya,�n�tm�߬&�imOS��k�F�����o�:��]s߅�>Ad���_k3W�Q��Ɣ7ޗy�ȴs�*��� S-V0�d8��xy��x�)�	�^�;�̕e�>#I�W���7a�M7cj�:��5�t`,PV�w�K��4���R��8On��ƈ�����"=�|��C �r��Q������:V�͡��y���e1TC�]�N[�?[��p%�!M�m����g|H�m|h�b�uBgI�L^u�mO�B�����ϡ+�~�i8]o��o<�݉��C���%RXE���4-1H��LR0Dx�T�&Qa۠�9�Q�.S����|����S���%�e���y�)�8kӑ�27���R��Y'�@���*D�0�;�j��N��"����Up�O�)�a�����W����L��!l���Xɮ����rW,�ф�2p�r��Mc��j����6��"�+ՕQ0���=�,8	YV~�~����oZA�5��J�`>S4lMn-��/�����O��_JG7ҝQ�$<��,�#9?�Ə|�����x( ��Pn(���v�%��:��U��{����k���b
�c�yb�q3o{�(��9��� S̽���!l�$Qc�C-�܇���TN��dP���>j���]�7L^u�mk�����y�A��MT�D��Jq%��^��n����\�ӟZ��(z��.��<��&��sê���|;�"1L.�A}R��l]ʋ}�"�s��w�����] TGjŰ4!��x)�.jr�D�V�'��aBμ L?�s������I��\��k(Ǎ��V�X�8w�sf�,U�z��oJ��{��JɄP�'��^���9�{ 3�M<.O^�W�����f�l��a��)��P!G�׬dj��.����:1}Oț�;	��!���h���v�q���x�ѽX��[�)�B:}OÄ!� ��
a1���_T��7s�֖!����^�D��=�Z�V�:���w�5�jgp�@���l���&ml��������~���m�%�)���m��I*UC!�]6�P��J]���r^�,�h\A��ʁ�K&A�֡t�ʍ��9�6Q��V�`��(���Q��x[+\�;RM�dn\��,��y(�\D_>{dK��D�]�W��T�1�����a/���6������O���}O|���u��g��E� ��'@�J)ܡ�<}���o���;�r���F菖x���Y|�*	i3ذC���	l�z �����j�u�BE1��]8K��`0e�kr�M.%:ax'J�B����s�8Cfv|P��ԣ���9�H�h}D����#����\a	a(���cQ��C�����-+t ���}��w�T���Mۆ?X�֬;e@�|%D�rN^���w���{S�LHy�����^�0�� ��� �ر�
��POG�'1ρՀ}\?ߖ�|nE-�8�p�O}�� Zx������'�Q�)E�g%�!K��յF� ���]�.�t?�B�[����f��i�_z�.��?uC�i��ai�T�gd�qds�e��n��C�󩤤j��v��W/qA��\ab��¶w`�����^\��8#H�~�+�g8���ݳ|�~D|$-�[V���+m�.�t�y����Q��Ҵ|&}�x@LX���V��oY�Z`��!E|6yP�s��70�>��ǣZ�F�v}.�w/2I0�L���g�Q8H��>�TA\�[����{�tO{� ��7�;
�a(y�RO!����i�j�BY���C֗�����H���N�`[z�S�-tY�q�$%\)K|��7��@�z�j���o�;��F�\�E[�&���-� D�(�~�����������I7�=@�IB���1��Ɣj͆R��UL����LM��%Y�/D}
�G,���_kH*�&f�&i$?�45�Ғ�Ώ�I�` ݵ�����8��<�S�p���%}���jJ����$''��w�\����I�Qd������u�ǑEW�"�sr4��l��
�2"�� s�L��9I|/@b�7oDG���O��x������3�x������~_
�����#�:u.�Z��G�Q���B`�n��Z�@���
�uY5����К����Ѳ�їO��O�"�,������-�9�RZ[���EKb���OH$$|M� |@u�!A��Q�r%>���&���t(������b�*��2��?#&(�\F��9�=χ<Y��).�!"Ԋ�f%J��z��ҏ�f�f��q:"1�I�՚&���S�z��m���$xT�h��7U�UV�eB&Zx	��_����h܃e�E�Ҿ�I�0�~�!�}���S_�7ě�xx�P��#ε���"�h}b9��a��p�b�;B�w���F���|��&3�<�tIz���|=�j݊����hp3� ��TCm�R���+���i��=T�X�E_��(�"����������+���,�Ѕ�)�����q�h~�b����fN�])�
��dj��))/M��n��/�4t�O-�֜)/�|jo1��O>zu;�$�%�FK3�6W_*,5T�p�_b�ɬ?hU��H�hG2ypp���v�S�u1V����רd��O�W�3���������H))?�j��*Ԟ��\V柿�3p)qx*���p�X"����|����ܼ��j�z��{�~|�S�������I�^����BQy�Z|Jރ����� r���#��hz*�ʣN0r9��N?[�Z�}q�3@��6���)��-��6t(יZݽ/� �l�G�z)��d�I�L��dw�8v��h�N��ȧ�U�Ǽ^��*���!��cF���Q� u��?�6 ��nI7)��:cպ74ċ}ڌW��;l�c_]�ixٓ0U��i�xu��p���S�����3��C(D�B*'ջ����X�|��[��J�Ws�d��|�#�{"�K��T;��z�g��G���H�c��7�b����c�X��@>>�����E�)`%��T��>mmǍ��Z����P��1�z2��W1nG,��Jķ����$80��C�
���x�m8v������'ܼFn�׍���˝^��QL���R�B)�T�߬�ԙiR%_�<�O^��+ԢU)]eW�������y��ر���h_I�ȠU�v�p�!X~����:��E� N3�J ����o�0�g���C�'��J��v8�D�������.OD��r�<*@��/����իp�0.�!�2����r��m\����Jj�D^�Z���O}TP���ĩ��ʘ�,9�||�o�fMU
>�σ9�oqw O4�єV�?���7��X�=E]H~w2�����y�Kw��ǽ�TpB�����1�C*&�c�M�O)�M�=��g±.7:���|A�|����,�	7p�����?�����K��,������5���|�����-�!��ݣ�q�����M�Ha��)�v+���Jw�aX�KM���i�~�V�/Do����~*���H�J�HԀ���T����ݪ�z����&,�F<�]j�Suְ5}�'��2��J��4�-�搋�bˊ�;6��2����I�yju�=��AxM�}��}kB�JV�/5��=@@-�N����M,�lгEn\p3C\�7X&Ӡ�ĥ8&n?nbC3E��9 �e�Ֆ[/\@0ͦ� 4	�K�أ����%/�;��"�:%V`����Y���f�z���`=P�A�wY��vW��>�Z�Y��sC>����W#?���d/"��EL,|�;���4��ThH<a��7H������^�+����JN�n�R��eL���y���_A6��xS�! � P<\�1\U��$�N�����Y��ok�j诧Ѝ�R	�
R��'z��@)�0�!Xd��d)5�GD�G�m'		0�q�U�$���	I����ς����1�V�{7�;����G+� �Y#�!�?߸J�?!��8'����)��8C�j?�X��er+��<X�@�,�������M�W��{�9[C8}Ҹ2�T9�W�]��9U󣃼�K�Ɓ�Q��@�O3+���s������N�6����k����8�8��~sH��z�Cq���oL�v?��\�=\�@�~l��̎�>���s��Յ]��G�GR0����rg��v�晝WwOX2�0������^��]g�f0��Hb�շI����h�tC�w$���D����]t���+>���3���6ٞƐn����ڷC�� g�����*ߋ�O����ٴ�a��	o�2o�2�h�h����:�6��g��>�_����1j֢�L�nz����6�I������j��]lZ�?K�8�N�m/`�gt9��
tzb�!�G;8��s�3�R��NmX���W���1��.�	��^|�u.��p�O����֫ϷZ����s���rq�NeL�`��HEϸ��)	���f_�����a��'����t0Az��o[�/D�@,���%T��T����š��!��-�MϓG)��;���׌��
�Og�8��rA�g�.�7���]wd| Y�b4R-pWӧ�?�n7B�֍�v���	�=��N �\����:�y0+�yaK�Cg�,����z��==�Y/����n��@�h�"v��1�6�$�p�D�D��#�1�!kbm�,��Ǐ���S�;���t�����8:8ǋr P�&JW���>�����'\a!���,w(��zD���F�k�>�->�"��IJ�t��8�Dϝ���BoG��*�<V��5
4X�_�����D�@�n��{�U�#������vͰNM;%�'1�	;��?S�G����ׅ�^�x��am�[C��,��)FQ����m(!y��\�\}�������O�p'D��Ψ���	�6�|�:���@ D��ܩ�h��I��\�Q��-&��a{�a�rA4O~��>�:Z�"�䠶(le_�8���'p�"�t�*��{u
����X=ͯ�"��)��u�j|:��?��W��EH����#� o����k&4��R��p*̆��p}G����x��\&RC�.`�j"F��l2��Ʋ���6��`�1!����=�,=�����t,;��h0i��sYr?jE�����[TVTA�c+���)7��J�q?X-U�Pb��ٯ̵zب�
+�X��
\%3��]��?�8��2=�JB��TگcFw}���r��y�3���" �|a����*����ʐp nu������6�0���/n�7(24�7H=0ח%BX�����Dpa¨G��鉤��[�o9	���v����3�M|J��WѢل�n�����5*<nar�'�x���w"�J���w��G���G1XSKx-y�.��O�A6*Z��q�{��l��g2�U+f�/��Z006TLXٛ4�gC�?Z3��F!s-�]~������P�W
�����H������� ���u98/_6��Fiܤ�wZy�]�+��uu��K3�(��G���]�?��-2��3��h��%,Bʎ� ��+��wv����:�&O)-N�?�B�d<���n܉6��R7rH�]^�V���9AI�;+����ao�����b���"L�QE��T�V��,���-�a�Y߃�L�)|�A��1�r�g׵&�$]��ۃrj��a�JߑJb]+�A�P=��@��l�sQ��æ�+�d&7�QF�V'"��dŕ���ؤ�I��E�|�F���l��\Pϔ"S�b5�._�R���.U��|�j�!L9��i������T4�%�n)>���MH�i�;����8[c��E�e��hF��3h���oWs�x|�|:ɲ+>K=�1�9�)&z�_��vo��kV]\�M!92�0
B%^.���Q2�C�9T>�%ِ��+�"!�{�@�Q�s?S�s��S2��;�qK���R��&��dus��|w/�J���fR��*��nGY��'nM��al�E���h�چq��(������EM�Ul�e��^B�����06��_
�W�]6�|�s�i�b6~���K�C�*J����mDi�r*K�V��˅'��ϼ�OX�dC	���
��q\�OQ-8]�o�+w�1|�s%lM�s�01�����&
���A)g~=��Λ���$WCKч��zŉ��A;a!r�ճܘI��{�Ɍ�57X�gqH�Z���=�4F��jc���ree����&'���]���)&��� XD �k�8n���Qlp�+�����V� ��9��2?�$cH��[�4�cCh�M��8��7�E��y�kU�0�:��z�8�o9���]>��}{��9��ӂT.��,sy~ؖ��~�������k6[?]�ƺ�m)�^
A�^�FCi��:=���:?f���ǘ�ɣU��W����X6�$���]���9L��ĩ��և,��L���o�����x\��H`��PlȖ��S�x���@�"��REg������*�7zcE�=����QoW���(�d���	��j�_�H9�컼�KO�I�Ls*gL��b�x����qIs�J*����|��uRoZۺ����U]�U�M��|��¾��֢���GG:����F��g��!�4b�Ԣf��NCv9�ߍ(*bu��݁�4)ez� f�@��!�A���������;�_cYd͋��g�Z ��j^����t��%u�UMH|��0�}�Z��������^|�̟�vǆ*C�ѝW��l`��V}��@2�T�
\�ٔ1��Y���G����{p�h�e������\�z��k�Q�S��B��ú0Z�S��>_'\�(����Ee�����J�X�n�C5Rt㝢]�U��{���W� z8'j�"�� �ɂ���EE ��������(.����`ae�5$���6���;�i�9��̚�]&�D"E:�����"c��1Zj�#�-��re�NԐ]M\ſG�h���C��YQ�{�*���Z��{�m;HR:�����S���&A�U��n���7�ξ���P=�� �[���Zs*�򞆄g��� E�f��{�n��snS5�aV?6���[�?�r�y���W��k:�\�p����w��L!�;��j��g^�p�����j-�a�(r�����5�f�Ƃc��{���um�'�6�W��m�'Fqz�s�1��8����8iէr��cH�_R�].�K��_Bq�Д�:P4Ţ�X��ȭ�6�#l�]�l������§������X���2���0u��s�+��;/��.nīZ��a=��L��7��]��E��y'4���I�s�ސ:�<Ў�7x�4���<�����<z�ɼ>���4��i��Cx6{@�'�	��X��3*`q!G��t3A��"r��m�?���/�(Uq�r�}qi"��E'�i��"\����Vk��*�a�P�,5�L��U�� �rb�O�j�JƫC�\���x�q��w�l�����U�tS��-r-�0j�e�������F��i�"�;n���(�.e4�(%��*� L�G��xDy��� ]�Pr��4��	����	ro+�p�S���dẕt��M����uY7 e%=�:U]bS>����A(�Yh�n��@���+������L]�)�1p�d+�Mg�}�;�$��?���nˠU&��9A�X$�˧o ����8��R�`aU�Bo����w��7�*�^��a������:���:b0�c~a$!�:�єW��a�%3R8vE�Si����
C?�S�ڮ�]��=M�&��� &\�	�����)l�}ņ���u�)ЫТ"E���Wb��}���I< �mM�d;�2�]�κ�lD]!�Ō����h�L� ��Su�ЛLo{�֦�H:\�Xd."���b'��ޤx5�)2L�ޙ}��k�l�&r��ip��"���n}��2��^��I���bY`��8�Q��� +���ڙݴ7�H�d���C��-�w���^ ?۠�"o�D胡oY�I2T��}Hw᠑��,d��o����'
�,�xb-��L��Y:�,�P��a	����`=��ܹãw��`�r�U�)��n�"�S|���\Y�&�n��n���o���4i���(D������#���R�NB�S��
mM֨UR��#���&�� �5Cu�3�x��-Pw������I��foD!��V��f�e��b�U�C��d��{ZNE�v�S$J~�{��`z��%\ ���u�kI����M�3CRr��s�mw��Z��|�0-���H���W�W��a��F>d;�8��ۂ�U\��̶����렍T����p5���Z�@�?%rx�<��?_�u�̸qeˊAEh�.�^P�Ӗ)���[�*�1���Jc[&�"�y!TP�]>��H��jKa���zX ]~  ��]�������L��l�~��;�ݛ�3L�~�Y��͒��9]�-sʧIB��[��F�^��M��v����U���ʹ�J͆@�͑��z�>D��6cQ������?V��ߙG�oE N�k\a$�fs��7�A��C�F	�d�5�=Ɲ���B�ٳ��~�C���UYG���y��u�1�鹢x �@�>i�<��>=�̄���p=�I��A� a���+B��¨�mi�G%��[=��M߄��!"�?��o�ՀxJ�����U�Y�����O�+�8�s�~^�����0r"��* C��4.x�H���$�$Er�z�p�u��h-�= $�F�������a:]������F�����P7|����g���,:<n�2�"*0R[S٤��H��{��w��6���p���V���ć"N�`<ޛ���N��
B���: ��R@�/��P%��F��@�^�]~Z���|�AZ�SC����C=�U~�+�|�du߾h���j��3�����"g���.���o����j<ˈ�; ��l�W�+������j-���0J�7�]+~��
x8�����#R4T���h)�C�����6�X�W��2����vk}=��ގS@)i�cw��-$���<��,'{HG�&�͔�h^Pq�%�2�)��a��#-#�$*���Tl��qHvd�U]�l��HJ�u�圱�S���*I �x��.�`Y�y�L��\ĝ�w��L�i��ZoC��db�P/:&*\G�x�P��eYO��P�S��EAC�b&n�6:jʊ���fA}�?~(���g�uWhfat��[�5Sp�[���nSq;�iˣ"YH�b��\���9RN�y��;3̮S!��ڢk?�(�A�����2�he*������E�	�z����������q$��iN����Lj2��l%�s��3U����]3f�&�$��u�8���Tq��R/����'e-�Љ]C��`˂��4�����B.۶w�`Ϩ���)'�"S��oG��wRu�@1V
d��e�S
i��cK�L�x�ϔ�ʗ�Z���̺�J��D�=�/���n$�EJa$���"6v�����TQF�jL�oZ㐟��e���E��Թ���r�(u����~��Y�p?L�Ǚ4���-�1���DKƹE�L"
�I.�+�0�DX�O����A�1ѕ身��#O���� ���9~��V��2��RdfHl�9���Y�\jw ��I��{gR&���1��Fp�R��K��}Do�hw��u�ja���G�9���
Ტ�%���\��>a��1���\�+�`� �	��$��B*��i�s���yˏT/C�5�Ħ}��yΪ�a?���j<7�>
z�O��,848�B�F�"ۜ��R��q�9ng��`�(�Ec�5�����b�|��!���'t�!�py�7"����}<b��Ǳ�_����5���_	)M���
�pP;d
���UQl���L�'m �t�i*8��;'�vbUF�-�͟��6����0G�	ʊ\�����ٵ3=zH�6Q�9_�lg��\=5�����{�z��������#n�m���<�u��.{�̸�:��>�[���+�8�^�Ͼ��C;������5>:��B���X���u^��"����y����B�K���ʏQ%1�FVgFvac#t��^Qlu���u!�@G�"�8�ʶ⍼�(�Y�7ΏY"�1��5��SB��14B���UX7/�?�H�j�����'�=����� ���M�������F�O+@B��-R#�R��X����>� �Zn��y����	�A�M�Ed�%b�ݜd�q�3u��f���̿zg�\�03	ٳV�%�>�,�c��������	��zp*>f^��y�
��!W�i��d���K���@Qɬ'	�!�[�4��xҊ�i8�+D�'5Hunv��ؖn�OF`���&O�X��������&�IFH?�M�cvG[gᐴ��=)	i�6k��{��M������M��d�|�n�R�1���X"̺޸}9!�=�"|��_��eݶ�a����<l�%@��	���sQ�
����x��1��*�ko�<y��+�֟���]�'��о!��H9�X�(���LT��io~e���*�G5`$Ƌ��!�ό�!Ձ�P�+f���u���~˦~3J�W�r��h�{?F��f1��*ª;Y�
5�41�|Vf %���j\��B���G��)"(��r�7P�,��g�x����m�������fD?�R(X|L$�]!/���1������P�����UV�VW�F�+��\ZEFx��� ��w�S�v&׋SgB�@A�.��\)T�4�����K*y�,�X�`a��h��D����E$������OA���KC�Ϥ���L�a��O�����v�.��\����̖D��FG�b+��BzL���֒���v�QA�H���7�����+��,a���I��~z�_��%�8�j�Ӣ�[�n�0U�g`�
_�p3�l��)��XC���u�ۂ���h%�:��MS@2�V�<���h�+���el�'�L���,�i��4�C�Eh&��{�����jQA�|��#Y'B�I��T*�e�.�,Ѿ�K|U�RC�'7ΔY6�h:�|��]��YZ���:7��^��h;C*�m��+���%�Xf$�����	\r�}�ԧ��&��(�:����%e������ڠ��2|d݅�+q�%��hh��� e< ����iVhWɎ1kNN��L$`�S�5[8�_F��v)! �]P��\q#��%�6������	�:=�n4ڝ�����9�p#��ҥ�A:0Pq#�w�UA�9b�ї���Hah�hO�r�L`T��D[��C�ߩ�
�i(�!���L]�f��t�ba(g��>�H2���B���p�Z��(�f߬H������gf3q�3	JbuÃxb�� ҋTkNlY�`�%�S�e\���$?��.8FP�R��"T, �L��p�/oW@e!䥬��XS!+.��b`�2�S����x�^���nm���X+��a=��=����)��_M��r��:�z������3i�Ŭd�n& ^[["~��V>�2�XM'I�>�@�	�dc釼�l�*����rx/&h��R��p�ơ"��㸮_��*�8�C�u����um�_M�B!�@���X�eӋ�"��j�Q�*��9(U��^6	�����@ �=<�R�*��	9�>�&v޽l-sWT��/`;K/>
b�(��Y��т��<�1I+4pӱ	�٤�tE���@ʍ��c��;f=�^g��D����М�^�
C{3�NXv҂��z��tYª��j�+�|p���)��ͦ��yQƙ5�M�?��������a�c]s����M���>Ru�@�l�<v�O�$�R �"xCK�4��\ڶ�����,�M�@�!�Ѡ���k����r^����*�3��N��^�������͕0�M�"�����%�8�V[�����A���{�.Sr�;4k��U�kz�=����wG���F�+�R��wL���Q���EgCFMd$d��ꃕȍ4�M�"B>����o/����
df��\�'����F~>Ʊl�g�_X�J�2	�󖧐<�oA�?���K��ŀWў�X�w:�ǜ��G�.*3���I�dL�:nϜR���/������P�Xe��z}5�����k�$8?�����2�ɹG�|��T�7��,�Kvh��c��8������!�W��!�@G�D~�u
[�y���S��R�5���ѱ��E�-�p�|ڟn�\I.��gp��°�����8��n�����_n|0�����N?����y���.��v�eZ��C�eM)t��cw�Xd�_��n��`�Ol��7��i��drѐ��?���G�����:�Z�0�3Sp�& 	m:v�u�=����7�*��������oq6�â~5��Bhe'�}����F����ˬ)k�}��'cg�^J	F�o�޿D�J��AX"�o~�g���}#F��f6��� ��}]��'����J��qe�b��;��>9ȓ&�	��Zi�s��>Hwѐ�fڅЋ7~��O�^��g���YX�A#=���jZ��*B~�E�9<�<To��G�-?�ڢ��k�y�ޘ�_����p���k���A�с喙#C/+�Dg�zV��c
����]����<����mL=������F X��{x86l-,��Mwۇ����$������7���iu�a���_R�J�JA�P\�{7z���c}�w�D%l����Qy�q��"�:9�Qm�g�n���#wj{��Ɵk�l��o�G�s!'�B�ݝW�h�K��2���/f���&X�3��PCm��J|��#�SQ�{io�Jmoa�g��U/�*!�C���#�L��z��Qn4mU\*L�C�x�Gl-��+�����R���Bk)n�M		��G�/v�'ꍾW����e�Xv���]���
\w�����Bq�Zr�'A��u~QË����2�L`����!y��W�-�ܬ�1Q�:kU�V{w�,=6@mF�
u]]�&�������I�F�9' BC*�YB�s��J��]��L5ARn��8���Xl�+k�T���_>�����{0w����	�� ��=Fԕ�_Hf���M�U)h)���F4g��Ɂ�/����*(��Or7)�
�/I��i/ˊ���S���K0�cAg��<ȔE[��N�3�}��Sq"�@��柝�#C���'
��@
��63��p�Ԥy'�J�Ff�k�f� �w-�.�- ���+#��O���r>���o��m�踱]u؟^K�d�� d�SK#����4ZU�Re9M���Ԧ�5ꎤ���M�@��5��O��=5� =�����R_�/AQ�y z֍���16c��cg�I����kK����{yR�@,�]YD:�M����s� �jӶo����K�7k�1�8���5P+�L��>v�{�I�$R�:���UAe�ƒ�O�9)�����yyb���LX���x�m�s�}r�$�t��>0�J����8�^NSzp��;��h�GD�.�|��M��Ȣ�����5�'��u�],!����2�1Lכ�B��g�9٘��\Z���9�t���t�y���;ó���~<R�@F�}J25�wK�����%"<T����&![�t���6�J#$vW�g�l����rϊm�m�Բ@w��E֟A�Z(�ת7(�/�a�1|x�~X��S��?wڻ�Wר�� p<�񳧊nG83�������A2��呼!K,���m��)�K�6X����y2�*��t{�LG��ы#�L!Ԅ�;��:z�P�D~ֹ3�f�R ,3�<���t�%�@�S�o�d����iU�K�!]pե�R�(H��c�ֳ0 ��;g@u*��	Tgz�~��:��;g�F`�a��0�����q�ȅ+��P:zK{SbM��$傇�$`����9��|z�!�P�h5�w) �� ?�GD��\Bqm6������f/�,��AC�X8 ��]���2I���>�"��2����ZY>�­���_M��(�O�4� ��!���U�ͭU������t8��#S>@ݷ��m>x,��ƤQ�����j��\r�✷�9?��{�����C��g�s��K��V\jE���j�ֵH�P�[%g�K獷� ��UF��w k�UH\A�'��ЃJ��N,�'��:��O��/��������Q(�v]| �
dt]	+�ay��+��D�hq�u�Sk�J�:���Cv�x�>��e���_j��� ��aj'�I���")gCM��5U�� �l��ռ}Dd��b���c�>��<W#Cp��wZ��'^�U7
�^:8�1�|�@�H�����[V��.X�)U�Y~E���7�k��SE�up�XW��/F�"��s�vK�@�Q�{�E����оȸ�	/�2��Y�0��^
�E��th'��v�y���Y~Y��ʕ�)�m_#^�ٺi>���d3h�<�ñ.?�O<x�����k���zEСS��G�)�9�|�	��]��!s6 � s5�n噃�9L �3a΃�Ǧ�P�O���2��l42Ąĕ��SE$�~��m(��(8��*J\���P�m�%�A�%���a�@M@��ށ�I�;��HǡB����$�����
���4�)]��ǀ(��pT�����m��7y{��W����|�QM��`����A'�~���&�MB6�[��Uj� I��|�'�G�UN͉�2u8N�-��� s�($�9
#ʿ�y_*��,E�k�<ً?��L)?�Y��fj��/<\��P�|K�$��W�y�t#�_	I���V|�d���/���k�ր�Z�~瀑jÉJ�Zb����
���[#���%��5��|�ѷ�����\���v�2o���4�E�)���ȕk��l��)�A�)__H'��]ܸ���"%PT���*��\:�\��a��S�LT�2)�z������C�0 ���)$��stG�lc[Ϣkq��	���AM{J>������dC/O��9�Ѻ��%���?�p�t����1���SVM��T�(1 ��=��ߠ���w��-	�<$��Hg�2�q��>��g��V-�Bth"~�Ĩ)osn���dl��6Z�=5Q3@�иF����g�	0WE�y�T6����]���!���N�5H�-��{�����k����6?v4l���[� !�V�j�v��V�K� 7%�����U��3>|�^HS�!S��7����vK	�]his�2�� ����מ�L����^�&��}9Ty
�6�i�ikȘ�!gK#MPJ�GD�$'1d��4�Hu�h�2���Z��h��s�7�A�C�8e�D��dE�	/��󅻼�I=�0Ź�xu?����8�!����lk y���yE��ݸM���eϾ�ׄ��T�t};rln���G1M9�
b�_���3�+�o��{N��;s����Yؓ�����+����	|��>��Woۮ0�F.��.C=I��:`l�]���v��H�3����-���I�Ҭ��5��2��@��I�zqI<q�[�bf��ti�/���q뛛۷��<%�'2P �\F��9������H���7��<���d�0q!Q���&�_%j�q��Y9�
�#�
���rA��c����^���Ֆ>6�Oo�6F�`���=�P�6T�LP��H�����~f�L��se�$�p����t������4D��g'�w�2\0�GN�*��K�,A!e(a��*V�X��W��5D}�~�8�-���ޚ��[qD[l������Æ��Ğ������X�\�̅,t���)�4������u�E�)�G�����y����E#/Q�amŪ��uĂ���|���@�^D�ϻ~U�Q�x�h�(�v��nx�0�~�C����L����Z�V"��[�r<&��8=�J�;t�X�k����9�"�
۹]���� �4g]���_���b|M�ɶ �\_�G� �yqn�R����ɽ�`�������HH�sb4�6��7�	����~`����ynȂ����aL*�0z���k!�IfCA��o
MH��*u~CLm����±�h�t���.K�� �ݜ!���4lQ�}�GT$��ن΄��s��rdK�^X��G�T�lJ�(�렭X����5ݓ�_V	z�S�D��l׿�]]NQ�蝹�d��3����Q�!,b�^Je�Գ���� ��[X��c����:��E˚�፥+�w��l>[��Q��mJy�4��WFo�F�f���&zC@k9�kЁh-��7ӳp�8��
YSK�.�$}&���͊ٙ5�B���^zG��P���m���$L4W2���_M-�8L)����ѿ�=}����ȸ�7��T���K��<fW���'�t����(v�]�P8)}�RG��fB���kvҦ��f���'Ū�Փ�D_b��جgz?�d-��C��v}.nߙ�Pz��DH�9C͏��Tk��v/�_8���j�-/i�բ@?����A��6k ����m�b�^����<{�Md�
�͞�5J-0Dd>�?X�0L1_��b).(dﱘ|tw�{���	�����z��Q}O���r"h��6� �I&������S��!I�� �OщD�Ӷ���B��޻��
�}�~�6�عƺ�v����&�������Y��� ��t\����؝'�Rg�;�.%��f��]Cݲ�����m�N_*)�BV?&]}h����5@��x3��`sn+C, ��w�4�g0Q�����@�"���k⾚i�i=���@���,<���H��K���Zy�[ME��4���s���!��?�5��?d�\��E�n��VF_�O���P��ŉCj�� ]:��x��l,D3j��I#3T&�]6�!ġ�t0�N�n�xF�fd��gq!��-�D�7��q�1"����ih��  �,�6=QT �7y��X����J�����ɱ�u���Z���-�HG����)��?�X7�����9ي~
�L�GmdjHҹ���~�zUt^De3:�� q�?e�/h6ŊM1��{�U�"�G:��f�{h@w�S<�!1x}�V�	��G�����8��דD�+v�����٤`�Ǣ�P��t_r���{@MD��S��^���a3��+���_"*��(�kMWm�<2�sy9���!`��>�k�>s�@^�}��c�,�y#4+:�*�Ҵͭ���� Gc'n�if����_�]'ћM�q�6K{|X�p6��dV�>��t�l��0���Ў�hu"����,S\�Y�ez۝� T@K����%��݈����ѯ�i���l�v�?����Ǘ?�(a�*�(O*"7o�	a~N�i�o�K�p[���l�=��^o���^���/t�s�%�ך���4T�- Ǧ��=8�/�Y��-��^M��V]�����6r��j�o�E����kL]0����`�����3ߑ������t�M��^�	�&���Hʆ�X����=�O�j^��IB�O���o�7EF=���9���xU�/��I���=��b83M���1bFE����GB\:#��~1��MT�G[�rG�O)�ͪw�)Ż��u����q��Тt>�)��!=�׍������*ƣ2�>4oG���/�����[*)�����<d�j�l�0u�$I�����x�v��v�M��"��})����M��^ ���7����7q�&���\�ȝ�W�箘�#�Ϙ`7�����pӘ�K3�H�~��$@�$���ރ�ї�k�7���o�� ���Qrx�#��ԁ	.�x��\(#�'SŪZNBI$;����]7u.&�|y�$MO��y����>/����j�e��-�� G0��%���L\<@���B�*
\WQ��|�%lG�jr��_m��d��N��G��u��+�����l2 <����Q����6�qo%1�b�C#e��8INۣ��`�o�8oO�
"�W}L�>&{�C���8������&q*jC�v�gx�J�<�/F�Z���O�U~k������V����ۛo�uO��Ƨ)��ˋ���[�.��b_b9��ʸG6�Lk1W����7�M��g�#l��[\VV�(��^jG�$wkˑ~��lt�o��Jx?�E������+�K���rvRa_8_�Yۃ �N�%y�F;m����浴UVvm�u���l��^�q-����[(�9�d������fse���)���Ζr�ݡ4��F�O�b��<U��R�,:H�ʯߗ-�湺}�����dJ�&wl0>]�-���5]��/�Ev���>��k�KȈ?g2��nQ/f>���U�Ј��p0���{������>�GF��M�B(R�̧������m,����b�wV5JVi���7$���eR�Ds2�	CN-'?l��p;k��a���ɱgL���R�-_}�d9���������b���Q}�	�.Fxn��u���mܤ��4�"�i�(�� a=�������~ϫ�pt��F 8LrO���PMݢ}�X_}�B������q>���ߍ��J�k�@{���gc�_�Vu��6���*]��n�M�H��y�N3�AO�YP�y�����UF!�6h>�Ēsji#z�Lz�avul�G1�,���\Zu!�1<P�ͮiw}�r����.=o����3=��-;��&�{��L֫T�&� �_�m�5�� zd��ל��0�6e=�����$�z-�ӻ�I��a}����0�Z8Cb5���oG�35�H�9��KJcp<���z�hH��g��|��:k��M��Qut� ��ӛ�Q�ѓ^��HfZ_<��t\=Į5�Ԩ�H���Ц�����U���B������\�}UqQ��E+��:ǌR�ȕx�>��]vm�^�-�0�q_lι�������O�6����Xs�*$�������*�n���kt��F����o$U
�m#�C��e#��yWL٫��A $�vT2 [|HP�t�6��y;��q'C��B&w;��>k��F�W������v@��]1�E�,zVeQ�8����,�9p0?�۟b~��uH5�F:Cb��r�O��mB�����1���m:�gڷL}��/Ydy/ �nA��V�0	2���\ImJ=���1͞w�A�-�x��x��ꉈsE��4�����'&�H*mޞ����0*�w�-��ºM{_9�<���P-����h?�����ȳ�C�[��$�i)���۬�e0-�1�_;$�=*U$y�]�x+gUVw�fiBr[�y��u}y���n�/�>X"
Ӕ.,w�]�H'ϳaUV�}�!sx�=���@)'�]fJ�3L�@�=�~5���O��C��I�Iű��{M�-_(�(<�is�_R�{��[��#�+A	�44�t�8��F�����	��_��w5^��+�*��@�Pj�0+��*�Y�U^��ʒ��(k������z�QXW�K�1Yߪ�b�� xP�B1#xLH7dֳ���sk��rb��:��4TW�GW��/+�8Ƨ��2�&F�%��g�W}���6j�8�pƑ�Ees̈́x�B5Fy����Y�w��~��Aq�#���b��f��C�Q�L8l"xjw"U���{r�(�@�!p٠�B�����b�5�V�[_��\�������3n���+к���Ō�X�3/�I�鍔1���Ƥ}���zV��F@/iiʌ+�G*\�^�%a2�s!N�Ji9��i5��?e�G[�d���0DR��R|�\O-�1�J�}����F��%yj��S�Ք�G JTOò�y�9^�8b�+��/=�P�������b'�����>}Mz�<�y�������/BbG3���������
)�b�2�ӄ������o7��*eAJb�mp����([Us8t�-�O�43D���׾Xez�ژU/#�X��V�D�Bdj�>i�_'L�@Ƨ��Z�S���0u9,��v��y�5��2��9��3���7�U�U����J	�l��n�h��[a��%�xQ8��l�9yJ����Rړf̶Pt�}��-d��D��|���&�K���$��H��ҕ*+���Ŕ���CȢ��H�!�"�ǌ��>����yrjp���bX�c�	@���|�$���ZDe�d)�w��l�����-D{2;N<�7PK�̉���nK5� ԰:3=b:�;���Z�2zT��Q��t�����pF�����G�m�u��)Jm�
�i�M�qS~�A0�V��q����as�W��@W܆�\cu�N�f*�����,�6I���^Ufl�����6n�N��s�������7�!A���Z�H�Z�K� c�?��	��t�If��T��,P��|�w�o���舆��ud���k��V>惡����>�A����Q�wf�\��gR�5�P����<��gTD�;��������I���\�,e�����˗ �@bl�K'۴?�;��k(��q��ưZ�_:O���^�6��L?�t���s���6{��thOp���t
�[�©#�&�fr&7�F�>0��L���oQ��d�����$:��>v�p�3aN���$��0�Z�C�p���渤�xR����)ź�/C���kM�Jⵗ|�N�k�u��W1'�4��e�+����s���)�У�C�=�xGB,~ 7�O����v�m�َ��F%�H e�^a���[�^O ���6?V)�m�������J�Ne���i�nіT��{K���G�4��ΪOҶ愅���G*`�Z��f�*������� e�ܦr�uzf�����)�7�Z>��
c)�⚟��x_jV�Qz���['������B|�$���O���J�|��"�$:y�F+�~ے��jR�C�z�F+����箉;�d�a��"��=	"۽~����4���X�%�;@�2���IF�6Ah:n8��>`��wn��E4b��P�7E�����5	��hZAq�jpL����:'I��?���-���0�WhO���svO�6-��*�������P9ַ���=�j����s�k���e۪�?�¤���.e�^x�
���%��@����0�s���-��3��_�;}�M�7�O%��@{��T���:v�o�6�p�A��~jt�T����w�AȬ�m�)���ꯍ�3E;�xF�%�KG��Z��V�%}rA�ML(��!��S���f0P]��a���C�އ�e����Ԕc��{�����n�J�좯D����7X�^�@m<5���ɋ|�.*�?��s�d#zh���B�����%6���Ƈ ���.��8�r�0EzlB�td��MUi,Ե�B\K��~��e�FW��nK�{l���4�^����aƇf����G2�b�0�`�w� �����d��}|�XBp�7]v3��{��]���
\jIz�#l�P���H�����'�玲9�A;r�v�oș	�9�?��Lz�.ރ�@sCt�!Wb8���Pж��!�D�T��X0�̪��]�duZ��M��c���i�/�PT�9߈�<{S,^;o�H5���/���	n?���@�*8�0<pW^!������M�j�xi�~s_��M�q\Ռr0�b�w�8U��%�^�`#eu�D�^[z��u�j��������ae���3�c��KF>�v*<��g'aCjP�~��&�����&K�n�_>C�e4��"�8�3C:ʰ�f�x��x{�H1l�.���D��?�=�ΐHb.�CN��辆�d�`��Ū2��.��U����}5
�E�l�D`6wU�m���J_��?��;?De�y�|F�O����-�X�O}��|s��ދ�A������&��������M{#�(T���t�r�.�J6>��'q�7��]�"��+��sԞ��	T;�.˛څ��@\�m;��Sr��Y����Y��9�i������v�O�Q4{#�ז�׽ �t���J�
N_��lج��M<��g4s�O�r/�iN�p`�V:��H� ��w^<}��WВ�s�KY��$/����7�
 0"�&��Bn�n�m4��ڡ���t�l!`Я�1(�)�[��%������<�H
3�T3! ���a�m��~-f�Tw44�@�_�����ߜ�L�%Q�pF�*��[ft��7oT���y���Q�!�o߃-L_ ��[��Y�5�.�B��v "�H4ìo[�~swh�aH���"���7p��HN��qq����K��{��ɝǽ�A��#�������v����+��A�-J�G����2L�qΚ3Ȁ_h\�j_��ف�z�i��?;t��_{���k����!�}(���Wk�ݏ*�-*�\F.Plliq�&�,���<��W��B�uk/P	xx��6!9pl֑����*�ْ��m��(�]#�%����� �fW{OO����d��nR����D�?ݑ�5����[=	����}2�LC�T`�_pq'���֋�r�\���D��OZ1��R�ZM�c�Bi:ށ��
K	�gm�bw��� b��+O?�� ֌�N�O���;m�w�Q��8 -{����O3_ϰ%-�4-�fq�7��!��n�����Qz� �v�;t�Mf���F��s禗{���~^,K5	Q;1���K�q#Ű	o�"���o�v,3�RYe = (0��F�D�����qAp�
�~%��� sH�t��1����Gͪ�;��$�f�1����Rn$pZ�� DHQ�u��DnȄE^���3���wv�������Be���Ws�4��R{n���;��&X:��I@$����Hl�!��mѐ��ڲ70�(���C����Z*w�)�6�ǽis�"��CB��9�'�#w'X��!��$���i����;��$5��K�f�n�ֿ�9�y&_�+\����س�Y7�C��/&��&^�v89J�W�o3�h1��!+z���#Hr��<��3�g//s��/�������\��r�yW���|\�L�s���4T�o��;f�v�-��E9\��G����J7�Vy����Р�������Mg�Vje`"��n~�V����[�<'���d�ڴ�f���*�E��$�Y���j��F�"�kPY�~�
!؜�C��B��)�bYd�!-�T�!�z���.	,8;�$�c�y�hk��(��}ySVp��62�_���ʽ�n6�ؕ�� �nk�5��Rz�iI���U.R�"���a��}�Ns�x�ฅ�c�Z������oFV����zU!�xH�/�S��χ���0��a�s2��@c�At�z�t��;%��������ۭd㆙iAMpT���k�%5� �qvS�k��7I�ܽ��D>�m�M�k�tܻ>)]1��S觴�!���g?F�QT�`|2�Ƣ\O,�I� ���������[ExH'G�6[���}xB��+ eN�"ڶf��,�b����a;�r5�o�b{.���e��/�0�Hsk�Ò7
LFZ�[}\d��m �����D�� �Ix�i��T�V����8~���^��e��"�5���'>���l���X
}� ��mUm���x(���L�zUT���p��S۸"��F��:Ks%B(wc?�����Êqn0CW\���lό�&�p�? �K�3nلr6�n��W�a����-t�������fyt�m�s��{�#�7���������yPV�mVaϻ �N~��x0�j�I�u�L�
 ����	}^��0?���"�7���o?ເ[�(�����?�p�M���Š��`wL(���x���o��@A�@4!,��W�!�]�"����gU��Qk��M܌�x~�J<�6vFy�ی��C� ��3-i]����!���B�֯^$����� �2���_'z��-'� ��)X��Ͳ��0������+1�[S���S�����MbPY�L#�b���h���/IR��������U�L�z ���9������^<�F�n�X1Ew$���|�0�8�׬q�`���ړ�"�S�6E�؆��L\��|Ӏ����=�U��"Bd�(w��G;��=�%��<$jTeTĀ�w�2�v��G���E(��s�q�4$wZ��+9�4��B[�w��VH�ٸ�x3Z}9`[���Q�^ż���iR������w�粫f������p^����ۣ�7��0d?�=�j�I" 7�M���#�� �B1�/K��hi�5�����*���<�^ъvӣ�<Ҵ]{�i��&����5�܎�.s��oʄ�O��RK��rX|F�Y��7�=�?@����79��
�-�xS��s�H�⚰������scz�>�Y{(h%k�&�
���ླ�	�Ai�Ƹ���I_ݐ2����A7��e�U]V��|��K�h���%c�&I���Ef˾HD3�a��gm2���^i�j5~��g��ךz�ތ��yV
���ū�&E��f�؏j��p("ܱ�k��ڊ><�YN�س��,N���2x� t<X��5r���vhh��!V��������Vӂ�Z���e��1d��m��P~��&@_��G�>�isW�U_�v��C��R���j�����<�OG����Gfj�m�����RR��;����9y��Q6��1�[n��� �l�����c�R�6M#��"�S1�p�]�o�_9#�e���(��a�[�&F���ۇ>�;���Mk�eI�T"���O_�@I�$�l�v�I��Z��m#��f�Kㅒ(c[IbO� �A�q�����)�k�z��\Vg��Y�ʃ>�,M��a%��V���Ἔ`�1�r,e�1�`�Q�|����q��BV���G�]��l��HrSw}��C5��P�� �<}Z���t�"� 0qW�P�%ty�;��|h����4�lN�1B�	�P�#�$��??���֢#��n�}���M*yi̲�m_��Tp]ᨍ��s7p����>I�	F�k��Й=�ԉ��`����]�®v�x�Z��}�tg���m�v���*�@}祚�ǚ�	B4���,+�'u�	���Bp,�c@��L�+�V7A�/c�{�GF��'5A�5��ڿ9�Wˌ1v��q�L4��	��c�&����8���k�N0!ϡAh�/��~<�|i#�b�Ar8|���څ`p�����0��"�Ƥ��h��-������	��l�gW�V��I��mB)���q��Y��h�����y��xh�PpQ�0�"� ���I��8d�Ю�V8�Ҕxm�B�R~���MW�����N�2�\���ȗ�L���t<�6c��6�Y!;s
�x��K�Lîk"��D�Q�����`@�p1K�Al�޸\7P�$��!K�`I6pQKi3R��9̵`�����r=��� ��5A9k4τ��ƨX=�Z�)��xf�ߖB���[����i�	l���T�����y�'����R����#!�֞��s5%�M�)o��AWp ����%����B�k��X���K�F�mU����*!Mjct��Z7�Qbq�,�p~d�D^��<��=}v�&�����N���^_��0�T�r/)5]叾�[�˹�<�$���5y�>�� ڞJ�u2"�(j�٤yjL�*�qEڤ?�M+M�9�-���?�W�~��h��[�A�z�^)1��,��y�RKmK���`�̐�*B0N�ۼ��6�9�O�-�����W�����ԓx-�����:��$�S��Њ[�,��Nw�O`�^+z5�pߓ�*7s�6������m�|�
T%g�`�������9�.b�?���ܤ@.z4��7�#ܶͦ�q��N�w^�(��$47q�BRm�׸F�+\BӅ �Q՘Yx�����W�:�\͝��xϢ���O/)�|��^�ܣ8G��5�n̷ؐ����!Z����걎Б=�ښNaF�7%ͦ�L���RX�Zz�D�!i�B�#�Zӄ�}���
����Z(�",�v'��75b �M9��TXv_ҥhɽes���|���O�[}*�O^Hlc���ëb�?A^	1#܇"F�՛�����A�t�ۙS\sY�����3����.}����W@��ݠK�>�<���@��]�u�p  |w@�y?�{�!�!�9V��Os��j�-jBt��g�[��jT3�f�Պ�H�;q/>^��a�s�69g�H,�'�g�5��W���|2I|��1�ͯ=��v��Ǽ^�v�6_�n�Æ8��%z<��i�1&���8��#,�Tcm|�w6���5��®~/a9�� K�����D�OpN	��SdϳpD��p)=��@�ѭ�T���fS��	a��^�LA6�n j��5��Z�͟D�}؟��л�b��!o,QR3�l#*�Z:�H>
����!�ld	"8���bDm��a������q!�����٤x?�D��[����c�G�y��)�m�t�Ă��E�e���?�BV�QQ�Z��~B>d8~7�;+D��Tr�p�+O]��fC񬃒zL�n� ����qd.��,�����,���,�R��iΤq�
"�䉍7��G}�1�#������|�"�Pya�P�6FҶ�S�b����A����݌h^;8��]�����
_k>"�
�$��zs+��.Wcm����N-|�^U��`v8�.v��#n�ε`�k����.8�Gd�r<�����d7 �G���li�^���a_n��B��A/2��.٥��p���&�����g[��7����d}��x�h��C&΄��C�1�8��܍���1p�t�
s0�^9Y�ŽZ�����������3�ϙSn��%��Ám� ës��lB2��k���?��WӃ�[� ���3�����,�Ey�.m%~7���c6��S��gX���<B	�����7	�t��Ua�_������t�:�ޟ�����f������ܼ�u�B 9 0�a�%10��@z�j2�ϫ�ۿ �0�O �*�ߣ]�|�y_N�\���O��`�~�N� zP�;�������wfAHo�m;6�2L&�<�]�"x���?]�m�!�>�v�����V��8�+�Ps�+1\�27B&��[F���.��h���
tg��:���L�ɿ���W ��8��HP�,9#���E��総y�5J�� ƀ@$�d���������ѱf�������i�bV��4���]�'�!.�s��xc`@]S(/=yƚ��Ǉ���h���Vu��Z�F���J�֦c+��@?�29Ţ.�@�Ȥ��A�F�6�Sp&�H�cӭ�雫�	1��R�ΐ���	Γ���»6��>`�2v�S��m���� D��d�Bo����W��-؅L	�u�n�{őS	�db	�:�������6�z��K��z��A*�����+7@}��Pt�xK/��,�yW*��͟h��P^��a�BUj��GO��p�� ��[i��U�$�eLgR~�fjÖ�-�l�I�!����c�W�{'3h��Ѻ��{:1��!�ri�fX�Ԙ�/�N��M�ݚ��2����d�ФfD���f�T�2(�W��#�~l�+.�.���{�a�+>�6[k��eHu��93��x�}�X"n�F5l�C��3��MN�X�
/�/:��jEP���Ҭ7О�4�6=���c�J���2��k�tO��-G���WK�l�ڪG��R��V�WF���:� �-o�!IX���P�R��%d��[�Rq���Z�F�1Z�_�s=r0���ٵ����0���e��t��e�����A0;�;�����9�^�$����چ���1ы��:Q�(����/P�i^ْ����[�VҚ�ԭee~�x����M�#�\N���Vh;�#�]�Y�G�锾�j ��ls��q��~��uhЬ�ϑ*O���EF<ʋ���GB4��4�j��WB�������D1G�Z7�K�LS�\���.%:���U�S �w˨2Q3��m���k�#E4���z������0R������x;�l�(7V�3fS�����d\�a�� &~�gW�!���
�%Ul�[��7^&�¿���P7�*����0��D�>�3��G�=f�P�:�[�F!�5�Ԙ"m'z��_�;�B��r��3Ԇfp�B��O 7���GR.D6���W_ O��B�4S����M,�"�Ӧ(�k;QʞP�ό`��c��yc�[�D�"�u��=�Zڙc�t/f9��Q��<ί��v֧�����J��ž3��]�,�kyox���]0�F��DM�d��-hC.l���u�Zֲ���o���MH]��H�t�J��cj�����x4�E+'!X��+'ĴUP�Ab��<-j��(EgVK�kX*mL����@.�D�w�����v'领�!�%��o�5��1��_/#P��yBy���/����Z��c��/�������C-����,�eK�0��-Z����xĠ}�G,�!�����K/��	��+�g�E&�nvGbw�;�+Q]�p��T9��Xa'[��*��-pm=�����������7���]��~�1�����T����r��RJ\L�鿸.0[�����D�������.%~_J��ICuΎ5�Rh��'�Ûr�4��� Y�d]�D�4�y�֋�R8|�/��������ؒ������8Ur`�<���W���TI�zO�#ut_ES
�W{�"�Z&B�=�~RE�b&yy��汞���X\'u��8��A�/ι��o�=n�HDh+.���3����hV�L��X��l$Bv8?����N&,Z�YFWC���;���\�v(N�a����9�	HGg��W��P\���O��{�RH��EN}�ũUS:�h��J\<��R��Ԩ$jT�k嶝����4`�=,b��l�:�w6�Y����P��e���	�j��D�u*W����ӹ���6����dE".Ϣ��f7��/��.�C��Y\�����FG����8�I��|�r�kT��cv��e�[*C/b���sCo0�B�έ��E�[5��R��a#��k%���)�L�vX6`j�h@�e��H��c���Np嵿��K1%)�W9JZ�C��خa��v��^@,�,��-��C�rn���nw�S����3��{1�SN&G-��g�����y�t��ONO�y�Ykm�X�SP���+���	ݛ���W���'�A� 4Ia}24oQ��Y����X��~���rT85���>J����b�$����4�Ɯ�eg�r�P�����*���*��H7��6u�*����<�~@�1<3;j�^Z���!~�NMM2����O:g�}�"��;	LJ/�r�zHA�*9��d\r�j0�SJ(���%�C{7�
c8,�W��C��~\���k��i�,���D��
7 4c\1�oKͩ��
Kh��.�S�q���B4�`ե/@��� �{Rsl��r�z�ǘ�s!������k����O�`
1J���V�:c���xh���'N�S�@���l+�q.�6���	�7&�Sc�0)	�>)��I�P�J���l��\p�Ń�r� @ ��1mFn�E��ը���?���K;��Hþ~vm�YPr��8�"�����e�QT�b�|hw��qA��B����k��Ǹ�*���.*�#C��y]�b�c�x6�a^�����3q���$�pޑ���M��cڴ`��i,T�A�4�TN��P�ȱk?��C�piS�NZ�l��Ԭq�d���w�N���P�k����;~9�8j�s޹�(ݾ}f�7/J��)�����pcF`9V�aD7��7�{�(Z�Yјvi����Ƒ�H`�-��	.AT�>�����]���Z�7<��
�^��B�pQW5���ä�?��*���I
��N��3|1g�S��x�ⳏH�ٿF\�W�AK�����i}SPs��h��fK׋�Z�z���ה���q-��=��]�+�`���&9�����P��_�J�'q��a4�-�2�+ȼ���J��(p��E�͔�/8�\^qU�p�V4�d�������{�C��X�[�71�|q�PYA����#Xv�AI�#%�Ϸ��!�?<�,#���
~�zA�  ���M�׷�:�q��z�eȜj�B�2rߪ�©[�8:��*��ag�u�6b���%��/wE?P�H����[$o_z��Xx��q]�x@�� ,��4��W���:�=#��i�h��h
��X��T�N
��U�	TҦ��j�{5`.��k�^ބZ܇����{�\�[%w�+L8�EKB�+,�ce�:���ͨ=��тFxX޷����o�\=���Ǧ����>�D.��`�Uʂ���a�Xb�<I��l�u��v[���0�R�8W>�g��B-A;C;`�C�Ɋ�/�5��\0gt��6��,`��������׷��2�9�*�(�綬��>0�'G��[�E@�V�.��2^�η-�-]Ɋ�E���)"q��%܈ղ�6��Oڪ���"���L�� ��B�\j�&�K���JJ��ʒ�/)�������A��_��FT ��z��������[�X�	̏��i5jS�a�d����q��7x:�&Σ�	�����7$��+L8�9W ���h}�~m|yS�N����%=�7��?6qlo���Έ\�rdy��<�ﭲ���o��ҷY4~�\�ZD�u[�^�HfP�
�i]�*�X����WМ�n?}e$$�ڸ���k�Y��2<jO�b� h��	�J<B�!N=:�Ӷa��7�Q~�yayR1�
{<��'�T��n�v���,M�r0�63 �b �����Ŧ�tZ߭[����|��P�4�X�CV��JK��������%sl����ܫ+��CVqΥ�1�Z̮q�0���j:#6S��ʲ������9?�OL�'���L�o���e� ��Κīh�a������D���
��'Z�p����x%�>��ל��,��K�ʦ��n,�t$���+?�d0�'�!�S[g��;-���,iH��\��#T2������|B�������OR�t�v�X-�t���N�c��X~w�o�uq��:��q%�jq�;̮6����N�1�W�m*��?Ҥng��.oig;*����y����Pw/�>iz-��a�@�e>3�T�1�^H��5�=�mN@FF�F���rT�	%��:]Ba��#U�@��v5��Mu�W�� X���`_{�f���8ТrG�*�<��@G7`�%��[�u�u^�f�g]��.
�����ju�u�&�:��J��l���;j�W�h��'9<8ߌ�Z7du����1)�1B���5l0�NUr����~N��NH ��, ���UENA�"��^��NC�� ���z�c��ش�^�kG�.�d�؛��P�R�wN��aL}�⤳�ƀF��rY��o
�s�Hdg���\�j�b�[P/z�<t�]��2R\��v��@꣬�M5ׁ�P�6�zv�:�ף��A/yM�S�t�藿(xJ.������G������{$�z����i�`j�|�/�%-����흡�;YO�4���NU�,���jc{:I�8�?���]��޺��>�;N6��g� ������4>M�`�{5 7�8�l���+�ԫ�fo⟲����Z�VNG��d���5��ɯ�����^M�z��q;#�HWYzm/�>G�M��~�\��!��2�O�/y+s+�F� 1,�X����º\��e a�˷Kн:�9���ʟ�
R����fN���ux��֢���
�?�j�Ǐ���{���M��u�MS���i6������CjZ\��3��`���P�Y���0<�FY9�4���
t���oĕ��qv���EkP��"{|��Éɋ�F��wNg��K-F�{�)>�����y�ǒr�#	�sĤ���:{��.���n��u�q9=�B�j.^�FNyԙ6�����Q3G���.�n=�@��{�4_���j�9��q�I����P%NNgy�U ]�Z�xiI󤐱�4t�Ш4L*��	�כd�Р��3|�Y��X��2m��ʭz�1zԃ㫍������� ¨IV84����yj���&��RApmB��b��H`�bԤ�ejw!��Ө�a�u���Ǩ��u�% �: ���fݩߟl��g��Ϥ��0����1�W�uj}��'�����_�3�uiͪ�[C(�O�$Sl^b����?i9ˮ'�".�&.z�v^�Uu�_�4
$��}�m{t�i��%a������M�ʯ�I;�f\��#kN�F�f�!�cdM(g�W�ߴ�����s�r��
7[��i��7"��a��r�I�����=�O�62Oy�g��185w�Q���b�m�O������7[ks�+��'�H��hé<>;�i�U���E������Ի���r(?�����Ķ,]�[��OF;��I�;�5���U��_�
�B8��l+4��XId�צ�ͤ���kMSl=)�T�� ��ΰ�����#RX�x���{�;G8�xH��RƊ(=X�1n��Č���O�l|��a~����D߹d�JƇ���J:6�-'�M�u2��q�O��_v� j�	+�?���l4��=���!8Z��I���m-�#O��W�V�q)#�l��^��,�:gYxADY����!��[��OM[��\���{�W&M��n�-e�R±Ƹ�s�t��_^"@+p�����\{n}a2	� ��:N�#�!��Z�Na�!�<���&�j��o	���CVt[�`����_�f[����m�7��,m�/���ǟh�%��H~��J�]3�������j�5�l`��>}Y�2����i�O8A�8u���N�m�k��^[x�e ��W��H*`�ZG�����8���(k��i�+ZX��;�a��:�W+�X.dttԜG��H�F���Ȗ�>%�#�/U"�	(����Z�a˕���]������:��(�WK��O�x�v��;s�����Ƙ.�s+V{�?9�SDޜ"uYw�Ɉ�ԙ )�Kau���@�
�KW�"��52����&�����`Df������!jE����=X�^��h�Ƅ�5}��W��c�i�^ޛ�'�w�Ւ�e�ы�	�
6��~��mQ$�]���<#�cU�����\�g���1�t�ihK��n�&4���g������)}��,���k�w{��l������&��N��1yviKQ�l�bM����m���}��+!�S��j!����p�|��$�;���3�����1CM�'����������em�D��E�I�׊��Z��Ե�H6G��!!���'�޴�d�(���-�����mqzmj
|�YZ�ȷ����[f{fZt"�+5� £"/����_��E-�;!-�:�<��	XI�3�-pA"�w�5t�d�(�Hr����N2E=�u]��_�F�o��p�?#�=�͎o�lo��W�-"?�����o�)��o��/4)lG���\�?�ȵ&�X{T�Do��z��F�:����^��wf���H�����$�/gP줓��%�7�t];l�����/1w�����_z��<D0���Fj��o�5�[B����)"=����)�,^��s��ν�z'Y�$c�ɏ�݊R=���,hzR���[�<���d{�BL�g撏�o
o�ӝ���un���\|��7W����(-	�Q�X��_�ND7��RR����6�M/u0)�Ϣc-m��4fr5Rvବw��~h�J�આ��X�?���T�A�_ޱ�����2����?xj��!����e��zb����da�aK����� ���@�Wj;�Ǖ�'/S���ig��~���g�H:[��G3�?
��&�*JFmI�Wk 
`W���

�b>����B�d�	��N�{���oE�Ķ�Ң���0��Q��}��M��0���"
�!�E߮������m�ϣ��Vzc��9ꚃ����g7�gZ��ߖ�ŝ�,f��O��-���'�]��y������~9�����/,�Ų�iv�W@�M_�X8�8l�]-I&sb�&�j/�	_��T���{񅾆����Qײ����$$�N?�'g
���夊�X���l���s���sn��Z>����q�J�Dʐ^8�@L�9��C�k,ir2��I�e���*T�k����PgO_���B}�G��a|{���QW�O�H��h����QEP3��M���G�y�0S���կ���<��|9b��A�g-�Y� o`��͗��Ov=#�T&Xc*:��yܵ{x�6��W�X�̓:�+�P�Z�Ŵ�|��gR�DpI���B�aoNI`�:aI[e��n�QK4�b�[`Q��f�x��1��Gе	B$^w��r	k�n���,���Tam��V�:�d|�؀���p`����3�!�����J#��/3]��@��k�DJn���th @B�U#:�������LÝb���{��8_��+em�uo����&'��e�쫈h/�d"�ׯ&������;n��hjd����M�o40�~]���$��:q����`�Tm�Q�~��if��HDҶ��a�h��~Ir�"�N��۝U+S�/H? �+y�M�M2wԙ�W�_Z��Go�N��m����|�j��.��r�b���8KH�N����!�K�i�+M������)۱3.u$�D��!��+a��Y2X�0��-��ؿ����9v��Hǈx�B����*fؗP{m��u�e�O�_�����J���Ӱk�쨍�7FZ��f�������t!���h�*R�����z��x{Y,��_�!���f�{�$A�zs���Ѥ'⇞!M��"��(	�!����f����oXT �o7�Xg�V̶�H��=�b��6䓊k�*E,`/I��AH�z�+�涜����>���ʘ�U�1��J?�:W���xB��wez@�g���f$�s�%7mYJ�Ig�sN� ��i�Q�l���i�~��|ol��F0�t�rҚ��c}	-
�}����a�S���[,��x����>v�DGh�y>;}�cw�~6��#(��c>��6��%��F�H)n�B�����^qޡ�`tL�|b�K<F[���O���j��
��<r����X���l-}Y�����S��S�5l{#��Mx��}nV�:��B���G�P�om��ך�g��3ڦ�pMB1>�a�[�t��s�t�v��9�zz�~ U��XT�D�:���P]цu�a����������x)J�5m�u��Uj��.�y�>�aQ�R%:j�&�ڈk��`�F1ݏ��c�oL�U��V΁�/����6��e>ݑ>"�Eˉ��.P����y,C'oS�s�4JtI9ln
G�M��ߔ�WmSG���L����I�u:é2f�~Y�!��C��2D�~c�hZSi�#��\*�w�G��%�>Ui�K���ڤ�n6��`����U�w��RQ���3��c���xF�tgM��m}���ΐ��9?��ʨ��������ڂ"%�s4@|�L:Ȍ��	��߱���t����HG�\�a��+��W;ۄzG��;�}�1l�x�s4�w+l�x� �R�;*VS�'���	�H�ؿgVtk.hl�v܇��^�[V�����L6Q}�����afĭ�a�10�/�&�\��i�S)�{0TC�rGuч�#��\
�<�~3��=�u/ɕ�yP=��{�.�:�-� d;�g#��"���^�2eH+iX���`U0�.`��4@�0���c��+j,����WN �-��,�zfVFD�|S���|X:���O������"CX���Y9��qU"�[�xzBͩձ�r7��BlM��2k�aa��5���<��d�+
�a�(z���AXe�{j��3YG.��#���0�^;�~E�AHl�Ʒ*X�mj@�{D�?�0[;��
�2%��:��T��hu\��<�U���������S����-���m�����'�΅��C��X͌#�D))l��U���{��d�)WK|\�;����A���<v�]���o�T��JE)�����i5�ZE���>����u>E�Q�҈[�_���^u���^kX�OD�h�ӹ4�:�nI7�*�bƆ��K����i��V��l�.��yC1F�"No��+p�K�+���ip�>�Wʃ��B�e�74{�qvێ{5Ⴛ��9�Q�g	)Ap�2]y8��t�q�F��L�gϦ�W�q1���eK��Ŀ9[x���f�ڄ����Q�DW�Z������Z0�0����Y�mŅ�/:
:��@8����PA
l���sGC�~u��a����.ӱK�4�Pa�Y�r��'����e�u3��{qE�$Mq��K$R�T,�OP"�Zɡfu8v�����<��/�w͜&�N��4
�� ����i
�^.~���n���F������R�<v�"�DS���X+������%c9��,�=�ӽ�ޟ~ѯ�l�^�oṠ܀��͡��j�d!�M��]��Б���L�� JK�n���|z�ޢg�dp��)�u��S	��%7��I,��~d�4�r��$�g}R�A:V�t�+�.6w%��[|P=�Պȇ�X�^�9��:@?*�^�&I�ۥ�X��3픝ݸ'i���"��2kɴ՘�_ �}��)�Ђ��as���~���',��%ɭ_�(\a�҆��Ƹ�N�<�vs�I�;��=q�RN��kuN��*�4��ҹyY
�7��>&x����r��Z/;j�<*���\ï�B�
���W��1-焬bri�&|Rja.�ʵ,��_hO ���>��P6�s1F��IHvh������c=p?�(�#�A��f <�i�߃��0�p���{��Y�z� ��5+Ֆ�R��d�8��J��*+���X�[��Zhb94�va	\���N��a&��-TUYe�a�[�c�&��]�JXϤv���(�����ț����m�j@d����᭤��\�O�Q��fo�Y1�=.�'+=�u28g�~��1�,�N`��FQ�[/���aH���9�[>�B�{�xQ���T4�v>Q͹P���J��0��[������2�:������㒱|ۤ����W��ҙq��Q;^k�T�\� ,_0�Na��ֺ@�#�)�E�¹Պ
5���D{��ǘ����w�����{���}��<��� ��~�ΟLE�?UD���beI�}�pj'桛���<B�?������g%5a����<��rv 3y?�9F``��; �X�/B�{�����x�@��F���o� n�.�$�UU_�+�/�jRe.�������|��S+��z�n�������� Q�:���8eȍ������%��ˈ�����@o���31<�DH�9!�!%�L�@52j�)H���k�g���qܔ7r��@�g�e��zN�7�3�
�~��Z�L_�D�y)��G����ɕx�R#3���;4�bgs�����b�8�雴��73(�c3XJ�H%�
�S5�8�k��Hq� <C�!bW��u�#`�\�Y�! 0�	�z� +���0��XD��n���@;)
������f�
fi�Jcfm�Y�W݈�s'��Cn}{k���u.����Ի���%8�G��n����1{���)�x�KY���_װx��x)���� ��@���xA*-+�7ak`�:�<s�i��`S&����LY([��cp����"G�}FCd}�����S���.�=1�:N[�)OkU�O�"�>�K�|f�,f5�8¿6�hE�>�d��/��@��/|5[���|;�'
���jw(�ce�n�B��[���{�H��-\� �L�Q��~�H�(%��`9[�i��č��M��R;welC^#�M\W���>cK���k�Y�� ���A������?��`̳|us'��疦V�b�+�e�'"�C����%��q{6 @	M���iQ��D[�a�\\�ΐ��/^t>= �����VRpW�j@�9�,�m�%f'<�%}B߈c/j���
 �`�4�)I����^�"6�O�d���1��5ʩz�)D,<�8��@#Qr��L��S4)Y�Ԕ�5�*�E���_���2׍��/��G�x�%�z.���5S���\�*b�=���Xм7��Y�2�7�d�T6l���#��ٜ�]�D���\��ج�CZ�u�e<m������YZ���ޟ (`+�퐬%B��O��jwЬ�A�kK{^�m�W��I#!�$�p�5%��J� ��!�&1���q�����*�aT�'��ug����l��b�F�N��Ý2��Y�����d-�t���Z�y�Fwŗ�e�1��֔o$S{T��F���/Hz��~9���o�nI:`��X�_�ESq�TS�Q����s��S���UH��E��w��4g��F�p���@�.�e��
{�9���6��A�/��D��b<)���ݟ|����4��E�A�Hb���:��W*=�k>�r�E�JS ��5��5t$���cX��_�_κ�:}�O�7\��!��`D����Q���1�%�� ���B_�Ts��%�VY:�粒*������<uR4�+���i�c��u�����И�����m;Q��p��:�"l�=tR��og�ŗ�N&-	$qU�Z�(�ܪ��`��9?;.\�ϩ��:���w�'�=�xA�_�׋�
h�0�ޭ���jd`�'���T�n ��.r�$e�W���rK��_��у��vn���f� ��:��_ۘ%>ry�3T_�C��d2q����� ��;���u>��:g��zr��Yz��٣\��g�%A��.��o���Rn)�R�V�����@��������-'��pb6�
��7�L^��ۣ���(o�Te%h[��AvJ�i�P(J*�]4Z4�=Ay����)�6��T���-<�F~����ʩ�2"+�d�X�껻}����mT�Tx����靝u@Tt	��=�>G`2_�'Z�n(Y(�͉�iu��F���ٛ�p�����/	ְ7� (�����VF�����p��  �g��� ��:��V����i�}D��yp_m�DGz4�)�i���������؁2�T��m;�LBn!�?�06�6XZ�l���ױ s:p<Jk�HC�B�e'}*��n�g��`'d����_��P/�bPEl,�����E���2�D�� ��$��,Nf�5a���T|�1��qXm�X�3*
g��cIɢ��L �P^�;�)evE�����qv�Ӟ`���1��R�r�XqA�d?C6�t������c}�t���a�����)�o�s�����R3�����1����7
�Na��o���Sj�D*��p��^����u�� x"��������LS�wQ�����^S�J)��GFH�]�h�I�BʄX�>
��W��,p��'u���p��ܯe%$oAg@ɱ�*R�W�Eq4��u�O���ғ��P"��ؙ�_�J�*j Ț�o��ѫ,��J:z=ljV����=����Ycf��}���6-���zg�N����Vn�����%�|b�%0�����|�=�#��[ӱY�뇝َ��Z���\Κ�� ����lEЅCS�nE�c��b��|V����Й�̢;��wg]E}��0g�)f�G�Z3�n�t��U?߽I�v3Ƭ	��EO�MG���ِ�R��������lbDœ�b���;|�|����dK�N�	J:>'�����)��{�7��f%BZ�j�^�L1 ��v�b�Zv�Z�h�g���ݤ�r�4;��&��,�x�r�f�)I��E�=���sݸKSe���ϕ������dd�?��7|^���Z�!hq��
2�Rv[���,��Kq{�g�	o�tr�V� k�+k�_���$O� b�����|߷-�|�r��kX�<C��WVhn&
eb�����Q|f�����_���r���[\"z��h�?��=m��D�l�V-]`��NoA�Lq����:�W��>��,�Ϡ�i(�#�b������h�ප���)�v�{��k��19�%�[�"�MMW#A�`x����V!%�H�k���y��H�t�ܚ�]ޠ�=r�.������л��BE1��ߖ&��h|X����7c���g�_<)����z�!0�m�������)ʖ��Y�ieG�T���5�?�s��*�by�" 2Z�s� ���~��9s�YQ�oU�`�<>�O׹z����NC��rq��AU6�c��+8�9a��=�E�Y�� h�&@�C=	tn��7���AGK��ܘ�-7`0�76 �,����s L����2�S�׋X�Ǘ7�bl����d/��x+�ӹ�j�K�H��0E��T�!?H�$;1a���c�W��9�c�j|����L���z���;r���2��aɜ0��q�~��^���	`��sJ�D����;�a�,k��sy�����r�Bn ���ꀴ�M�f.I�d��_�����E4��-.l�
�!ors�膾v���w:-��'>�Ç&iq�g�<���^��C�m)�������k���tv�~�N���<�[����~�I�LDJ�@���pl�7*J�\y��}�����D�s
�Pg)djn�$�����a����Q8��P���:��6�{�g/@� ��H^}|��س۔.BQ��Bf�o	����sʄ�YFY�x|\:�������^rTNs�T��p���L��sW�X50-��`)#��$h�D�iXs�����{�I̤q&I�?G`f|�Z��SeJ06����u]�C+Z�^͊ŉ������"@l�h<�>��ϼ��Q����(�KQ�ᕸ�1� ����X"�װ�`6�+R��E@h���/y�����6����r��bE��8h\��B�u�J�?�b9�zu	i~ss�������r'՚l�Nܕ4u>�|�\I*e�?z�����S:G̀`"X�2/]ȫ�D�CMk�Pz3��#�	�Ԓ,�[27߽:�bQ����PeD�[�=�ie*�IZ�?l����JM�:��L���M��,�����N%[��~P��W����׭w����J/i�38ȩ׾��U�y���+�S�+�~��G��T�B���ܔ�鯛!�r�t�R@�tJ��g�:����řWϝ��+���A	�2����2����,-�]���_�2����e.j�7���a� �_R���i`��������Oou�7�D���&ѳ�&�"�*5����/Tì��S�������ǈ/����=){G�]���A2�Z�����5�T4�|UL��	f EC�$x�ZD
y�95��~#B��G!*�#عZ�^CYRC�2.�]���xU�T�U}e��e��V5�ƌ�P�!g��/�#AǞ��;�6H��Lʓ�RC�uYX��CБH����_x�=�W,��ƫ�z]t��l8�#i��Tn&O�,�m���DӋ��~��[�{�³o{�N�g��(n	�y�M�I�l���.P#�|%�1"������/"���/\}i((�Ko{�}/����<!��k��~T��_��n��Ӑr��I���?������96�R	��4��E�5�A��Y����ָ3T�� yC���-<�`��n~�i�Q���?� �f��r���Q6%��4Gx9b���)����
�	C��%�>�	�9�+���:[����f	%�@�]�,��1�i�GK�̨�Z�D�R���w��G2�NkͤX��v�/cW�ۗ�=]a��"��H��9ѻ����b7��[�c#���;WVn�>��wPi�\��+j)���bH�1����^ӺM\�`�w}#8�uK�:����ςn��/a�+�y\��#2�9�{ܐ.�hL!�#�I%����y|~}�Ӱ���p���Kף�'X�?TV.�2G���%4:0�����W��G�U��Z$�dV���A�*�{�/�S\C0n�<hjL�鶞�*I��:0J��-�I��7��`�=�߽�G'=� 4J����_����,���s��!��*���j�oȔ��3�u��	Y.�Ú8�i��֫x��Gu�]��)>L
�4<L!I]�����J��)��� X<�*B������KT���餦��*&'@�H�{�	` ��a��(o����_�>Oj#�
�j��[��	�@���*O�|�+�A4Ӻ�f�_´oQ����z4�����o�4�^�ɬ]���U��D|�d2U"!`�t2��h�)=�<�ܟ�ω[�:#�Sd5/1�`�>�����,d�5�nw$=T�=�J�\�k� ҉O���fqL�EV���S�o�6��i�N���"WKԃq�-�	�ű��>�N�O%k����`�ѿ%�KC(k3�S [���~Y$��e8N1g�Q���"���[�B�gS�n�#��#�>`5���{�5E$|�sʌ�]�����Vsv<��d����'sG�+^L��=~!��R�6�$����������h����"k8��x�(��t�_]�Nz&`��-u�b�C�����{���^n��.���|��P�N?���zpաT9T�J=@���oʖM��kۑ %���F��.�s�}teu������1]`{N�0��}�[�I�a
���?}4DM|��X�"a�}>JIЪT��J�a�Ft���;�5�+����������cA�v�z&F9�����`!���M�S�Еr��PX'�跪��~-=�P�KBiI��-)֫ۥII���\�Z��@*�1�n�Z��58e�"n��L�Yi+�ns�!1�R�*���e���t�k�w�xj�� �����{_T���ؼ�q�f �N=�;_��K�:�.���X�z+�&F���xZ!���3R�������jdJ��eR�������zas�|p^M�d��0e��O�3�dl+�QY�ҍ���>�7�o:�y�]V�x�k��P�9����{q}$z�Ԟg�ܿu��)<E-p��}�0x���S��I!��W_��c�(d |�/�%�?]:ړ�Ц�ZW�FtҜb��=(�Ԟ�0%�}1�`),
A���Ro�t�,|���p��S������>[O�!�l򍀉��E��zQ����w1N�a�O�i��V*�˥2N����n��ip�!�<�Y�eX}.?��,��SrG┴�C��v8�A��� E��[�I���I�-]&��&�{=�sتz�hrm'$.����]ޭ�?6���	�fA����<S�J�;	�^��{��P�o�+��ha�"T3��X�|�1AL>O�S��3����g���`��!�a!�dx�����[A��r������cc�J��,ALn��a����嫟q�Q���jX��s%�*�T��ǎ�l��ɗ��o���\��L�W~�����(&!a���@ɡ�t���w횯~$=+�8�;�`�J�����2��}H�Udon��8����C�����\_��*��\s嚯�Z݌�R�:6��HN�|���f����[�?� ���zd
�KwX�cN�`�GP;w�z#��C��t�?�I��;�C��A�z-�&��If��ZA2s}ۖ߶;�P�h��Ad��3ԩ�H��P�Am	(���%���u�ޯ�����ڙ4�l�.���=�7��1o,N��٘�me�u�F��Kl���k{|�X�]$ƚ�hl�OgǱU_��1�T`K�~@�]:�8t�A���b�hW� /_�Lck�}� �pXJ��*����I�,�sH)���L��ivi-c+��{��l�soC�0�V��� �訝�S`͙�Q��&4V�I���~�����Ϸ1�~"����b� O7s6ȸ8K�Y.�����~2d5.���X
�Xq���"b�����|�7����:Z�.�
�A�i<m뮃�q����S*,�M]G���b|� ؞��o5���l�^5vf�ʔ� ��'�~\X
�,�m�YFQ9�'���o�
�ǣ�]ɀ0e�QE9?��Pܣ�.�3��������%++��ݾp5՟�4�6�ߘ��(9����Y�x@��2��o�}��"�W�M�;��X΋�g�!�����F�P\���k�U����]$̍/�֧s��!��(ӯC1V�{��N16a��v�@��Rz^qԿe�w��0h�2 ���I�m��ܜa�DY,�~%�(n��c��&�32Bm��;�~gߕ7�lٓy�Ek��I2��L���YP�CT��&X��k%@쎟K��\�2��ns���8f�H�upL�?�����������SkLF��Ľ��.�w"����׆Hm�g>�L�*ׄ�|K[q��L)�#W z�
�����~����R�������ޑ����no�w�=g�1ĭ��3�C��7���R���k:�f?0������`�J9wÑV%/؜�J�ș�]�4j=�*T�"�=M��3#���lH�u��Ĝ����8gΧ�͒<��G��"LgbZ�)��o�B�dT��SM��aۗ�:�A8x��Y��oϝh�ښ �M/)�IK[�n8�J�8�N<�P�e��ޙލ)�Hq��@�A�;�L�����*�F�]���Ο�D��A7'�D3DqB�L�?��O歚	FJP���H(@Q]w;3�	'ն�c�p�_A# {}�4.��ℸ�"{���$�A��\#~Y2x&�W";j�#~fJ�8	�E���:P��G۲e�f���;X�G��E8�Z +�lg�#Y#��)�y	O#b&&�m$5{���Zؒ��[fu��L����&B���褞�������IYJ�����z[)[��Op�+��6���d�.�"�8�V}ugЦ��3}�yW)j�p䐗bw����Q֬?9E�(}�aqe��g&pf���t_���a�#�&�fX��<��ܫ�l������7&F�T7F��j_�+H�si�6+x�aj3ģ��a9dzO�A6�T�"��Sjv�k�����4�&�;<�^�V��˪�$�n�����w��z
;G&���$�c!�a�:���A�ʨ���vu�^��؞v8;m����4��\W���M����J�W�(�(Fϕ���~{:�p8�ʰî�<:�	szU+�&�^P��@�����n)8��g �<;�r����xJ�� ɹ�r��9�Y�a%-�A�������1`\�	b/���9^��'��F��dp7w;�^�9S8Q�`( �l`D�n9�^��_��'����^/ x(�x��1��x��T��$������%z��CEv]�>�S_�*������D�E�s�,�. ���&{d*���� 9�&��6C��
�,E��F��9|� `Cm��H�{�RdZ�*��e�[
)����`P�S��%�����V�I�<2;��]G�aCs�y8)���h�R� �@{�#�K?˥w�mlB�k��d�Jx�fV���.��b�� !�.�]�E=��� ��8��yz�y��P^�W��U8��J�w��<;]i�ψE��mP���Oԏ��@^����6nA�b�j�%��1��u`o�$��ڳ*����y�z�'��Ϸ�}���	Vel��yCY흽�������
��/�����LO[8��w�N��P���(T����d�`���n�) n�2�GIU��}���4o��!�K�D�C4�3{
	PV-f��EO��dI�Y��������;'�'��셝Ҷ��s��E-�l/(��)���@��["џޮ�E3g1��b��y��0�	��L4r����fF�aYՇ����漫�S��h��p9v�b�0���)3�F(F�$V��eJ�Pte+ .?2؏�䬢hl+$�d���C.�\�-ݵ�w^� ��S��T�Tz[;�D����=��R���jg�!�E5G'���\�]��M�魏��ri�c1
G�R�5�6��4-��$ZŹ����>�V|H�'ֆ׊��kE�������� �L��VB��2EJ��7ꨔ��	�
��MO��Р�ׁ��0�v�d��qe�#�����y��r��WӜ���y�6c�&Z��t�|{�
�`Џ�����[�zgkT__S�A���`_���>����өȥ���Ǩ�8Ep���;uH�Bݑ�]�.���*~�I۞�-�$�9G��|�:4��4qj�W��i=��Z�J�pjI\)6��9Nb��S��� i%��0X�+��#�m�Z����ݟd����g��02�U����p�1��2ZB��wMH�Ȋ���.s���*nh0
���$%��
�W��B�-�8��LG\0�2�|`�$���V3�@ �������{�RD=��P��/�h7CWf�"uE��4>oc���؊ň�X�k!�:�ε6�Qj~�aW��
���!��g����b���+Ȭ��.��DU|K}&�6<$;�ݱ���`R�o�{����m����b����MG� �E��;Jy���X�Q��^G�]� I��\�f���R�	݉�)�΢t�C��o��ydp�к�=~6�d��\HW��S��E߄ZF.*��(��TV�������L]�� ��bf[�Ԙ��
��E�E�\f�ڬP�Yx����'u.E���[e��J�k�E�ȱ�{Mvܜ��� 4���{p�Sj����.��Y�!�=k�g���F��2�1g�+�����uɇ|��\�܏k�eS[�7t�߯N"�a1U��E�~-�j�Q156|'>��w*O��'(O���Ϭ�/%������=#��~�.�NT�  DA�i����+����E�f��jP�Μh��k$��J>Xc@C�o����,�N�}�i�����o��#�x��zNN+մ�1l�w/	��<�7�0�J ��� �
�M�E.�I�5 ,��n�n��L�$7砂t7L����⓭��@$l��ˀ����QL�{�*��`�5B�}�ɿO/o���bkW��S�֬�؀�(޷���:��K�4��%E�i󱓂}��W�xJ�"����x��0�ݾ^%�]0&���OnX�u>g���B���!��js�F�r#mm�����.���5���9��j訊p�c��W`��EkoIc>5��}��~�����t��=�����l8c���c/-3ࡾ�w>)C�>���˫K,��"Xo�,���J��iá�CLy�}\3%��yX~^}�����bQq8IR��~�L�3��B"®uJD>4�����J���b��L��0��ϻ�w�А`� ρ�I��~�-E��FaS52��P��e!�򘫞�uD?���f�M���aȷ�_�UH����S��	���;ҡ"ȓ��E���lK������]G�(v�^)o@��"5����ci��n}�A�6Lo��N�Nm��>�j"j!0��>�(,�m�{��� �*7���5�N���XeF`�w�"i���*��P�[b���3>,��q�ht� c&����P�n4��3���6D�?	_�}�ac�� �$a- ��2�L����3�d~ϵ�c<�\���K��t\�m#�oC�9��F1���S��	��4�H�\���}��
��X����NR�|�����ß9j��(qF�z������=p�U'�r��#�d�>K9@��>���ͫ��.�}����G��\f�eȠ>��9@�R#�\���'u_�W�A3�?� �?$����r�����r�- ��6�#�
4����K-�	��4/K� m��G~��z5_�2)HH1�Y�&�3��@��9���A������9�'��ZJH%0�]Ҹ��@Gm��<�BT���~����4��P���S�8�.��U�-���꽐�K�N�G�RڱŢZ|Q٩:����k�����b.iƃ?j �V����:��ۦõU�4&Uw��M!�V�b�W;b�Z
*ts�������#��W��e�gN- �N�e��k ��`�ȤB �J?e�;H�Nͅg�z�(/��'c�U���o1��j*�S�5f��h�o�C7����J�8&R�Uq�*�hJ�EH7!E�d��M��֦7�k�eez�������DI S�����΃~���AO�l&���M��2��g T���9��V~e�.ik����*/��r�+�	�'�j���f�U`��A���/ɫ0`�>��]%,lKb�5 5[&g}/�;2��D�	~���u�ջ<C�]~��������Q�{����B[�n5�Џ4{CD�
�����=@��$�5=�;��v�O�>�LߑN��ҧC/�0���E�Ǒ
��n�M���(�z�T�~_f���_J�S�B����K<"~�.`���$�y�;�g��b�!q����v<�$ewP5�z�5����Y�}+�|�����-��p`�T��f�4�L�]��F\���V�.
�W\_A�:8����Ex�'�ۿ�ۃS�(���&�ց�x~D���SL�#md��w�y�;��}�@��+ދ)-����tg���j�w���aA�n��J
%��\���bK ��!su�'8\`�`]'(v��*���B�F�v&7��/�|��)]5�}�ɠ�Yl�7�E��`~�����=���)@�%�w��O֖���3�G������e����8`���p�b���%.�Ń���;yb:�G���Glig,:��Pf������Dlk����񬕴��;�Zq�r{�`Y�(������P&G�Z�/h�������1qSª1o��L<�(����N)Ñi���(sS��<��[_��v�k��i�dk�	9�����y�F�*o�ͻR���Rh!�y�a�سx��/[@��a�8�m��P�{-F(N�|�� ��/���U�(�(	�v5��$a	�u�����W����+X&��+�Qpŏ�2F�ʫ$_��5��ۤ�u[��.f�J�F�{��e���)0�j���np��!�z��gb��t�I��iM�(f5���s"��ҩ�z��B���]*F�Ù��}� {!��f�0J�<�	'�0NH�C����k�����O�U���~�[�n��s}�s+�P�G-ct_������މU/mX����l��� >��^F���N6ӆYFc���_��F�8�q�>P&�Ճ�]c���HT�EB�ϯ��k�kM���P��p���m�̳�v(����A+��� 	N��i��o��A��F����� �9��� z�U(�j�`/��=$��>����"UnԤ�
� �����2%b�4�����Bt�L@/�D
��AV��2֛��1��K(��e_!�[j�3v�K�:�4*�ﾩ���lOe�֮�����0�h`���z�Zm�\W!��k�%�3M3���%����3-^�蚗=.��)�W�kQ����*��f58#S�@�;c�n�̱r岙ď�"�%�ӽ�*�/�v e�m?����n��㴘9�p�����$�*�h�ƀZ��,<.,h�C,��?=�i��!c�#.�'�GS2�p6F����:�=�*s�z�'L�臈 0Cx Qp�̧ ;����.��ދ[w�q5���8]W�z��_� �f,�[G��\�ڨk���x��!���w�z����+kh�5�R-Sd6O�o6��k� �p�,�����h��7B�o5.�L�j�Rꠁ��h ��Z�Y�y+��~��cf�j��$���]������HP�Ze�[����c��,�Vz�c�C��[O��"������<8�R��J���NYiW�m��'Ɛ�1�+pZ���8-���P�Na��$��v�v�Աyf�4שVbM5���ޮ7����ge
Y��Wy2C�˟S=����=�4��f&��G+B�#��ޞ[}���T9�a�.�/�F3e����0~�##�U_��	�i�]�F�Nx�2��z���
�6ʿ,��L�"w���L���7m�mKNx�ٞi��I�ҩ
��-L+#`��3�m��-(KX�Sz6m�p�4��nA��y���4x|a	��y˅��&	���n�YƢ�~��v��y�4Y�X�$�Ò���{t��1z0����9G[���|�y�����? ��Wxb< kT�8�,lPv���z	�}d:C�/���v�M�����r�j��^P�N��c@C�O���=�����<.N�<�פ J��^cl��Zj�y��"��,1���Z�3���e��<6+�Ti���Z�����JZQO��b�pʞDq�)��v(-��E�L\�!�!�,����[`����~\�)�� ��R�C��e�|��.o9r����ص�eD����>zH��n'���X׶v����� �)������ɿ�.�GG��[���d_θ��%`�j��(�}���Y߉��b{���^���FR5�6rC��a���D��K��4������N�q�f�C���D������.���9���V��\6'a=s2�?���ɾ)�DBp�ITA+�[��ɡ��s�:~�pcƓ�L�T�5\�*��ϖ�\/�>�7��吕�pi���8Z����o{�-�����jg��TqA�U�l��ެ�'q�lc�	<��F�枳�A�ѓ4�n|�~����W�H��F�ұ�,"��n
����^��̬��lxf�RĻ�s@�����պ�Ď11�'H �q�����  �#K��?��p���:���:�Zk��n>�"���
��JY�g4h��7.��J���+��e�%������G2%r��`P��@'��a.#ѐ�i��Tr�j�f�8p v@7��5t8�#
V�bُ�J������cf�aR��VyF�g6��b�u���J���?H�kpѝ&�$)%^���!}����J_jg�s��6�X]{�Ɨc[�J+S��\�?�œc��W�~
hFP$ ��d�U@3�o���b�?�ы�1��B�ƥ���E�^6t��7���$z�GDa��+��/��V���ͺ��ʕ��YFc���,h.�b{R�g&��V�������h��k��JSaٽ��*���3���Ԩݎ{=D�Y���5ả�Ԙ����!���u�,6t�8�5)�yt�-���jyߑH얗"E���v��a��+V�u~5�P����2�/A��W�d��$��� ��E��w��7l��.t� $'���I%�c֑�]��X��Km�H���.�:�
t��3Ѣ*�ءH��)E�7
�+��x�t�9�z�r��?�U�3R���G��[��7ŏ8�p �^^�L5˃�O���Z����C�.��h��K�Uc
�P-�s��c���,i��_W�,�9fq�MA�G����qi�q�ʘQ���b&qA���`~��MQV�Wk.X�\�-�����~^߰k9MҨ���&�x�xC����hZJ�FC���4��^��CLA9����Ѫ%�8��2ި��z�;�5`���ix����-ϟ	?��/}�qݢ��xE�t��c��Z�K2���5-�S�E��s�y.ny']���;�w�;���>���"�^V�GD�]�ub�H���)X?�����-B���*����ӵ��@6�ǭ��N���H�^'��[r�KTG�J�{�����K�����M���ҕ*��I�Q����N���D
���bEm�$&�%�U���)�� �}�϶��|+Q���q���$����XG�	3{]-
j�yHN�	�w�lu4��7�AČ�5g��r7��y���o�vb�F�%X�Qx($B�v���O��A#�2R�`B�	����35���3���z���Bc�:R*r��p�K��0!�_O�y�_�'hR��54w��I6?�Ť�k��1ɯR���[��K�,jbD�z���j˗��r�>���&��hy���3t��4B�%�E���I��m�������4���߹�P�|�J e�
�U�c���%�jM0�&���q�J�ӊ3{��`�,���jr?|�zL�b�mޗ۳�Q�g��?� �;��ռ���:�*$z�C���)>c�]\����~1� ��M�����?�2�W���(v��G���X�X+����@�"aU��KG�H��!�����3}> �0�
�_r,G=/e�Ù��b���31Bio�D /f,��S(��_o��qpU�V��,aq���Զd���|*���x�ڡ29��JgyA"A���c+N��fE���|[K�3��$��8J'8�%���c馵��Ұa'�� Qz/�Z�Pn�:��P0`�V(o�[�'� �F�ڠ�@�*u=�	���̑BиwHY&FwI��ku+�E�?��@�N�9�C��,vo��D��Ϻ�fx0q������y��۝o�U�r��!}�����X�q�~�v��W#��ٞ����t@�@�ʴ��ց�2���?��\D
 �������",�y�D99������	�\v�q9-b	-�ޘ�GOh�1|��Mk9tgC��[��+x�[?�"��O-�1o���z���j�{c<C���9[8���	=*�����;W�����'���DЇB���8�T�NI�>B�I�*ӭɻ��'Y���v��b�}�;���V�BUe���`9o(�x�b�_��?m.�ѹDU����:CTq�f��`W�V5��NC�Y�[�E�DB������`��gi�����
�����rkk�mt�F�~��N&ދY��������8ec�	��`�볤�Zj�\��P+ᨮ��-M��W�5!�Ä�]�6�7+�M�8�-�ѯS�����鞶Zz��y}�K��*�e�nb�ɵ��f��o�~`($i���澨��/�b~�#B���Z�!}�c�*�qp+�����-�����ߜ}~���ar̅�#�!�T�� ��q�����A{?��Մ��D$}�c#�ށŋ���BG0
���
 ��y����`*��`�^e����4P���~Pa�P�p�L���S��QZk.���ʷZ|V�B�#>Y�"�J���rؓj��5Nq�[��u�!4������0�t1;lW!�����;&���ܝ�f����؀ ��l�� ��!u��h��	s>U)�E5%s,o���UI$^��3V�!���HL�+��0��	^?��-�Yɮ�h�S��aP@J���d�i�gWY�$�/���k�d�����cȇ:�u�>��N1�[��?")�8��V"o��T�絞�5������R0��|����YFm������jX���7?߾�Yp�GSq�/ɣұ�z�L��MMYj��|n��+0�Q����c�Z�j8��h��K�O���k������C�~���	M�w�@?��)XBu�C7N�T1�?���b@�߼Zj����k">f���SyƷ�N���J��v �1�wt��KrQ���(�Om�pD'Y1Q�%�9�p(X8���{�}�r�@7=L1!�R�9�'Kظ����|5��������E&�񏐵 RSO�P��=�Z��2�~>hc�Oı�d����[�cLC��ُ��^"���7�g���x�*�����)Co���p��D�i����%��]ª���_���=#M��@�sݪ�&���y��䶗�`PM�����>�ˌrቖ�û'�`>'S=ؕ�{�",�:�	r�b��|�eUk����3ǥ<�����<�&���Am]Qi�O	�F �6�F}"-r���z1�F����k*��Q�뻩�V1��ٜ}���&�v�-C;�9\q�:�{�l�/��Ʌ�ԁ���8�,a`��C�e%a�qPQ=%�e_���н��������][�!%��Ú�ܧ�����T/v2�!?fv��>q}B'>2����[���ͪ����a�&���>U��1����g����;�Tn��`�n"A�vu�V	B���NE�������9�9��U)4� �Avy�+A�2�۞�Y^W�Cd�cG5"��Vp���z`�o3#�ӺӦX���r●��b�F��'2?��y�?l~M�w��PV��Nkq<�YмŽ��I�fe��TL~c�E5���Tb跞<eH�O�b�����ی�B��ŵ�n�+n���g�|R?���E3��ʣ����c�qt)����"(V)=р&��xh֌eIKq�GI�u��i�ͶiNLT��������B*/5n]�g��J8c<�?���֩�mY��}�DJ�;�"[K�T9-9�$�"�g=51��r��C=Az+堚��������>����I���jO�9�З�7�+3�4��G���^�AP��='E�7�d����Yr}�
��)�l��7PZ<� e�o�C�c���K�2?a�(׳���<��vK�ʵ��~8�}����ֺ6[��.��u�Ғ�d@v�+/��L�,��c�|��(��ˡ�)0TQ��z;>v��_C���,�o@z����I�~N?�!q��rx@�n�����>?�席P�$�b���rq}�i=�����Y��[d�2�,� �|o_<���|�"h~�����S�bkڸ.�鷟��Z��D>ɠ���\���PW�}Q�c��
#-�̜6���"�h[dUUo�����Ê,k�{t=�3׻#[t�*��aL�*O�i��/�j�ꁟ!�f)�lABv^�<H��l.�oݹg�, NvB��ERA_s����O�Um����)7������*V'q/�����q>�D�y�V�z,���� k��/{R�f��N�e�ӟ��Te�B\��a�Vk)_IQ�f�]�XjgQ��9�f]�O�Dj̞7	g5����l0ot�+��p������+)��80�M��|���"�(f��<E��^<��h?�곃��J�$@�dl6�ܫrp��MV�h��҄^����~=�²�.�����@��j�R��뽸���R#�Jka��mSkdW���Se�\����kf/Þ~2���ͤ�?i����i�#K�g�=���e�#W/�,�\�gd���^`��|UJ�'�\qĆM���G��e�U����-�鍹���̾��-���؁<b�T%�!�K7˫4���E���hd��pZ�C��4H����:�ZW&}��?�y�ϒ�M�0�O���	���/s��߿�C�I�DK��9'+����9�Mvv$��T�'�7XΓ����:�7��,*��ۛ����מZNd�M;*��m�-q��'s���*o�w8�O��a���]m�,f���p<t� P�G����0�̏�,nz���aY"$Z��LcM"�H�����Y�q
uhØ)�o��Iװ�e��b1Zm������(��K�_MO��kq��n]����6�]&}�c\Mڀ�~>�?�V�Jhb@���{t��rw���(�N�*�e�e�dm҅ŰW�GA�,����<!!o2:.��xه�8��p��<j�<Q�MR��AE�ص;b��/z����Q+p�yI�O����\� w�G�Nq�3�7K����G� h�f�� և��t-�Rs��fD4�I5>muM�B�@7l0�jr�$_K����O�Z\Gh��7��cY;XQG'xR��V��,�}��=��a��Na�d�Oӿ��(H!!bg��Y"˯�M�Z�U��@ꬆ�X���C��fT����B�JP$���VBn>)����7�qE`�W�������*H�SbՒ���4��@߯�ӤJX�9�ϯ�n�;p�a�x���m+�-O�^GX+N�f$�7��v� �砓F,�I��ý�x�I�	l�&�)Q3���;�bX6�2���ma���_ab�8[:���z�g��.mw�I�)`H��v1u��̌�"dc��W��L7�5��B�g��}x.ώkoF���?��>�Z��j� UAl4�~'�>�'=%\f�/q�Ht�F��v)ʁ�wb�u���qG8i�铠%��8��x��O'�H�5�ig��2v��������ڡ�ϣ��᫲��s���E3�_�@/J8�T�W��%H.�D�� :_�����tڲg�@.���g#(� �'"Q��x)�8g�akLӱ3n��7.|T���TB(��X�A�*p�K�-��hy�^��k��yyiO3�a�hu4}HH)U�*�:I����Gv�����%3jC�`ErwqE2�1,+ԥ�2M��V��cw'U5�߄nt�p�� �œ�uC;�[0*V�h�$U�uI�k�e\͉W���ҡ�
��8�p�:�e������ꀺ��:�G�K����anIY��Y�z�����vOL�E��;�����,A`bo�������	�U���Iᆁ���Ys�"�T�/�����ͽ�vKצ���~�m�k�1RT�L���P�i)*ƋʍSV���݌Z�^��	������~*�+�(��������}���lZU,�3���Rsը�PM(����d0�����}ߒ\����k���5
!����y���e��D�W��bO|[ j-G�_��[ h+�A�D�`(5=酞!�ޛ��(-u���m6�SS�Gd��k�M��^ٷ��o�嵓���iQ�ӬD��
=�7b}Gg8�y�Z��-�B���M51O-���ڒw7G�aa��� �˱��r��u�|��(*7��h*������y!��2�Z�]��p�U������<#�Iqi:�f\�iE���M�㷲�ϙ�Z{�j`�U8��1�V��,�9�������BOS"�J�E�;^��2%rlh���g5�bF�"�ҖI|��<$ӎὠ���
�o`��qi�z���D�W&Ts�p��������2HB��r�1���4w|}:��VJ�T�T]��ժ�R�n)��/�	l7�-.��1d������;b��%0G�7S7��ڞ�ocP/lt�A?�t<?�,=����K���u�_���\��*���[���!!�L]	��Y�	���zaV����Y.��:2Q#���8D��{%���tٞr��C���<�&�x��14�z�\o�簣썮	��:����Y�	�v���)��۞/�m�[_<׳qKI� � "~r����"�P#��6�}@S%�K���&� ������{��.s�
����}�J]~���6}`ķ�R�{�pL��E]�+*�a��dp�@&:��Vo���.��#$P�V�X��zK���4F��*`C�g��iM��y�5�뮲�ڨ�g�"d>ZL�t�xX�R�Ɋ��+߸��Kt�5��˞0|��ˣ���C��m��ێi�^�4�N�<����]&Fm�'�{p~�Ȇ�>�����0�.��J�N皹��ֿ��(�ъhnP��b��W�.����_^�ÕE'�&��1LH,Re�!�X�EB*R)�RAf�[M�T�;�C�y�l�ǅ���u?�"����,u�(���k�o@S�U�����Ry6C!���A��Z�w�K��%���'�K�r@4QnӢ�~a�	ܿ�V�p-�<P{G;n��f��6"��6����`����u�K_��L(]90&6&G�ˑ7�T��Pz#L��9r��`2���:���/�Q*
�������K�<<��l�M}�S��i���a�7��>�VZ���ϸ
Nv�����jNe����0Z��n}�v�y҂1��Z_n�"�����m�*f
�'�S9�4��*�=1����%X�'���h���tS9�ſ%�/�w{VA}��������������1��4��W��4���i�ݾ�ˊ���}�DQ�U���� ��RT8GA|�w-�i	��j>x)����赥z=Sg���7t{�蓴(e�t�n����n�����6mPLi��#�QD��(��m{��g�y9��c��J��+�|*r�^���`*��}j甮�ծ��^��s��m����_�@̜fI$ ��w:�g����R���Z�¼����^�Y�{ևE%�������5턢I�L\$��X�Ϸ��m�{�L�y�]Qs���<@�'���-U?n:��sh���蹫��x�\�����=d��[Zp���)�����Q:��3G��%h����P�� MI	�I]5�����j�[ 3,�;X�A�p�6�}��2q~[���`�Jc��GL�f�*v�p��_��$2,���������FE���4�)��`=ML�����Fː���?3�����SL�	�[H�D~�H�jc�sn�b�����Xٔc,�}����_�nva��np?p��,��"��̖��~�����蛥�V��T�zɒ:���� 6�# �yF�^T��4�6?�����L/, =�ǚ�~���2d(�Ť����|��&-}��:�=�$k�cߋP���#ZH~FgQ���G+3Ԣ�RC�)	�e/x*>1�Ey�ʣCP����`�^)!�LŔ-�m���' t�����~b��4c�Y�֚��~)>O�嬑l��um@{���OX��P�S��#��B::#0��rp2ue|Kdr�Y��]P�(�I�{ڼ���Ԝ�W���hQ��/�-�?�B��m�ݑ��B+�H �}8��C��qrqK*h��|��9�񌈬r����>En�gx�-����c;���f�����|E�|�ќ�V��Z�^�*_��I-�����Tu䩈���v��}�'�э��O贷.�U�h�sڲ����7�_��O�|L	��?y���7�J��ڸc~F^�ߊ���$Y�䟬�}�_�䊌%�/R��c�~�\�f�ܕ��,����J}����|rZs�H�p�q�ˍ��EY�w};�N0�j��kcU�k�.X��@ �u�y<zo#��4�o��������;mc\�C���X�V�2�����:=��Xv#�S�~,Z�F��-�p��R�ҹe�f����u�����':N�rȋ�GM��1<7��{5�Y����z�݄�l�Ta-����� vK�tK�Rl�!��E<�j�oQ�Ĩ�4�"k���y���8b�2� �LR��$Mn����{����O�7��n���'�c���u��Q�Ln�lFE�e��/�S*��lϏ����V���d��S��b�&�ĄfH�F�,T�Pj0�'@k��^�l�n�Y�F�ɚ��-��H�v+U0�w�(L�|������>EN��a9��$� �f�֕��:}�ԍ���E	Æ�n��qP���/�i�+q�'&&�)yOEI�]���xQ-���VSTq�Nw�v�>7R�/��ƧI$Wr��E2�܄�Dj���H�X��~�yͰ8��T Z�?!�vVՑ���a ��GUj�e��є�8�l�R�{��Bς�ieJ�Ҏ�uC�����U㣜H���{I[�Զ~9���d4�Zx�.$��wF7�� �����!p7+6����g^T�@-����9c0�@��g�\<�}Z��/�7��*��-F��(^�[�j��������PW������ױ�)l��FAg�V�������I��̻�]ƥ�����d�����u`�7OgXA�d�Ê�/n��q���r���wf��(�u�r50rQW}K�KAKP�P�O�D��D��Z���}b�ir|�������<���;����`#z��pko�i�Z���(�u�W4����J�1�e�!�<+�V%�h_�9(����d����B�d�1aOrX�q�x�F�z{��6��{] oj�_���5-@;���(;u�D*mw섧?U�̢�� ��4^v�5�)� ��sQ�lM���u����b��~�sH�?R{u������1FM�ƈKNr�āT��0�Q�L<OFG ��� �$�?�4��_��j��;����͚R��2�t��yF+0����c�_ņn���LL���!��8���+��"��G��������ނ��h���Μ��u���rLU�[�'��
o��I'�P�o���Yuz����Q���;����٧^E@�"�q};7f>A�:z���}�j��� ,���/���2��~	o%x^D��G��F�l(M9Ƚv�@���ß]�X���vI.'�#=�n}!7��z���Ҍ�D5�?���M���A� +�Ι��J|S���BF\cBS��P���b���f�ܢ�~+��៪ 7�i��[�`x�7��)[��k����}� �0g��?�h��J����\D#��J[�K%�=f�".dQe����Ͻ@G��'f)�~�̷ΠP���`�NLV�) � ��v����d�S�x��e�|W�̋=�\�����'W��͡�M�$AP�F��A^ڲ��H-�O����z���Q��zE��#�:�� J��������%g��$�g�f'��m�|	���|@��p����϶��`���v?���#!��+e�/��s!�����A��z���T�k���M����M���� 1�������W���86���K����)j�bW� ��2��~��!@;�������c�{=���:��W�c{�بʌh/��#_�d�WCrnW>˞m3�)~Q�$�W"g ���0ఇ��ڇm$Ou�,w�H�����W�[M���`q����0{X	� U{`.�L�D'U�-�(�'���n��_ ��̺���!�=�F$T�9�՜h��_� ����x� ������3���.��^`���-ك�}
W/G����� |<��i���7.�^b���+7�z�'_������
B'�#6��(+/�Ds<�E�DL8k���lg�?�J�8]���X޸����;�דA�N
TSE:�nڇ�c���ژƖ�3j��`�]�IL���3���S�$8��:�e���n���3�:d�M���,t�e�v��1�i�ό�MfK�5ʜ���?���z�WS�=�u����o��U@_����kAHͮ ��Zu� WZC�V7�e�=K)�ͯ�}�,˸�w���op��ʯћ�2I�p@/5����7��eJV��!�j���+�[#��v���W'Z�_�Om�n�Egq�V�ZE��|*Vc|���,ߓ�ct�l��5G f:rb��J���v{�x��J�:$$�sV��>�%��ॉ�,;�~^�L�y`���ZK#U�@�ld�����"���!<�=Q-g��b���j���s��?��/�K��V�l���>Ob����m��e6LQ��)��46��eK�F����I�L@�31��f&"���t��'H�_�8�l�@� ��>7��3tpK*�O�ӡ��/S?�wR����0s>P�-�DGt$Y���b��_=і����F��A�г�s��È�"��c+5��Z��8t`���ǲ���Y�l$<�\R�V�nJc����2�A\��3�5���3GJh��9���70*�j�
�_����>����O(�[{a̮_�{/l���5��hC94�K躓��m��:�G��� }�J���)��Z_�[�ZК`��0���i��/�0"���2�c���Ӏ�� <��<:I5���-��\{��@��E�S0bBڼb���IG�O�'��?)e��j=h4{�mT��ȣ[!���ɀk����[�B_f�P;�i0�}�i�������jC30�3�;�����T� $�y,t=28R�4Dz^m�_�1ז%�
˗o�7jO/���M���'��t�������b����l3k�e�4c�v>[P��OE��s���.`7H��W-i���P�?�y��5Q���^�T-N��8)�jVx_�5ʺ��#������3'͢�ult��7��̛�|ƞ�QT�Er~@��3y�|�Ѓ�1�@����P��Fs�K�uQ�|/@V3��&ȕ����u=��L��02��������˗���^YF���{�� �z��&�ۤ�ࡣ6��4��@u�D����[��-=E�$�����S ����u�~���÷y{���ʰy�}{f6�T����-{�rHY�5���9����67��ǉ����MB��0|Z��{f4ѯ�&)�q����܈*��_G�ֹb�4}<�N��Q�L�(�j�Q_| #�h�8����@�i÷�i�Y�oX`�>��&e�W���?�.7<US��^G6{Zc���ѐ�>���{iH���Gw�!j��
�� �{>6|�ݯ�x����6������)�����-*��;\�'P��Zhk�ә�e\�)8���c^��n<T�$��/�DIN�������&`Һ1W�-n�Ľ4�����O�W�X1*3$]���jq��r���uY�,2���ʺ�#|Lx\�����4�]P{��Q�4�����ZZ��c汻O$�l�ɤ�B��֠{'x���59?CZ*�Q�Py�b����m���-���6�*1����'�Ύ��xT�����U�G�T�f%���0����﯁P�%k]�Xϓ�L���_���Z@G�݉�գ*N��<��'i�7��#����×嬹�R5t�;w��}~���2o�ZYcك�a
�t-U5+�Zzk�6�\�s�w5ІX�ཨ5{���w�i�pN7�o:��)�b� Ԇ�-�k�M�GP��Ϯ���MH>���0n7��X�[Jj �e0ח`��G���V�u�����r�B��91��'m,Mm��ʭ���͒\i�F�}�5��7Qշ2+G���6qѩP�����W���X�'fXM�R/,�d��~��[�2+f������|\���sW|��N��u��A�G͊�⒃T�8�E�� �d[/��k,Q|Y�C\V�%hK[.�1�R����7O^�]q���^��#0���_�a�?kX�a�Wi;��n��;�g�h�Q�[��Ѝ�"1������W*���z�����5'4��
Ԋ�t��,���}7fC���h/0����{wB^�a᧏c�r���^{��gV�x��!�'e�٨rS�=�W!�Q���ք;3fh;�;�8��k�C�9����H�pD���X��R���T��ӆX�"�v)k�&�{0���w�\�=\Fpb`5^x
�|�	�����D��fq;
���z	n����t�iB��n��Y�4q�9̳aX?����*O��9'������Tt�̂9{7ps�H��
��SΌ>�ڰ��z߻�n1c0�<0���=9����/��	%�ǰ|S��n�W_i�>�3� 
��	<�4%&�;f_>���:tƧ�/Հ� ���Y�f��x<N��И�^a<Y�!~�L����`��,@�d�j�,�������,��V��g�`;�w������;+c�����fH��xӗ/��4�E?<7B�JI�6�d
��U���n�V����Z	��,y3�uVz����1�/a_2@��?��d�2�T��ĴoK��E'���<�d��%�gM��Ji��x vh4�A�"90C�E) �2�ة."|�n���iF�/�UP8TS
����O$R�tH���n�Kc��8^)��,���͇o��[G#o���lÓ�[�<�N�@�Ɩ�_�QI��n���#�iu6�4�ȝ�[�1����w'�mZp�W\jt�ǰ����Mp�8L��m���<���`PV���0i
2��C1Q�"��no����k�[Ķ�{��.�T����*J���:���
&��L��~��s�����a)}��������_��\ʬ`���Ne2��W'�զr$މ�P/Ia�C�:�&�b�[i�{�ԫ�q�w��}�e^���?B�ʡ��IEK��X�R�!;v��:�+���3�ܗG��R�ڪ��N��dp/���,��m'�%�V�ߵ�Z���H�.q�,�3砎�#��4ГS� �JT��7U)N�ɗB�I�m���PԮ^U��3�;�bC�I\��"FG�m��G�oiͿ��������DdfX��,!5�K.n�|Z��;��Y��|=ܛ���Wf�˩��-[,Z��Q����R�\���ؘe�~xKt�i�tg'���g�+V�:�z�o*����Fݏ�hGV�`�RT)�e�s��,�_�6����?x4-�af��DJ�Y����ʵ/���������n~hs�j7`q�}���4O�^����/Q��7I�C7bP�Qzؒ4��7��$�C3١帛�<J}끿e�P��i_�Ikp���@6?�׷S�Q^����{�^�P�*�ܒ?��'��9lZY�#�}�vև��zB�a/�8���R���*�v��y�t_�l���>��-����֛��}���9chyaͫ4�"�,EZ��ؓȦ�X���ѹ-��?�WM�'>ͳ���Vt�z�?���G��^D���{�O>�x�x!����l8�ڷ����b@{Gm�I5�c��2��L9GÕ�L��	���ٔ��Q)2(Y����=mѹ�~���w��A �%�6ߪ��>3w'	*O&ŕ8#f���K^E$*5����|x����2W�j鋞XPv�!2��*4���P���V���	���h����<>�)@��u�/�:�e��}$ȷ�"��?~u�G+z��=���԰CӦ��wm�����s�=lC�Ў���~e�|.��&��]�'z��N>ї'�S�Ƽ��tbtZ6=�����-|��.ȯ�$zȈ��7����$/�F�g�p���/�e��6J��i�0Ij������3vݩ�8�J%��]��L�
IIW���I�=rXjk!jϔ, `���tួ�]d���t�z���	�u�qe����̛<�ċ�oȦ��7FN����XN�w8��f�,�����M`���r��U ���&U܊k\$�2�UG5�����>*����)��R��M�/ԓm�P�|�7{N<Ʀ[�u����y�� ���F�#\c�W�z:��c����~4�0���ث�O2��&�-��7��ȕ�C_���N�p�ƪ/������RI1� W)1�+K���������K��a4p]q��p�b+�-ҕm0�9�J��2��v�dx��#A����V>�M(�h;j�%��i	r>���o[�E_W~On��wY"꾽l*M�(^����=�UV��s�c��lZ�].�%�1�^�����vR?�`��~�����X��c�:��;��=�7�f9�]����\4�r���N6�6X2%��\q�	�55�N%�{�t�?Q3�C�"s'�s3 :/m`��FϬ/*_��-��'��!�R��]mh�K��������8G�79��q$ÿ@�~x���(Ho<^��l�@��l���vd�ƚ�z'���w�N��q'�0}cy��;0����PkhIQ%���`,��8�T��*SxR|�+���@�q��pdv�e��
pnhTW�p��%�1����7J���sI����ط���k�q�nD#d�==F"��O��Д+�b��-���rB��{�~�X�,����:����ɏb��
�H������v7}o�(hRt�âr�!�;aR�ÏE��e���z��|���tD��
��o t�	6��Ok�e�e�?�Y<�z<!��νѴ1��u�W%����;���Z�8���G��r%:���:A�#G^u�X���h��Д]��k9�9��B��f�ȉ=�t���sn�ƫ����Yu
�1��G.� �������8wxߵ��0�<�_�z������ދrd��zfM�r�Ģ�4=�h���ΣUԔ�������%�3�ҶN:�t(B�'.r>Bu�ӳ�+9�)ѐ��,�g��c�_���ț^�H>�(BN9u].���:sǤ�_�m�q]Ձ�Z�a���K�һ��?C���@�obh.}�{q�z-�Ü�1?/�9'G��c7tZ4ܘ-���S��J1�u#ʒ��?*|��mt`���� �<&��r[@d�|�0�>��G��*Ã�l2ڽ��N�FC�f��� ���Jͱ
�ʸ��,���[x��[GOW�c	둅�;�3Ͽ7�����g(�M��aM�M���}��H����>��<tE�b��<QB�x� ��h�-a���U�'Ng��$��,�l�Ef�;h�gF�'��*us�38�2ݞnND��#O׾��/�,'�L�J���.ks�����J4���D�c�ǂ�#}����<d���Ms�R�y����9L-�%�6�ӆ�k+��?�b�vWrz�0JO�,��(hz�(�ו�$X���E`ƨc�/�{ �O0��T���U#�L�>��45)9��Wk�u�Zŀ+<E{�Δ�i����.�/���78r��aϚ�\��ؠ��dӍ�r���xe��Wϣ�;�[�ỵ��{�}�_8�Y��sf��bvdэ�π�(�Ξ�D�<������t]�G����Ȁ_QQy$C�<��F*��l�{�v�%��^BZ#Qra��A�[��QY3ל��fa]D׹��Ķ�j%���P�Q��`|��5�v�yhz^Kkh��u`*>����c,.����'�O�m~��`�(��T��xJ��Z-￹��"��JӺ|#�n�kLd��!&#��i�=]Ύ��I�~by£sZ��}��w|�������"�= 8n����⪹�	�8J����}���L��Hb��Fj�0���ټ�>�)��{�u�82ja�
�Ԉ���d]ƯA��Ʈ~�,=!L��qD�)��Ɵ{�i�f�罒��	��4�6OŤ$T��T�{c�J�N��V�F�}�XS��w�!����ZH����~b���	`��n}rX>��w�����|�3�$��}|-,=�W�,7��g��8�?V���:�<&��&p��!��r�#����/V��c^��	1 ���$@d�u���`\��M��+#�YC�'fB���K���0�����mA��
�DP����$-Z�dȗ��B�ִ�_Gb���Ru�9���+����A[,&L~��č����j�)r[��� �T�n��0�M|��`���� _�e��b#����8@]Ժ^}Mϟ�������?�[� e��x���/Z�D�D�.B5��l���X_KaF��.����b�7�|�:�A��g�ӵ_�Y�>�K��Ϲoc��̓�a�>��m0̜��r��7�6䰱x�/"�e����w�Y����ڤg���!���ihA}z���T;�{q-� F��9�գ���{y���#�7v8+,���L��M@�wnZ�������1M!������[0�)��CsCm�G���B��G{�R�&��P�2�����d<���F_����4�鉹b��8�/Z1̙E�^�I�l'rP2��S�/Sb�����|�]�r�Dhgg���#���:&�D(vV�`PԌ� ��q��홉������z�|����w����W.�j?(v��@��"�T7)��j�R�|�~�9��h������s�R���l��0��1x���	����U�*쳻*ς���	w��C���D/-yqܢe4�E˿����}�
ג�t��A���KLA�}��A�6����)&̌kH���t�6�]o$�V�;:���p��m������`�K�Q�z	�����a��$�������A��>��{��o��
�o����5!��F�U��1C.�$�PL���g�u~��or{��I3Ưo8w+J8�`�S���g��"S�Q.;�8���hM;���~�F����p�ԓ{�$��A�D�@8g��A���-?�X���g�]��sW��N�U���v�VU�]lg_c����!�[&Nv�������5�C���^q!n��;�q��*��un��:���e>���d��������H��7�>��k�B
�I���p�ε��p�����M|�b``	\Xi�yp�yܥh!�"�
��^c޸(b�8d���z�Z���R;�A�Hc5�)�������c�b&��[��S��nV>�̝�k����H�\N����ē|�s8���PU�Ql�s�U�QC��^�*7���u=���E:d�<�k�d�t�&}����SA��j�ZV^��	�@�T���9E�����YO���u�ɺiѰ�V��?5�`찁)Дͽ������W5�0~5)J��I(��#�X������+���9x��~&�r���w�N=�N�!���X�e[�ϵy��H�jkZ�C=J�Սr��N�m'��n�����a�T��x��˦���%��#π�;��'ԘJɒ��E�i��n�7 a/ԩ�z���eT0e�3�r�g�f�72��z���se��>A�qTO��|f����=��<�%��S�c�� �K?ut�Z�9�K]׫��˂:a������k�W��rG%"^v�����;�i֊��r �u�[䠐��܊>���������y0�InmS�+^�lX���w�cq;���\dlS�~Dz<�d�P
M���l��!�����':��Q�@�/��lcdc�Xx�B���qxQ��vk��|>vP�O����so��ƿ3��Y���t�U����2�8N��&�덮������,�Ծ���k���FNE�H{;w�9H�FJ�hޖ�^tD|��̱�.�\�(7z�;�2Dv(��hJ� ���m HW��GZ��8���8a�9V1�m��%��v��PgB�#kŏg
(�Y{'�%3eƶa�V��:^@h1&��c?�V�ob��iB;!ʦN?s�7RMi2P.&IP��l�6�O3JĹ|��n���_E�/<���q�Yn�����ʄ���!��o��)룝���j'�mōZ4�_B���m{�P�_W�H�s���]u�P��C��?��5O!cab�����U^���beWC���G�3��g�#,04��V�q�4��o�,Š�[Ӑ��'	t2/4h�Lb��{6^i����Ι��`.ؾ/�C�0��u�.�Vw#�HJ�=jJ�����g��-Y&sq_�f��v(��eqO"Ԡ�k+�s�N^��]����[{�Q�勯�)���
�B[�����J
�9��!sEClʮ�/� I5yl7)>�,�Jaa��2���f�G���v�ΗBԖ�/Y7�t\}^Ew���+Ms�#-V㞴I`YdG��](pt@�"`}aww|��{������v���������J�!бsP���q
��h�7�/�$����>(h�u@1�x��d���B'ԊxI��$5LҠT8ݔ$hُ��	Br7����2��N!�? �v�S6�A�㊇z�����L��l������|P��P}��I��<���g�ę�o�~����b���.���i������Xui�Bd(��n�����X�Ш)&Ю�𐹐ln��pt#��%��&��/6�K1���]���fSEe`��Sa��l��Ȅ�\l/�{ ��P�!��ʿ�]=��+~��p�G�)Ũ�Z�\�~��M����3��C��q̻�{6�J��2U^T�$B�pъ�R�T��n�F�eR�����5F���g2ԅ����ma(�q��#� m#f�v�K`SĴ�Tڌ���}�:i_Uc��,���!(H{vc��LGtp/ǎ��&�C�8h+�E�'�ry��)*�M�jTv	�_[�̵�����q�!�n�̰�p)�n���<���$�8U�̀�_ݼQ��T1�����Gq�@�-�j��!�H*�V�I�l�&w|�ع�������)��γ�Y��n��8��1d����%q�䨠}��������s�j�un �fO5ozI���[n��Z�W\Sh�	�D:ls�K����5�D˾��}��*���o���Q᜕o�����ur�7U׷J@�E�gM;�=	`\s�{v��F����ȇ�h�ͤ°L-AE�_�VC�lz�5���O�0���zA���N����؎��� ��`��q~� jM����������e�j��#<GW󳜑`�j���5���3�,������[�]��]�C��
�j��n5/�7]{h�?��pB5�יs�;FF�D����BZ�������_�{K�2P������w#w�8����Z���B�,rw�s ��:}z�x�w��]@+�ߍ����6x�%�8 ��?��C
�\�"��E �l��q��R�Yժ�X�p 5�T�ڮ,�����nc�����O��LoH�en��6�|\$	1�m���{w������>�ޕd"�)�\ �it��$
)�$���0>s�)[����p��SL_�0+��\������(�q�}������ES`w�����Fc�ƌ	G�4��dzԿapx"��u�3!�a�_8�WF)�M�4Q�k �+P>��Ǆ#`�q��\��j�ǰx�W|��	��5�8Y,�N�f�6Qֻ���e�6}k�V4w�T��2�xk-�Bm'�-��D���B!�͠NZ�i�	����_!M�N����XI9�Y�rXW�)"%5l�Ƭx�c����Kj�:�n�<[(F�-Ú�n-�yZw��!���phbF��X��
G~$b��?l��31�!��ߛ�>�I�kn���>?��j��dEt:�D�b���4�M2����Pd�I�h�Yq:�yk�������+��8�sO��-�,����&++���fY��x�O���7u�zAKK�mӖ:�:�<��ً]�>�k�I:�j}Ĵ�;�&�/�Us���'�~��M��u;լ�Z'��h�d�����x���3b"�X@��qN�$#Yr~xO�`晤}��N����<z/pI���g{���PG�����K=����ɡ���PgL�se(
 F�2�L&yt`�fJ��Y�I�5�˫�\u ��܍��!e�ÀI#���%VJ�����b�a΄l�x�5�Ŋ��}�,|G˒����+����U��QR[d�>��5cU&ȥu�}#pWz@�P!���.�G8C?��z�"��T��(S�r-P�k�����,�������4��]�M�H�C5��cꪫ�t6�۶�*RPM@X�B1�1�������2�GF�V��"o:B�=���V?ڣ���_��c������$��si�[T�5�o��G�i�ec�c������"�WE�k�k:TӔ��3fsԮ<V�KG�
�_��@�PK��j*Q;�������x������*R0�w��k��ˍ�Hp뜀!I02�a����*��1�OO�|�FZw/cp�\���o�MS[`��8�������������K��ˏ%�>1B�n�h��r+�Tu��^G�c���zC)�pQ�ܒ;uv�8���������l��f�	g�9O# �tڨ��W��碣у�|Ip���s\�t2	�7�,>�y���-o�^*�=��F|�osh�P���Lޢl��	���<�:���o�\��Zj|}�����廚���K�f�c� 4�]�e��o�'�.y�������r��w��Jؙ37�7^��$҄Lq��\E�la��l����}���A�&g��H����($��b����*�I�V:i�Bk�gX��fK["����.?��.�(<I���؎�]�D�6��*��3�o��T���!�&v��D|��[��u�fI�Ftӡ� �H�iв���pj(�@��f)Z��}��p�Y��G;|#l�݋��5^���!����+ޕn���ML�8���QU��c��