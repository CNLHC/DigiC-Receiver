��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ������
�(5�A�	|���ϝN;���>~}���<����DY����s>���j�tL�KM�`ٖ�t2e�ޱ�*��'��i�����2�b����X�lV+��b�[3�_��`�_߱UF��5��.����5�3��e�BR"������+�����9!6�J���w�W�)Nn����Ԓ�1C 5r�������c����?P�ד�<���;�~c�L�"�K��6�+�'��J���m#E�߻��I��;�Y^�=��;���W��-U�!�OO_��Z�ρLK�o��v���6�T��B�^(.4�+�M�h��TU��Dr�d�91Gۚ+&�k�f��O@�-l�xِ�ME;�H���a^�8b2˝���|t�b�<�7�[�L�N���$�~O��)o�pb7Oj��pg�2���ֈ�HK��*��|p��&Bg�<�,�z�ݢ`X�4J�iIHԂ��}{wUt���g�iD5�l���.�s��7swq�h �A+��s(=^lEū��?�_�� H� TC��ۻB-�H���j-�������9_��b�b�����A��{%� ,� M'(�{U�(�Ɲȯc��e����x+��er~c�B�<��S&^�m4�,f3�X��M������5<�.Ǜ������D�w��� ܜ=�0��~�oeU毜��.�\? ^�.���k;n'=w+S�alaj��_��O9%fHe��玃��[�e�0בig����[ ��L�W1Xs�p�����F�E,9k+)�%S��� �@O�jJ-l�C�R����!���9�~ߵ�7~����R!��Eh�h���L:Vͫej�.]!4�4�u�+�,)C��Y��*�3t�`0;�G�od��^ۡ��@�F�ԭA�N7R���)E� ��)�I������I�()Α��N�O�U��k+�k��ٻ�t�d�"JW��QÃ���!�\�e@��(2 �_��4�� %�o��ـ�Trq� ��y���M¨Mz?%�6so��!�x�}��f�$�C�Z�?Y�U�6�鶬]��d����&�s���'�Q[�P��������aNG��r ���f�a(dӴ���w��C�u�jb�P�I���e2�ٖ~'�;%��@e��b1!�h��Sk�ݭt���k:shn݂Jey�>���>��+n�B�j��nW��b׫���� Ԃ�DEܮȆk9b�aZU1le|Oq�ES��j��	�:w���[X��_��i#�����<�Y��;����_���J~/���^_����c��#���/^~cd�P��.��y���{K5�'���q�p�=l9I�##�Z� ���3#Q	<�p��J�w���l��	M.��f_!�J�m����v�3�t&��?xt��{��k�DO�%t~	��vCg�$b�FtS�6t�ʵ��K�׆]�ʇ��
[�h�ަ
�.H6%��єJjAiԓ�/W�+5��A�f1���`H������ʣ���@Ǳ��5��d;IgkFn��C��H�y��>���\l�2^��7W�jx8�F������;]f�j��8V�0��un�}���%�6���Yo������A�BB�;�5aA�&�
xոJ�d�w�hnWq.���Y-�~���g�8!u_	����ה�`pV��~?DFo�ҁa�10�A���'v�%����U�$����S=�Sg��J(M�	$U}R��=g�2c�yM���8�4O��{��b�7Qhe�r�k�Ӣ*YD�8iƯq��0�e��9�Q`݌�����8�L�T#��E�e���6jG�G�C�:�S>���N5����Bb�̒t#hT�v�d@F��`,��?�ӥ[k�|�|M�9�at*.�DP�����H�l�r� º����
2� ������0=hos��9��ki�Q�AZ�ƛ���,s,�X�I;<�T��3���
`�*f���8G�~���Bي�o��|�c�T.��b�V�� �~��l6����'����{��������q����I�҂���e����Y�C8� ���Nq�L�t����TJ��&1EҐ����m��9��)^����h���6(��=zu�(@��>�ȻW���d0vzl��Ĝ��,�#Q�E�� dQ�"�P�~|�
��?KT�F��}Ъhod��W(Ώ�,\ !��:��i�d�|��(���>�V�ʧ�:�@�h灦Q � aɂ�1����b���.^^C}Ts�����w�D2�|��ğ��/�X꤂Q@��'.Za�3�F�V ��z���x��	x)o3O>�86cط�@.@�hN��_���qA`m<�QG>?Wy1���x���aI���������Fp�JU�����RZZ��/-��]��EYi���)n{/�H�Bq�[�[��v�9����cA��i�����a��If�g,��2n����wCd^"��)S��F�{�Rj��(�e��B� F�c%Z��Oj'��3<:����Y7Ȱ�X4�嫃T�j#Gwf�|#������3)��3�?��d��@4K20���݃ٔט��^��5���Z����c�0��^�� ��;쪻�@5�е����2T��45����W8N�P��U^�h��Ե����9��^�h�E�Q�����E��@�9�ϛ�����m�P"n]��We( �τhI�mu4zp�2L�`}��Ä������VM1���H��d�w�ݵB	��@p���.W
pr���O1*@�Q&\�:�yw�ƭ5[�}�H]v츢 �= 5$J�R�u���lD-�.-"Og..�v&��.�����f6?���"տ��c��v&��n2�W�'�QQ���E�������=��hu�Χ�"p��P���`����.���N�G��A;�`��}�����c�*�R�F@r+����I����S�r�D�F�����N��������(��7tz���=�n�#��E]�1];�Ǐ��8c�z2S�)�~s�I)�t��hUX���V
	<�*3gh+��\K�˰�<��`�b�/�2��(4.e{2�S�i�,��	Fi�)�BP�.��,���]�B�acg��Dn�H��>GoS�6!U�M&~K���pjq=��賎�yL`;��N� d�W��s�����s�޶�3_=D���W'XUW��_�2�/��a�QlWKY0�-��&[#[^$��4��Zp�i(�]1�3�rC���X�	RoŽ, %�;%�G�J���+�Hekݲ]��h�Ѕt\)��,m���7�~��Lk_e��򇲫��\��8�N렗°��0w)Du�7��F�7r��7	��	L1�Qx����Վ��Vߖ���6�R�t��Dr�-��� �~�v����jPƙ�jFU�nm<�;E�+N���4.�������+��=Xƭ_��*A!
�wy��P(VS�W���Mr��,2i�y��'Gf��t�g�}�a���3��3�W?-��Do������nZX<-ړ.��QR�[|,��0a)~3�5
�mr���7��Y���^ۋ�����i�P��N�ǂ���}��O�GG�-�gA�D��X�bљ3y�k2��b�;ﻬ�D��e='��ܳP�����C��Co���~k��<��&T@U�Q�W�)dJk�J�����ˑ�3�����5��~o�qB6c��&+vԿ}����vMK?e^pʰ��	��pUQ��T�����Yv�ʔ)�%�/N�n��r]�S��N��}l�ӽ!�:��Nz��?�h9v&r����({���?Y�E��3�m������RP�9����2�)�'�v�j�[$u�݂��4�'F����5H���x�����4k���]?	���(sMV�~��(��M"��4��7����0� ��[x6`�֤2&O�<�왆���i��*��Fxx�E�Ab���mw�_ш�i<��ɿ��Y!��v�[�'�©׌=T��3������=�l�r����r����@�����jb��g�hY��1>��F`~��߀߈v�rՔ����IE;��]�lѼs���*ZE��5��V�p�a�����ƁzA�<��%ZE����k+�>甃�[��I��$5�p���qF�VP�4V�=?��t���t-uYR�D�"�ыWk���^�1��������Eן؋DǷ^gH�\�+�h�F�V���zv�B ̹w�odv�A7U o���ac�@C�z�&jNL�~,l�����"D�ˋO�����y�Q1r��z�9�&�ھ�*���*��{QiWKm}-�6s��-���0�UC���H'�G�� ��wƻ����x�"; ��Ej�,bd9A�YL�M����9�CLQ@T�n��3�5>*kV��gd�-�nM\c$[ʬ�=��r�\�@�H�O���jw��:	��*i�Z�-���U�pz_B�P�B�#�=&삚�W��g��l���H���e5�b���>m�4f$�� ���Bfs�o5�P���{m�p���;����|�.}d�4��)����h#��J���EN���T��5!d�a��id �WP�
�"=��V;�&4,��jTZhY/�/M��ٰ�OK߃��w�T�����&�O6[i��>�)�TJ��S_VK���X�/|��_P�+;4�[�6�^,V�o� Lި<����;!~{Ɨ�����I]AZ��v� ��h�.B�R�2��
4p�Rͺ�!H^t���Լ���aC��������{8p�V�W7'_�H����LRO�m� ���I��?��ʁ ω�Vc[I��NE�j��5�Y.F�7��Ň2n�&�%MY�%?=fTw��MLJ��|vD���F+��r���Y��8�Hq���!��(_�;A����\��q6��ND�Z�A��II׶a�9�Q�1��_r�@�I4�&X�1��޽�5θ�w�E���6t�d��!��dt9�D�����,s��G�t�ⴝ:S�mi["ⵣ}M��_����T>����M�i{�[%ߥ@
"|?X].҈+�Ćy昔�Q#�������X�釄xƿ�Ii�Ǜ�cɛKVn�|�j�Eρ��<ƽ~�����r�;	ަ��9��#��)�UHu���\�4D뙱�VQI��|��X?+?B�iգ������i"�D���V�8o�5-�=�B�x���q(꣒��/�yo�M�?�?]w��	�<}FU��`�Q ���F>m�;8!��ԇ�dS�HUlDC������ ����k?C�~��� ^QZ���Ȧ_��Q��C��0�n�eσ4Y�'ӗ��ŋ�M� 2��c#u��!�Cc�1� +?U�}R����Ǳb>d�/�ƍ����(!��_���'��Vf�������zm�x�(1),�A��h��:�=��CA\�M9譩`c>55h/�.!sK��r������������C���a�M%��[�8��-�%3Jn%���޸��)mzt��<�%�[�my������ �A��{�ݣ���᧼��n����z؉���f�\vv4�.��-b�Ȃ/��_�*��l_� �R�1'�<�L�6ǕH��NÙ���
<�0��8�%5}��d�u�e�%�5�0}X14G4�+[?���s�~��w�y�A�/��Ͱ]j�)��S�>ɿ�2A� #W-kk��Nڼ�l��`%�m�d��\�[��F1�������]O��#J�t�5U��]��^n~�\�"��hhP+a]�:y�l}I�ˢ6�맬�,&� ������o����E�N.�}.Z�_mhM��ņ�w�O�=Qe|�E���"���O	��S}k~\-?���Z���J��������X�3�HDO�#t�o>�׽�ف����
�R�.�����8:�>�r�3r�Ӎ i�o50�#
����X4��W�O�s��#���Ē��T�V0^���d3}f���١��4��.��i���Ҡ�3����>0��F�q�(5�M����g��2�l�?]�N�
�5Ω�O�ԃ��C]�^y�%�d��~͕س?\�v�Z�LjS���rY�=��U�4?>���1K>��y�N�)u
�1Z4Z�n���}��ۃJ�#L�Gu�7���s6���vo7�وb�yg$���'��L��Q,�V>q�&7kB��lǁ��U�N�?­�̖���+�e�늫�p#$��rb�'�z�ц%�""��EC˚��h~�	�)���n����X��TiX���ˍ RU�G�F�`dc��љ�'�z1��1��V֨���ā��������apEc՜�Ged�ܡ1������CU2��!�	^�"����Kg�m;��fק~aMn�/
���$��!�H��#K�u�3����[��6A�Sz%"�$eZyOc�Ų���~/{c`�cx�q5�z��l��-��L�����m%3��l�B8��=ɢtI �@W���h�x?����w���O�Jpb�d�)���1bO\���ԟ��z�J��l��{�P1�������o}<����Q���h�=���w!_�s����t���ic�(�S�^Bis���N�"VU��F�yl�m2�/=T��\�J�Q�R֖`���n3�j�a��BMp���@Þ����Zٝ$[�q���"BC�
tJ����H4яE�*π0����3�h�l�0p��Ζd�O��zD3�̟.b���u��`�w��dS� �����bcv��v�J���iѐ�	Ch�֨���>Ȓa�&,x�8�b���Ia忻��@��+�T���\����:-��2Is#�\��������C�4�)��MME�O�Ҹ\{S�8:Ǹ�|�t��Y�֋k����li�yƖ�&]�I��o-��K9r�k���j��-�|������Sz�2�͹Hޣ��3��-���W>_l!j�M����B�7���̆b���s�>��K��
�;g�����]�Ӕ��SƑ]�[!É�c�`3�a�XO{[^Nl�!��Y�DJ�Cd�.�]ը^�p�U����*�HL�/#��P}x���q-8-	z�^b� �ӽ���.�����,�"�es��B�J�`��=5���,�Moh�j�I����-�)�j�_ {�43I���e=t�%ɰ�i�c"�l���\�h�8�Ï3^�y�zs��k2u G�|��^-ZlRS��g5_�9�ˤ���CH�cܼ�6�t�)�o�8�Iw��xZB���m���{��!XP=�i3�w�r3��&{����@�q�qlyj��0�/*�Ԁ<@�t_Y9F2@O�&�9�M��B�]��#��H~�3��g\D��!}�vf�=�"�r��CI�.���d5�!f�>�9(�&T!�fL���f��B�yg��gp�-4��,�yy'q�����i�ۡD�R1�\ja�3x�Z�v4s�&�Q��Z�ш���	gZ�Z���ѬxƋh��R&Z� �����t��n��VO#؏����{-6	��.s���+�oۛ�ZD����kȿ�>����!�pn@���Z.\@ �B�v	�e������������Hc��gS����J�L v!��	u��gfҀ;r7U�(iYEWۡ���wo�LԂaDl��F�>��T)�J;��#�.��_�8���C�}\��9t`CfA~A�u6�HI�s��%�?/]
i���-� ����	4���,�I9��q=(�b&G�j>��*���q���O���cE87lmw0
��Q��O�w7�_v�`�);m8IC��B3^�B���d$�S���y�
����M�>Iv�tm���%;tb�% g�&�����D?)U-�@�(��ZIIB�ڟ-����I��۟iY^X�p���Âo�3��OW��+�����V�*Vk�jE�?�oLwJ���yG� �؞.$���Pn���l=�'��bR<�v���6�^�{Ì��yND3�	�#��=�Ɍ�/b} ,��\̥۶\�9��I�g�Y-:�&,�f'%�f�2G�93g	��;�!��79�#�9��q��mc���
p ��=vY�~�E;�I�2ڜ����� �Lz�\��{Y$�;2��ۓ�������iXD�ܸ�����`�%d�hi4�YC .�v� 8~�H��Lݤ��!��$��m۠�K�Nb��Y��d��M]���j5���g%Z��N1�E?����d”�"o�SV!�>Y�h�w��x?�)�
������V�`�J�p��\�¡�� ӉW�=��BQ^�o��L���.r?�;Hj��_�L�Ʌs��(fnӎ��~������7���&�Z��t+
=4G�§Bϯ�F_�_v�.��њ�����%�%&W�/@j�dV#:Hʰ�bE�SI�v�<�h������߯
�V�����g:��@��J��B9m��Ѻ�q��p�g͉+F[J��P���oAH���.�TE5�k����^����ɚ�Ә�;�:\r��Z}c}���/s�˿�NO逧�.�vG[��RٖS�ņ��kW�:=K�qP����fkӰo� ���V~6��Gt�SZ���-����y�?�0��Z�<-l���ʰ�)+0�d�+�fdp�J�Yh�A�xC�m�i��a�^����ש2S���˳�;��4��7�刀19)���?��ʹ!����=g;��v}�0|@�)��튃���J&B9��m�A]ۚQ^u�g�f�
8��"���֚a��h�#����gtm]�����ew�2���D�چL��
�eG1���