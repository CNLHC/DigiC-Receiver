��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]i��n��R|�u�2�vi܏��Ns���5�ؔ���O	��A2��Ap��:٥Q\d���y��> �<�?�	�n����"L@��}�w_�b)Kq�����k|��c�`�:d�R\S��t�h���r1�%��ap���*?$Ȗ��쪜}֑hw"�x����~N\u�����7�k�$����brJ�"��^��><�)��E�Kw�w�n����JȒD�z��������ZӺ^貱��ء��j��>�l���b��U�	��}@ ��D��w'�O�������擻6�7/���[Nf�S6,��H���T́�d��+
��¥W���r_=�`�	"����¼�8SSZr�ŭB}9�
�������M���MKL���{DL;�U���%7\ӕw�ZZ�S��'/��d�52������f���j���6�b�ݲ��hP�s��i%C&�k�����$�C�t��A&
@w���O֍y{���Zb���=6O��;���><��rHY.����κ����N	��D�z턾|(�۸�2�*�R�I�E=G���m�0��a慵�����bjPbd����)�?�Ш�8����6��J���ϊ%`?#�U�KY+�)�o`��)�gկ#�8�ЅI{i��F��5�P �{!;l�m��(�W3V�%�]4�#���4v��I�pa�a�|vS{#9�Ҋ��|���#�N�����\���B!���M��.��j!��i�N�\�?|�ܓ���F����$Zh�]���>��8Gn�y�?U��_fk�HN!d�cO4��g#䷶X����ZP��>t��l���v�y_{�wե�!����4^rVo��m�G��x���g��Hby�s�"�5�$/W��>�i�{'+��4˖ .#�o���z��}��hz��%9ԁp�n�$K��_���K�F��*rl�d��u��)��ئ���o�����a_|��|va���p���:p0�u�;]W���?=x3.��+VO.,$�D)+`�݊w���'7k3Ý�L�5v�[�l���t9�ne�>/��$�I-����� ǣK'�vb��yI�eC���g����6��郜�L�8�q��r���N~�p�3^��UT�:�6�*��P���7k�̈́!oR�$� $�JZ��[��h3����8�-8��@����&��dw^�]߳�^�_
�g>�/�`�%�--X����Rރ3�2[®�=��n:���,�k"�2y�Z#'`�3#2C&��b�k��l�v��l� �ho|��j�F5hv����"��DW�b:���w�HMfϟa��vv/��D���Fݠ�$�	�k����"AP��P��pK�������g �Ꭻ#[�)��}3ӡo=�c�~�y���)Qzԯ_��S�`t_�
8�E6L��N��p�j���ʅ<�FM �,A��@p��܀�����I�������Nhh39ߋ�~�M��Ɗk���}7��>"�7����%� ���}
0T���-�����k����=^c�6\)~El��y6i2�.�i�U���Qb�ǝ�~&���rA]�]��Ț%�n�?�m��Ϊ�l%�G��d4�]�pU�o�L@���ؙݒK��7CND�E2X�?]>�jv�*
�O,ck��e���J,s�S�O��r�dn�`���o�\K�9&XJ�k �4�!�{���
�_�	%�/��l��CR� ;@�����u,��9�����w�&��E�3����ғ�dhp��d;kX֮:����=&1�[��se%��N=Ǔ|j�������T#���㲘0��*�G�Cr0�io���[�s[�B�Yv3�яڛ����ëX�V$�O���/uz�x����#��"��`$����O��N�A"���Ø
P�el��Ǆc�J�,�a�7���o��R� �R'Q׊/��0����̮%hx��%���s�ye��]�c��<�6h����z�"��Y9�Y�Q��U�7�4++=y-��3Oc8ٜ0����a���f	�<n�=�U��Q���B��6�q�����7}�x�[M!Ċ.N�R�h�Z�	o�	:Uר�d�_e���^����|�1N�u�x�ph���^
g�p��`4����)yb��5��֓����~�:��>�e'MG?dt���4���J'>MQ"S!)��uR��A��Ԧ�Ss�FQw����i�ј�+:�Nd�b�9��G�^��)��:Í@(�R����*ĪQ�[����m�
&~�����L7����b":o�29K{|�׬3�ُ/�6�1$F<��ٶW�)�b��d$.���g�Y@�P��k:1�w���b�֘�d��Ӡؔ��?��U�4sɑ�?�*�`��+G}�Rj��]�`�$_n1�7<��p�4�7b�ZR��*�*q�;����qI���/��}TR�=B���n>?�d.��X�$�.�Su��N�Vg�BI�bK^ �|�C��q�&0u�o�z_^i}
��Ӹw�M���W&�jI��;U���oj =+��N��������ì�� }��}��Dc���5ش$(��<(#v�yOׅ��raM,� ]�=&f����٘{��s�m�1�+�F)0���N��ʯel���s�8$��J�����@�1����j