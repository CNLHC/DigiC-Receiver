��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ����u�SM{�"�Z����s��`K_W�]L���KLv{�- �-��]��k8*Ƽ�Ruʖ�!l�Y�^9k`O�����Et Q"H����mFf'$iB��k�ۨ�]�� d,���>�������7!仔qN�Ɉ.��WWrU��:���|�rY��E���ڠmyB��<P��R���P1����LۍH7�#�u����;:���G���{o��w�m���9~$���D���g���rH��SA$�Z�N��2]Ѵb,�e�6�G�0�H���A����;����a���L-�X�9uL���fR,Ӏ�_9ϵ{:;۳��n�6cQǵ��ڲ���k!<P�Z���FT��%]���ru�}1bƹ�(�ͺx�y�{6��G�d�<i1�� �K�{�m ���9���yz'nVڿ�w�p#�{*�����[�Q�ԝu� � ]�9��B�e����{�:4ʚ`m�d��|j�C�����W�s�6��	�^��R�u�e��lL\D�D��y��s�?	Of�Tht%�������4�+ۏ�.9A.pE8 ���DH�F-P�l�'Y�<�Q�y��9�Y����d������Q��x��Z�QP�K)Ǌ%�F�?�
���i��>��F�w�8�c�۔>�`�>ę�(����	 gm�=JOW�L��{��ue�g"E��,��u�N4���� �mpYp	kv���E�S�%���j:��M��<�ղ��>i��ċ�@}P�����	�SE?�ѵ��4�(2(6��B��e�$`伈^ۻ�&F��&��fH��'j�n}<_ux>����`�߫��g)��<��,��7�o�V�\L�0�i��t�+�J�6t׏F>��?�HL�6v�4ҏ�~�R�O�����vl`f;�c+��z�}+n�f7፿EZhf��N���62�"97��_�y�٥�~NR���ex�C��8}~�H���j����;�4Z6�����s���;E���y���=�o���%ՆZ�p��DJ��[��6�U;�V
l=K�h��3��»�Y^��Z�*��'ay�aM@���"�A�E�2�����:�J�v;-�	�ܼ�5u��F��c�� s�3�"��Z,N�j4PfY$�Fn2z={'0�j���4�O!97�3d��Z�+D5b�D�����J7Jk�Rƹ(Q��U�O�5���<�X�%��~5q�����R�JYp1D��f���9��
vCOG���Г~�J�PM@ ���M�#,�4�*�;��vh�z�U�{�:��Ն(�*!P�2�/�Re¡����JA]H�[�4Xx����z���-�f].��Y��C}FӢ9ϭj���;��)d�ב*U	r7������`0�
��Wٓ&�ط�m[Sul=�hp�Z����p�&�\NH�4�{ <�H����[���*ӕ�z���C0�F�=�TE ��a��������!��(��Z��ɼ�������"�'vXl��R�`%����E�x^��}�b[Υ<<ۆ��R�t��!�_O�m��+^2f�R8 �UP?Vu��N�����Q��xŰj���k����cQUo�(�a6SC��r��9Ք�ݱ�2@V�b���~�4��L}l��p@�G_?&>e���\��-�������P��#���pf-˂S-f�ٔI7Q�a[���?��A��D�}�.��l�P��u4V!�S=H���3���[Ar���W��T5Q�j��F9��\8�3MH�b���~��g�u�2�gջ�Y4�̥G����E���nW�r�G�`5bG�ċM������N����7.�xT���_�/�	"o�l?8"��/7���I�{!�;����+,���gxn�3,��2>B���*5���%�ש�ʔ�����ټϦ�t5H��⅔�;��E������.� +7��Ɉ��D�cۅ�.m�f�m���EG��H���Y���po�v�S�S�ܖ��:ʋX�&�����l���t�-q@�h�LCÂ��?�����N�����0�gR�h��6uP�� ���ɪ�<x*�y;��5r�_챍��,��$%C=��>O?4��-Er<Y})�s�����3�m�Y�
x�^'��8%��˼6�sL�m�����ɥ>F�ƣ������D�py���?�$KlVi[6�!�t�]~�0��Z��H�,����&s�
��Ww����^�ڊOh���P���VT�z�������:�"�`��m�.2nנ3�4n��f�����4�?�:��s��9%�}�\�w�3B�X Μ��e�?�����P�fJ)����kf
��*\^�ܼ�^�Qb棝�m&�����T>T�f��t�X?b5qd��Y	s��G3 �$�Ndkm���9���ȏ<Ѓ%���\�)j��m���V_�yn�j��L�θg3J�4A֩��#U�tdƀ.���C�5*kQ�"�+-���?��K�f�c���3]QZّ�ߵ�����WX֞�T�$���S�ǧ�����|p	4Qգ������1�U�3C����:�s"�X�\O�R?�G}u����4JZ.���+z�Ӿ�!��2lR�`��B���7�a$����1=�$��q����c��P�`�گI<7�%�C��Zx��l�Fq�AQ�=C[�7���4��'�`�\��$3\/�aC������h���f�*T$CEF��
64�tҐ��U�*��!)��v4A���\�}k�͂��&4-�6h���T0��)�OZ��#ŵKO��ٱ9�^j��
f�8��SW��O�)�o*thB�A�@3>���J���<�9��Ҁ����򛼌H����7,d�,��x_̪ڴ�Ѧ�Q�qޒmC��()�nɚ�v\U�8!�G��GJܴ��L �x�F�(t���U:�jPe�L����e�,���#ҙ�3�����So�.l�v\Mb�,^<E����(�c�(��g1d���(�﯈G����ԥc�(?�1�٤��ע=���Pu���d4w`S�s��f"�T�h}9������X!����{	I���K"�:�E�H7Q�BN�e��-�b����^�-�^��1*��Ϋ@KB��a[�:�6�9��EY�,`�m�u �0i������r�:�!�����׎R=�3�`�J
���2,s�F����+I�m���Sj���}�2�.��e'm�Ӭ�|�ϝ&%�� ��5��!�`��@{��SYִn�m*�I�mf���ħ|7$�Q,5Q�UqִC��Q+�b`������C�
���4�5c��k�H��|y�5��?FJr��D��c�P�� �%Ql�:�sXΥ�Ҿ�^R��uM8x`[�>Mϒ3�Y���z�nH���}��R�U������&�s����κ�0z}Y��.�!dC�q%��Q�xn|���Qew��n��(`���yZ�b��n�ߺE�����U�uL1���m�	L�_ʰ-YN��s���
�Ok��ndŽC7���Zn�Z��>�l��i�߸��_<
jrrz�.Oxٶtr�Ke���G�K���T��.c�r�C����ɦ�yl�DS�f�1B꘧w�9���/'Z����\���+9���r���"���_�oON�����S����iu���	[V��И��Yg�A����%�����(`�ɓlBE.n�`�
L.�ĳK�&*�SO��(�O�Ҿf��R�%��%����"Z�넨�x��m�L��u�4mZ�&�X��OCl��c5,0�_��36�{���ҸA��?��R�C��ڣu�8*�aWB�R�o��~~����b��|o`�|fL��;��}[\v��W|�?����*�"M�@7�[��iNr��
�P��/&��kIk��S��;�䦸t=k���(v2��e?����?����Ɩ,!֯�� 7t*7��53|nj*:�XL!�������"��%{����"%F�R�ͭ��ę���þ*ۡXE~Q�cF키��5�A�����Ao�eB<��������TR*��c��аЂ��)$%U�{<!)DZ�Y��s?�Ri%���L_I�-_NÙ��_6O�e$���m	�k��7���Z���14OŇf�ce*o��%]�u�*�kLfДk�w�J���Uk���z��⥥]��$6�d���Wf@CQ{t���"�΢����@0YE��g3ƽh��:��rYJ�� _2�T�����.N�(�'Q��B48HJ���݋���hǼ�W}�[�k4��\,1��d$5�Yz2=�U����~mu�ƛ��h]����=����/��/����mw�kg�<���-E�
��r��R�7;�]Q�蚐���%ؼ?C�bJ���@K'�v�&��F��}J�����ȓ��|�(13�i-J�����'7p
����\ ��I��F\B�$O�=���
�A��/WP���\�%U��}�ة0wn���2Æg6���#������(�&E�5�M;&�H�CX"v�n)���@��8[!&o����/���A(u�c�I�����5����FzV�eZY�
���V�A��?x�I�t�a<]��!��6���_���YN�g����7�[˹�������j �u����7��:��p�X�v{�K?�`m�SބvG��̂!��Z�8џ{k�B4�Q�,'uk!�R��aUǗ��gh4Γ���t�z��``�cZo�9f3��l@���R(���`dB��#3�5ft�;bs
=^5Y�X����	�l�Z�8~��S�wmvp.��\�ʳ&�!�`7t�0��G�����K�{��w��^8$��AE��*�wŻ����3�=��iT����ү�V,�mYy�$~f��7��݉�%��R��'|*��^:wbɛ���*\�I��J2߃;p��8����Ż@���7��'����+����l�6�:�\w�p��jz�Η�B?�H(�nnX{'˒��`x��f���5�� �k�W���.4���������!�X��莐����E�2�^ֽ�4���*H�Qn�� ����G����D&T�J�%�=<월E�*Z7��������Y�Ͱ��7ZzԒ4�����ӂ#�K�2 �B%P�+�rD$���o,v�_J