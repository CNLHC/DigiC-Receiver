��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���������V�ċR��u�z����;wjH�"k*��� ��������eA��^d��UP�/O�OɁ�L7�i�lW���pJ4�}����N{,��L���>�e�T��j+LW���Z�z�ڄ!;#����a�1�S�g�����H=7D�22��Ԟm\��y�d�S��X57��Y��^t��&�X�P��)-�`��EX��.&��q��T�����ӏ�2k�����>�M]�&ش�{��]���A'(�W�v��sS�e����3��2I�V��>��_ �[��<ń6y�$h�u�/Q�=��!d}��L�֙>_�M�;�FQۀHߍ{f0�T�:�ؘ�W�΢����9P�����>{�������G���� ��D�����p�F=_Xd��sH�Ve�߹�&N�p؞�@���7J��:�Q11H�z�z�!�fɣ��̸E2'o�_��s/Ƴ3����a�]/�p�B=��J�mOM	ld���,V���t��҄B1�|�2�<����ـ�oC�(�*VݬaƶHf���hS�gJJd��g��{ӿ&��oٕ�jn�#����!�<\4�3U���u�{}�vL�Y#�_����
B6i���;܃�k��`��@~QU���Əq�T:Ř����v�wV��Cy�d����/B�b�uA�NUg�R@�����KJw�np�E������55K���}0������5W"u<��"+if�Z� #���t�M���/��_�Q��Jb*ة^����ł��,!.L��}	��v)Un�wTQB��gC�R��&�fV�ӹ���V�-����4ע��+#�"��ҡ�o+�3��쌹�~��/q*�[}����}���������P�����d���&�o- �(�\�ڧ�˄B5����s����ud�8-3�i��Y�)�O``���h�6��E���*���N��T;�q���u��qxt'Jj�
!���������>2�N�:���՚�zĈ$�$�/Ǳ���{�*�%��N8e:5ǻ�-*mI���=�R�#���R��Jt�^̜��>������4��Iu[��|~��,�u8� ��7K0������j�.MT@����dDWDC20�;.�p9�s�������='�{�������w��`
���eA��Ji��c8�2t�cmt9�Y�wڷ��O;ːnh�!��Q�[Rb������|Ǉ;�n���yk:!�W������<�ث��2�5����%�X-I2�ƹ+h�.��-��LD�#�$�p:�2�(������x�	��a�T�F���&���#��s��� �=_P��G�4�R\�'
���Jv��#=!d�QIb�	
]Mót�m�%�rd��f��7n>!�e�7ڧ$@�
�N`�u�����ci�=܁(��[�߾��F�/6m�s�	-�"��w7A=�i7�t:G7$��u��#�;}?��Y��T�զ��ve�KC�S��7���Z�'�fxܾ�B��� ��Xm��k-?�)��٥@��m���6a�]�(��.�{ص�4���?w��I���
�97����4���j��4 Zl�BF��;��L�2K��� �m=�j�\�)c��|9�� ag?skxRi��"��M0�N�h8ᵠ9�44-	�?��cY8�l���V���d�\q�'��1O���ҔK�m�,��6�$�	�H�z�u2�����ߨ����s��^F`Ly��P�+�D�m~}����UkЅ�k/��j�<\��T�י �K2IF*��!���x��P��A"k~����jh�f�����+%�uQ�6�:ɉ������j�Z(��h�ǒ^��<Q�Q#�7��R{�3��O�5}�5�LV�������v�ɉ�>��Nz�����s���"""d� �&M�FDs<�F}��e4I.r�:���0�I��L(Z�ӊ�/�'5-�I�k�&	���(�IӲ���q�V�� ��ڃ��zk��|�A8]�Y,?<�*���Mc1КR�����#�_� V���N����6bu���������6,��R[
\"P�c��o)�M�j����r��V��0�_S���=w_��ls��Ƿ���b���\%�	N�4`,J��O1$tB��!,��0k��3�(�kDW,�Ć��}�Bx}�S`�mQm��ڠ�, &��cj����e�ӊ�#��y�b���,��0P8�m�f��P�`�\G�� ��8�2�����W�]�S�[��$^�'Ta���H���.m?�"�n"��*�M�U���\���R�����n�r� ���G2��8��5$��&��&$/�)k�{�.��� m^<%�9��-�9��A�W�P�A*���=%�J��/>ɷ�3AA}����4,�k�kj�o*�nH�y/B�0q�f��VC.�)��5��߉��3�?*f��	T0ϟer<��8����V�`BL
B��Y��ٱ @�Y�/�E��4]f/�.���a���U�0yt��D�6��@>&��깕��zѼ������|��gI���yV��p?��mn���<;)]����`j��b���._�R���l@�κ�;|a�l!���u��}��"=��V]���_�T���N� x����C5�?����,��a����)����)�	���U�l�Ϡ���Pk�Sx�зp��<!;����4s�r:��?���m4$˕<`��'uq$Ͳ�H|��X�QSyE��QR�qll�4ɈMD��n�"���:���sl����6�oD���g�!�fԳK����	�(]���ka�'���X^�"q�$A����{�$��P�1rZ�ZedL�A���� ��/����3��$����v�˯���_ECn�2>�r�ȼWk
&��U���\�4�J��D��~����js�!ޥcRׂ���J��J����نfˇ��6��M>�`�3��z��yV6&צROﮇ���9a?+�����BQwe�1����=e� ���:l������U��/��Fo?��H�fɳ�Ep�H�Ɋ^����[����r�ki���xߖ��z��e�6����Bw;�r��Mw蹇�S):�a��d\��w5�M��ץ�e7�۩˝�n�p��E*�0�&���O�C��X�`ر(w�����7Ҏ���A*g1�$v�'�lȄ��鋃�Xm��4?���L+��1M�!���o�4;r��x�(dlm�W���l�g ��jm�f��[1ԝ����݌��Ħ���K���T�k��됨����j8�jqHŤ�ƒ�4�G�yR�)�|�̾���g�)gA��[<���tLg��ia{h	l�wKٕ��/�Df��.��^)�d�&W�5R�/��]���n���(t��c[���2=s/�K?����q�5x��h"?��@���_��s��9^u��v18��V e�V9��5�'���Q�A�9�\{uyJ5j�����G�S����6�^�B�}ކw�9���>��|��d��W�1�@�1M�V���/�Y|E.Ύ��f�'	��Co	(gn1�gC`��x&�k��X.�F���ڬ����k���Q%,Xo�Q�aOix�_�����}r�(�iB_�e��7�8������2�h�s�&?l�H�u!2�RI��>�8c�Yr
H�!']�W�Fh�I ��$2/�����z-x��^�� v�g�-J�X�qv�u mZ�tT�b}\�ϔ���WYL�1xYV7��P�Ù5��Т��4�ä��s�>y����;���b}3P��p35�í�D�~��ӷ���U6Y����tw��W�� c%��G��"�hC���}��<vhR���*�������]\���)CwL*~��sƘ�a���LwE���i_�T�v�)��>0�qǗao�nd���?5��(�'��n��4}��Y}���>"ᒦ���n!l�E�<ے��L�����^�]O�n��Ƶ��6]�d&:��m�Wކ*ݘ�p!���5��Q4m������\�k���FQ�}���_�`�?���%NS"~�W�S"[�3����̸Ѕ�oV�?���H�!ҵ�I�.Y p֌�0G��: Z����zeG"*"[ϒ{��"�S0�����=S�(2�R>��i+���z�@3�t
-��� �����_��Nq�8ٚ~��՜��b��E����s��]�P��h"�2S:�v�˒=���!?�f�C�7����*��ᰣ�?y�v.�d����AF)b"�+��a��_�����Ŏ'�&���u�V��B��Me	�׮��t�A���ZB��gc/&��/򗢉k-�5e���		KsuZ��I��v���ӟ2*T�%U�v	��w9)%�$�$`*	�h&��ׯ�A����muc�m���pz���ș�:&��ߟ:Ʉ�a��$=�Dkx��x�A�݅�
��*gղ����Xsv9�ۊzɧsf%ľ9����X�*
(��W姂���n�7z�	��}�Fz\MZ�v���"H��4l2:Y��!0gQY��"q{�SO��I���t��X��������|2���m Y���5�$f��t	鸤�����lXi8��>�#����$&�:��p/�Ш�v�U��A|���X��I�,]F�H&q���FR�寁�o�3��8�9w���Ĝ:�mXCZ�`�=�4���i����0�*�Kƹ��ऱ���1uH=�/H#՜�MC�f���u�ɲ�@H=nz�!8�����yq}��� ��5AP�2��fl5=]F4�;B ���LU,f�@-܊̺B6�8�d����/���t,�(��g?�������:�"�vr�R׌Ě���6��;��k��z��7I3F8�֘O��.��/t	w�pX"6�ZG��2m�7���5\'C�JԢ���ʑݚ�	u����rt=�_(K��>���_�s�_�Q��ÙM�?}8yu,O�N+�<���:C,�$_�]O@�����1>L�@1E��^���HX7A�v�}��ڰ҈����L|r��vr��%���oovkz���H�}�0�;�Ц�"� ^xRV3�zd�v�����5��!�-�9�k~Cƭ��<)�$Ȣ�l���R�9�4q���,�$'�Wo�1>Cn���Hw��&ꢌ�\̳J��w[�V%T���6����Ω]���� >�nNRġw2��ɭ���E�<+7�gx�����Fa\�B��r���{nk�$���G���hY�5W�K�%�	����a5X@V����5��=֑.U�0�0⩏muŁf} ��M?ٗ��Y��rK
��H�ʮ(ꩣ��W��7.5������ZͲ�l�iP��5WRJJ��
'A�D�ށ-~��}p���Y���%��=F�ŷ��ſ���Y���BB��	F�\�80YZP�m �����7����������k�֍%w�>����o_�_Mb����d{�lT�����m-x�ZA��W�1��Y�~A2�/���Y�$�t�����L�I`�ɝ΍M_���N�d����4�b[�"K鹅�C��u
�9G{��	=i���CG����;�t�AE���5I���D,�GsY�pd"s>��z77��ޏ��`� 0(�	�=	h �xѠ~G3�*)x{�xч�X���Jw����+r,Y��u�o�XYЛ>��-x�-��D�	l�_����%w�g���'��IW�e'vRI�GR��@}\P�Q���J��ؑ?:T1��ٴ�K���{(8��u�DL�G2C�1A|� �~$k�h���$�e�_���P��M��a�)�č��1.�����mV&L��M�ښ��Of6��;�c��2����[P�Ff�X#�(Ҳ_��ztT����_0������j���Gt��<z�!c��Л��Cy�uLx����[-��A5��I\Yڻ⠤�L�=�7F�?Ϙy��|ݡy�4�2!"]#9AmĎ�<Âr�u����F��Gq�T7a��3&�,�ҝ���W�f�2s4��0�k|�Nt,fE��WQ-r:4�=n;�Ҕq�8NV6��.��0�i��<&�"O�>r�CNd	��n��F�B�Q��^�v�9g�Bz�s�E�ڢ�o��wxhJ"G�= �\U�,x.CU�v����qj.!��J6��֖���@J���,D�P�N���b���~BDp	tpNN�)fD|AD�����Q���ۖ���N7��7~ڝW�P&j��t�,�e���i�������s%ό q�<, - �X�""��zD��Sc����h�M�R�
����Yį��ʉ*ܮ��,�J�wx�"�������z�W�����=���i?N1�g7o�_2�j���?� 4�䕇����R�zZ�V����L�\�}��G�
W���c���.�25z�2p��m�r�$�x�.*�lgłegخ
�B:�̉�_��v���H
Q6��D�y�2%d�Ia�$ �*u1%�W%+U���8��ه�;H��,�o6ꍮ�w##FY�e&��K���r��<�+'���.��^�P���:;9?1������I���S�Egj��),��mU���I�����H�� <��:�7��]\v� �:��d�x7r���"z]��땙��$��z_���l����giO ��D	)g��V�Q��坉��y�ޥNӿ1�-͙�m�V
ҏ ��i�f�5}�P?�x���%u�*�0�=I��]��N�Ղ��XTr+�S�=�	�kq9}���7L�c��G������-:3��䗛���?B㛅�`�7�0ME_}� Y�T�a��_��Q:�>5�ľS�!���Ԗ�i�-�o?�~�=�<�r�z����D�E�@���m��܉6{�{��G|�3:��ʦ�S��܇�|�ez�W۵EpS�1A/`�UU�����?�_�E $"�Ä��.� �����Z�.x6�����Q*$�i�S���ܵ�� �8��	�/N��4�,����y�XeSO/�nNSs{�5t��$y	����i���o��c5��z��zϹ��%�MU���<��ё,�������]�Sb2�s�v��b�������@�Ғ�l:�~$Dg���e�YX������\��.���<zG��}�����ՠ�o3��39#�~h���'��X����~���mt���Q\�HI��g�d�h�'��ǫ���$��s�V�!W�smH�I��y�_�Mys�o�.�6�g��������`���₝��~A�	����^e@������q]&���e͗�X�>m�}{Q+������u�I�J����s$O����_�p)H���!���i<V��"9�~)����O<�ZM�K���qNYYbhU4Hm�s?8��j-	�R�RN'�<_��y6��(D�q�6�,rp�e��dM�E��*4-޺���r$ hQ�z���*�>G������E��˵���l�n.<��z=M�T�j�T������
f�&|�x�!9�� CI�v��.�\��#H���yl+�謉����ע�!D΃���l��5��w�ݨ��M������}�;���`"ev7皇l�x�q]�ǧ�о�
�� 3C�*Ň�*�&#����mH�oF�)�A�1�
�Q���DJ؉.ֺ�V�͆?�%rSV2ߡ�"?��}�/��S�