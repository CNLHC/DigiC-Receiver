��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]���-�p^8�3 ��TLM��q�"��z�����`%F�zU��K�^��3��}]��0N���������E|�+{��O�z��Y�%��l�d�f�����M@'VX��%�����F�\Ф�E��h[gǅ���0#���5~@q�d����r>�<]|[s���&�*��H*̩�OQAQ��%�ySbQ6�� �]��x��=I�Ɉ��q+����c������:��ȑ�#/�	��P"��-�����0�X��m��U/A�4��R��ҡ��b���ݜ��pq8g���nn�E����~��z�r�	��W��mF?�Ŀ�{����\�\�*��Z��`o��ݏ�&p�k���=Ѯ���cN�� p�2�p��.�&�a���U���ް�hn�ߵ	�'��#���!`O��gM.K	�0���zI�����J�x��/�*��Z�Ԫ��2LW�{����G���Ij+Q�\�ce����um� D"���\vV�D��@���}� S��u]���4���7hߺP��2 �R#~w@�6����w���hʴ����tbE�]��6�8�ު�b�O�ѹ�b=)k�"���Y�Dr6̢�(�#:���T�$,Kɢ�4�]Z=�o�Ly�������W�-�NF��%u���Ô>����xt�9]�Ҏޅ<�����ôy���!�}i�OQ:QɊ�o5���v%�퀥�9B�f7t�3��-*#���� d~.T�F��]��2f*Y�b��rCp������L�v��A�t%`�#s�ԜӺ7�js���k��5�"��t�K�>�|7f���	Mö7�T8l7M9���!'q��J���l ������ѣ�y@O�