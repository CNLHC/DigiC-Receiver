��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��$tgi����	�v��qNo�qt�I�<������r��F3�iG]䇿×?���~��m���� ss}6�� e�M Xe����[acC�=�r�sθc9�2�Cő���xeDr��`�{����4���t[ <��#��2����J���>7|i[�Ω�7Ű�Wr���aXL�\����$s�HςZ��&����g���m�.Y`R�JI\���I?���Sd�=�)I�&o���:�r<���������o9#k���&'��F��rƟ��3s��ʜ���05B���vv��HGDUkԱ�����&���VU��޳�OEk�����x`Z��A�5��n`mP<^z5i5`���:���� ��5lZ3�26'!~u|]n��uX(W�g��w�!#�8	�v�Q��(���+�T��m"��ʀ��3]���������+�!�j�ʨ5}��j���c�-�+��f�6I$Q�O�� ju4���K�욋�E@�
(cV�feˋ)w�L;0�bSz_?�J
��c���{�gB	j��\�w]��������#��[r+�:��(#���Y̯DFy�ǡr~��b��9�ѡ6a�fL� �+�3��Vޥ��Ec�e�R����|R��>=��A�e�|�MI�cM�q��O��$GS�6�})�8�M٧f��^��VʍNpa��\�@��&��a���E-�R@��s�����(r��+�D��;>�'�'@D��jh��֩2�巁h�/�p�C}��D��qn7|����֫?�����>�Ū���Fr ������#��5�O���c��ld�6�e�ו��$����T L��᥋�F+3���h.E�	����G�Sm�V�E=SS�VU�Fr�w\2N��������|H<�οs���!e��	˝����v�p�`w�'@��O�w��1���PP����guH�Ĵ���`��ku3͖�t̩r���{�;=�8K��"}^}gR��a1`'ږ'���+io�؟�cm��:��0��M�8�Q	�/�/'� �B�q�{�����ע��A�t��ü2s�9�\���߭&�>'�ʲ�q1�-�7+R��,���&�CۿR�; VP3L�u��A�bx�T�fq^��ny�#t��3Y�B}i�����K�O8���g�Z�S�E��D����A�k�}�V#���e���O(ͳ$N��q�+Ȭ��/�yzez*����|GK
�@�\���#�x\ Tl�6{f�*9�[d'v��b��v�k��E�_Ӣ�^��2��F�X�̕s�g�3��'��2�[v��'w�4�.����<���0���)�����4�n.�"@@�lk�E`�M����I�Jf�3

c��)L��-b2��[	���M��@�Y�����iX�@i������W��㣩������q�}^���xh\(�X\���5��-NH���>L�(\���3��;�":��1"'������]�g��xD���ºׅ��5D�S�u�/�pC��Ij�+�g�;TO,N^q^|����~-�-uV`����MH�I��s�K3���K�S�G�z.�}6h��+ꞛ+Ŝ7���43W���SV�0Q���tM謕�v���"�sSj�P���>�{�w)e,�ҳzF�
�N��/���ː�JnV�ŌP��	+<(�U��p�N�C|�zQ`���u���"�C���x|Z1i���_�ܗ*�Rݨ�%#�Uxi��Ǒ$*B^y��ܠ{�0��#9�m�S�v:�Kd�f��X�"�#Y#�ق�~q�-)B�����1/\��E���}�QTf�O�����fi�4ݘJ̰���q���Kz�<P��d:Y���/*��(o}%ϐ���������c���%��9E�W�C�����~�B���v91QܫR[��]=�O-拋�^��X�Al�Z�jCl���Q\<h$�Va
$&�)1���&��）;p>䅻��:���	���{�G~���Ngev�F>E4����ћ�/��
�<U��Na�٨�1���*m,ʟ�H36)�$m_���浅�̜�6�=��*�U����L�oKO����>��"V+�*F���������KpG�|�E��C��/�O�٩�����?��P���-eg���׳[��hY�@�(Ѳ�1�!s���K�||̠��n��=�2��8�+F�E�n��t2��X�Gϩ=�ߝr0 f�Mc�]q��������8���C���A�t�3�`H�k��ڲ�^��OAG��d��ӗV�~jˆ�Tf��ڿ��T�v�C�������b6�C�ɠ߅:���b�-$��ʷ�ֻ^��N��O��j�k��s�"�Lbь�A`}ȭ^�,��Ss˽��[�e�)�O��_j�Y�E�c�Q�h��
&�W���^x����0CS�J�N�X雦<�J.�s^}���.��5��q�����6���4���7���n3�e%V3�y�t01rQFÔ%�<
I4r4��<.�Y�q�P��D�ӟ��	�d`w�f�p�k@�o��"�Ϧ:�ØΘ�F�_�/�U������)Γ��B��G:���*�\��;�;��0��'�f�U�G���ϼ�0&�.���/�SÓ�6�Syp�7��έ�����f1�(~3���>S�ES��GqZ�E�t�h��R �*|r�(�c_��$���j
@��ڙ�M�WU�9���Ւi�u	�i�DX��S^3�����8��j�A?p����6)7���&7P	�.
�t��+���M[~�*%,A�;n^�!��b�x�V�5:!lHu�@��g�<|��G�s^M��I{�gǴ�#���(���O��А���f�	��Dxcm)�sk��61"�P�;��=8�e��t���w_��E�2���ib6���`�#�$ʐ�a�H�J��f����PZqS\-�R�������?�C����<ۓ��F���'�.0G�_O��K�?b�^	�������1x��������L��7�*i��1�Z6ML�؎A��0$r�0�E��)�����Z=�	T����Q�z��w��y���d����SF����nW��w,��7��0k즮糓t��1�Y��5�I��3���1�ھ[�<�DuAY�A���[�kG85�F�Ue��%����W~'�u
�>�k
��"	Dj�&�ZV���T�@l^�z!_�i	��,��<r��x\��ʝv�	b'�h��F}��^���O�c���Ԋd-�i�7�bE`h�9��⩱=�F���
�1\u�>�m�("A7_����9u�@w����7���d�Kо7���"�[*�q��6B�Ox�r��agg�[�2[Zh�qk�#<�8a�TW���5޷Ж� �]<�U��/���Зj�M�+�	��bԅuj%+��f��_ph��U%3�()�͑��/N<�:�(XgA����&���u�I�I]��|<{��a��^���ʠ��xv�^�f��0e�b����˃5	�KKPf�ҟ�"i ����LSHK9���W����z��Ʉ�u)�0`���i.db�p˨���������k�=P�.M�;���.���t8�ޣӣp�u��ycyw���b^�H,?H����=�9զ4��Kc�Xe׵�� �����G�-6����#GE]��
acd:�f�)�ƶ��jn�xp#HI<�e���vf@���;��~��W1HQ,��Tj�w@H����,��[;��$!�N<o�R)k;H
� �0�m���힠m�*gm'l:xt�/���(�,�g��(y��h*0�[Gv&-D�`�T��sر��~�e��w�
�D`c�� .Sw��5�HēA ަ��K��n	T(�q;���~v��3�h�L&t#2����<�z[�[�6���%z�4��.]q� ���r�f�3���6��vt
���~#^�*�~�_"����1�"~�#]��zh�_�a�i�	�&�<�_���,ύ4��庍޶Q��ͱ}����R�E؝�FS؍,[+}f ��٫
��+�W��i5�I�wH@�R��MeQm�m��c䄛Dl�Qɭ������3�Z1sl����J�c�*�R�6��+��tzs��A��ijE)<�^�H�P�y�.��Y�k����9��36��๡iwb�{�������n�O{k�fȒ�z#�Z�#���{��5�S��>�O����m�itu5T�qƬs��[D;���{���m-�3����tl����yE�A;Ý7k2��L�q:�7rJ��y�%�iH|ũI���<@Q�G݃�Kԓ�����*7�!�U�����Vt��.Ə�n��w��3��i���9����R]��|������V������K�!������K�u?����#��A1Yrw�\@��qf�b�SNOG|#�ѓ�R+%$�N���OJ���6�-\�P�n|���/- "Ek�X^a @kF�Z�M��g;S���fDq'߄��qPПA�o����Rr�MO�C�K+����\ �a���L?'��U��\�hu�}��7A�z��N���TD�m�{wPU�qf[y�q�@�KI����#�z��טm�����6.I��Y��O zzz��X��
�X]���>����ĳ����)o���;Z����i%p�am!9qPa8Q���&j;$���9, T�+D=���0��e��,0O*J	�A�Cw��� O�ß5��9�c��@ߠyq���-���oj�B_���,e*�&z�6�L�����v,��@Zrľ�G��^��,�ϛz^�g��U��0MfїP���࿺���lʔB`��th�*��{�wTW�&i/�?_�y�J�)/C���H��o�C�6eB>���Ҹt���Q(J��\����O���e>I�s%����� �Uq����q׮�)�1R��2���r��O j�@C���[�������Vc8�ɮ��?���:��ҥ����;~�c̈́fm&m(�6�70���2��L5��l[�,�c?s��MU[C�`�����:�R\x�,I�g�6��ߒ6W\���6ii��~�QX��5�a�{�H6" ���{�8�i�~}x�>'��n���E�g����U����-HA`�-��~�����U�{�Dp�`�Z���o�.�!q�"TYm�}n�Di��z��t$@�w9KCǟ���x{��"�T������gd�(�4�<	y�O��}3#L�:&6d`cZ!t�i�[��a���rB[��H��Ļ���/u�b�
㏼<E���ϥ����O ��!�%�e��YBҙ(�Kl2{E�K�2��(�/F&�����=�����,4�[�!�ˢbbfJ.�G�76|
�����2������*W�>+~@�|�;f�:$�7��c&�F���A�"����4�w�<kDޣ����GD�a�:�IPy���C�C~v��O&�\�H���@�ti�8iP���pJ�[����<ȂM�؀E�)yHo�wt�48S7d�d���|ԘK<��ެ+��� �/I*<[��ܯH�uC��<��P�,T7��ñٕ�<3m��LU�7�>E�|�~�Ab��l��Y�(a<�e�)8�~ݒ>�@��"����ƱW� ��hɉ秅}�1����~H�b�/��NP~2�r��`�F�x[��c���J�hTw#����RG�\`L�d�������_̠��z�a�6��"�z��&���<4��Իm)f�m������|²���1{�$�v����o�TS�`��������L�D��i+�Hz�J+�[�..�����~�c�Nd�L񸱟��c�m��JÛǈrMi�����Z!t�����g�����~D)`��n��:�o�i�>IUI�	�IueiV��~��{�Km �~���ٰ����� ?�f����%E Z�ߣV����l/�~}��'�	�dԯ�e7$ڮs.LMcr:�4�#z2�z|���c��p�;��R5���y�;���!�7T��>q̟[;�#�#S+��,x�B�͡!��I7U*i��)��XQb�����z�����{�Q����3~L�D;�nM�Y��2�.�e���P�?�R�d6tn}�D#�[z�ɪ��j/�����|�I1�n��*����6z�yن-r��RM�e�°��\Q�܆�yϊ��/�)���M�%��=o�RÆ��3ny�:�y���ƛ��ϝ�w0G�9%tl���Jιwy�9h���y�;(ӡX�U�'_i����_�ƒ�q��qcC��ږ	&���'�W}%�@�58�:%�+q?!Qu����s�h�§�a�Ӆ��0�ПV��<@���C$ff��$����o��������/�.���i[92|m_���ZE��ɘ�qǐ��v����3�xp���!�������7!�f�܅��̨[X�O�d6�z��T-塜��5�����6"�;D'���k�&5��'��ol('�P\!_S�˾JW��o��+8���VG�E}A�@��%)&{�B�~��(H�L��/�x��K����U-5�j�� @B	M�<p�� ���=��y�'�V�A����5r
��C����5m�]om��.JŔ�@N���2f��zC��Pq��w�L���fX��Rk��� �����N�EV��B����h,	��/Ҿ��������D6x�sq�
���.�_�*?���9�07b��"Ϭ#�bh��{���_�S����Z��𾮬�h�Yr9܆�)ｧ���ssy͇xݖ6����ك%��>�>��Ŏ$�N'(��!��]�e2�'S�
8�E������Ϫq���QUo��N���$����F�b�3\=�, ��<��Z6�u�؉��-��
���ŜR�y��&V�*���B�)��̏��������Oݘ�yxD)ӰI6w RG�^
�=��i�򟔫z�Q�Te=rX�7}��Ajir?�0����H4~�q���X�F�v�n^�>��۬�lm�������Y�����R��L��r2<9w۷�ʟ�k�7�A��IP֪�N���2�ė�}����v9x������0%�mw�doI���E����4����VH�z��`���IT�F�p��eQ��v1̣��Մ�����YN`%:�`Y��|�׊�a��;p��>u�ʓ��@(u���M)C�.�����T�C��i�:j�C���ǈaS١O�N������*WH@BZ��Z�P�Z�����rH�� ���ȗ���Z�F�=l᥋=���zͨM���OX���Q%�1���%��%�٦<v�j�;B��
�*�ó\E�S_ҩ���|s�y4d��Q�mrš�U���e�u�sͽ���ճ4q%��'���a?͛�zb;�~�:�ʴ�n ���	����>SL�T��0�5N~�ʭk���ݠR( ��̆Q����f� A��߿����+���r���LQ���A�׼kij5a�M�ʥu��_�z�vtkYF���h�ڧ�����j� ۃu^̘|M�IEFB��x��]�'���0����	��D�~r���bzh�`���)��a��5�&C �h�/�sM��+�a;��u�ؽӥ�#��=�1�¨O:G�����[����̸�n��}ڀǼ�k�_�	
�qf(�S�R�"�Ұ�6�_��~���Āh �8��s�����gR'5�4|cY����]��N¾��8�K��pWZ�禮��hXM����<��&��>s�����O�.@��$n�O� �M-w��U ��]��=��'<M�MS�(������;��ON�jh'�6�奪�����;�]76���p�S��!�ݢ�`Ӄ.3Q&ɜ ��q���e��1v�B�;�Lx�y&r���V+��+�6)��q���P�%�ƶ�G1�$�!DO�"�L�M��7t@c>����A��w��p&.k%���JZ�U�He���ld�F��� ��5��s����z��)Yvj���PdGm���1G�!�w�7O^��7�S�g��k֝������I$ntvM�.w���q�*'������@�q��d�o�� F����V���]���R�C�#�7A��-���Q
��t��� pT50�QK,a�I�&e��4s�\i����@_c�W�3�䙳'���UN/� �s70KR|�6G
���g���z�"�
&yD�NB
���Z�j��<�Pw9���m�4k��m��6W|�����AfEF���Ɉ4���*��S_��}{�"�N3.���]c�tئ����t7R}�ϡ�;�@f��i��)ɜ���u��Hj�,�WW�һr�ع�:8����UXA5��86���۝O�eAv����y'���:�!��ښ���"�'�zU���vl������0 ����촎�.v֔�0��Z��~�����_��Y��	�K��'�w�&���o��M�"�b���a�@,�.0����Iȵ� ~�F��c��Ł�B�Ǣ&�W��yR�}����ڄJ���{�g�<������i�Ն�I�c��|ےP� ۝9��_7?�Y�ërp)VL{V]^ke�d�ߵ���ଔ�ܬlO�M+�z��O��{��~��B���3����Z�>I���O`N��s����)_�=�-�@S��Ӌǋe�ጻ��r�=���+Z'���"m�3�"Ν�q@l@����;�KUӟl����ໜL�X�Y� i4�n��R��� f���~Ԡ����j�B��?��A��EY&���W��2R�Bk��i)��;c����-�E
����]����?DI�z	��ū���^�o�X��z�6�sn�"B�.�O����јH�N���H��aW�P��F�A_vd�b>N�I/���8?�7���f�~��J_�E�@�Io�4�L-�*_�����lc�ֿXA?�O@�F_��8�����C^�:�;���?�C̀Q�rUCG���,�=���;���rL�
��C��Qݡ�~��5r�˃<o"{�_��XN�/X�%�������s�8S�LN#�*V�T�|yc��nzO|>1�B�)�H͸H5 7R���&g�zf���L������(<|s�K���m�թ������ܦ������ٓr��]��h�fi�v�{�ώѶ�� Y�ŘD�3��l7�$��T��i��'&���Ds�a��Oy�MGZ�����⪸���R��n��� h]�>�S�^��ү��C
A���! :�H��U����'-�G�a�?��>����7���7?^y�M5���Fn}�N
g^���� 9 �
��O4�*��̭O�cC3ѿ�0'�k�$A��(�<�2M��qvr���e:t�0����2�9�N�˔1�9�/m����.#nQ�c�w�����ޣ��s��
��Y�L���ۂ�ɜ��p�y�AIS�cI�I�FV�i�GPf�@�7�N�q"�$TR�Y�>�7�m�6| Bs���q��X`����O��vɑ)�,��<-����K8���x'� ��9�Ȕ{].xtS$�b�I�]��D�x��{��hEc�F^T8Jb��B늗�b��j�fW��;P�࠱(�K1)�d��N@)���UdѪ�;���(����>ߚd�A���5��xii�<Kp:{�^��w`-`�ؘ鲆�|�k(�$��nI-��U��Ku����A�6�ko'�W���>�`�\������	_������I�
�p������^�\�J/��-�v|tK8O�,��Ľ,�8����&���9$��k�t���)����t�rE�����[�]�p��X�N�n�^��uX�O��ꪉ�LV��ǧ��G��d�_�i6��"�9��q��OF��W>��re�A����\�ͥj���I2�
olL�<����������'����ҜԲ�5^e�����bj�'�)�؜��g��7ƌ���6��~�4]B冑l�[� R&
�.uqb���Ox���"���s��ݞ ��Z�5�ީ��p+�����4 �Q�{���V�K2c�Cu�=�&F����r�7�&�i�Hͣ�Xy4:Z��e���I������(�;
���H+�X�-t�2��ʢɏ��y�j�2o��@��%'��oRf\r#��1��i%�B`f�Ri��}�c�j`"���I�%���ӭ��)sQf�&j`	d7;� ��͌$�\�#��^0� ���xk���{9?f53�Ƥ���� �Wfp�{DcT�D�0_���0���ϥq.2�ZE����V����N+�<Ǉ�|�V�eɓ��U���1�>0���ƃ�|��z`��C����XN��J>��V�i��,_�q��%G�o�э�u����/>��Sm &������A�F�- �
I���*�3c)�$|N�~:I�b}�s�(@�`�kc~�"��u�j��X�"K��K�C���!Х�t�bf���y��N���5-����|�|0~C�T�!|�Ó7
m�̤R��P{	�$��n"&�`�#���gR�&a��/�iOJ[�l�$���* �
�c*j�/�)��t�����Q�G�Q��|�0J�}�N�as��N���ɡ[(C��CQ�u���(b8pTxg�T���yz��RO�B�(�sPL��M��r�~�A�UhDB�`�}�KXP��G��(�� �4�R�Y��\t1�	J_G�Y͚��$�oь�dc=�F��iDWRj8vc������h>���nF�T�w:�)�S P�h��]�l��2�>/sZݤ�Y�.a*#���*�3�?3�#?!�������A�2���_tW/%!�
U�X[��N~,!����2�E���T�3�/$�d��/�O��/�$JF��]�E�oq~�����Ȧ�&+ŎC���T#����)��ZB}K��,�ho��N����Q���o+WA!�9�89���2ߩ���\6�����@��O��]jR.��Ы0��^�t�GjYt��.y�p8�����G/��;|mN�$ R���	�&�|fzs��2?W����^�"q5U��z�Ҵ�M��A��.6�\�ڮ�c� �W"�^�`xV�f�w=���0.[0����/�4������F�j�շ'⢈߹a��dnɸ�&�Cl@	wًB�y`��<�a9�$�?�4�&� ���/��~R�̌����좑�4P6C������L���r5���8:��W�ig�j1�4��y�)�J/�V���OS�z�H��﯅��r��f�7����ӵ�՜G�������2�$��\�t��K�1Z�:7#	R�pEdO�̤���hTv�K->��iZ����1�_o�x0l��gF9>m����^�n��l��}��KI���y󌼗!��l�9a�&̫S����E_Зqܠ��ǄD}�?��ap��!�� �?�x�����*�������� zsa� 	��O>��H>y�Ŝ����I�����N�c���M��=��h+�#�l�	^�"��E"�<x�S>�0�? �V��� ���T{f+x�y�NA��w<i5J#|4?�>@+�,�5 XTaat>�ﲮ�4�׈[o6奺���Sʗ�-I���pB,*AcI�lu���P[Z�d�$�~�d�PO#�Y;�6;hs'L��WnS�����'ҥ��
)�7cU����(/(S*n�N����[��G=�v��oo"��e-��d4o�̦鋖\N�7���O�4��u�4;��=����Nh�,�0yZ�%���Bخ��}�]M�ʷu�&.�.��[��綣�A���ҿ�Gc��#)zib��d<��F��X���l1V Bj8M["�x�Hun��je�K�Yy��4����w�Z>Y�Ύ�"���[��ͥ�D~�}��x ���ʕ�q�����?W�����(B�Ċ 7�{�?�9��w��ʇ��"m�����sF:_�vy�;Q�V�+��l�ͮ{;�S9x�{��V�&�Md�[����^���gP?�a����	�C���ݾ\+��Y�D~]��a������n��䜋���A�Pkz������hN�V��#H��{��J�vo�X��F�:��x�/�A˱}�^�pw�ٿ��h~�[�@��/r�T�..������*5�������Y�(kG{�Sۥ����R�^�eֆW`B�6$�A6,}-B<^��"���,|����'w�V��hK�T��b��յٷ�ҡ�9�'B��&�&��h�[�:
�1����	"��Q,:Z� C��h��h������T9�&����y��Q���Z�qR�(���zy��\��o�#S����q�RiS�{� {"d]qt�Y*l�T� �ʜל����ʞ�����I3,ѵw�[�t�\ƅR�%!b=�x͇�r���oЎw�^���ŏhf��ap�J�Nq��n1�B��J_	N����t��6:�Q�9�l�M=��?Zé�d������"�P|m{��Ndo�<� �!~c��I�J�������W^��kh�Dܰݪt��6Q���n��[ΜL�GH('�/'ٞŬ� #L,N*y8�#�Cc<"��sZ熡ć���!uԥĄal��Rf�����琒�/W���J�7�[c�$}���*N:��^wԠ��\�� �W���z,���|W��� ����I�P(_w&�G@���ۮ�&