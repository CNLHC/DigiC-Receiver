��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk������A�砡{����'�{6�WN��U#�]Miy͍�2��*���N�R���1�*�)rv���̎kf���Mb)8��ǵ[�I��hF ���8�s��d�9�ҟ��a��*K���qN�z��+�bğ��2��|=W�*!Im	e#����FN�*,}��Bݏk+�	�h`�u���p7n��법�5�G���+�Tzܾ�q��5Դ��3���Ę	��<�ѲTA�%���78��M��yd�Vgk����u��F2�/S���9J���������qF�J���]q����9C$E��ֶ�2cz�Q�tZ�ȋ��x���'����k�T3ķ'B���,Oh#,��`�E�F/I���P��I���;�i@��j�w�>d�v%뀂�oZ�i�_���e���E��0�V`K�k���U�L������ɥ�S��WfIt۾�Q��=_�u6��L�������W�bW�6me&�x���8����D郝o���t ��d�8���A���6��%�v̋�� %�4^6���}��x#6� 5xZ@��h~�7s��2^�`���f"������t�����	e��n�E5޿��4v����b�Gb�ӟ���POhO�rƿ�?��S.$�_��J��(@P	���t�I�BU�M� �H}��5�[	�@P��;�	��e3r��=�򝣎Գ�Z�G������c�G�__H��'�A��PVw�`lP�K���@BC]�?�;�5[z�}�������:d7)��I� ��>�f�����󒠗D�-��x1���C�,�����^. �����b�?.QTf =����\�Y/Ӯ!��N��/X�(��������ـQ�\3���	��ƲJ ��p�w9�����~�D���¬��zS�4pRj3�>aH�ףҥ�Z�U�,���R�����״���X��pvـ��F�����1��G����~x����g�ӹQ^2~�WKc�,��5���������Q��f?L괧����)���(��`s���x��b%jΌ��K�l_N�L����V�z|m@6JQ!z����xi���x�{���'�����b�f��4v5�	o#M ?���3��.�ʘWl%�պ��1�r�����5,RK9��Ly��B�=�~��3.�GKV����}|u �r���f��s��2i�������d�);���"��C~T�������l�qj�
�H�0a�Vs�i�olG��������I��ثh�G�����;�8J6�Zsݧ[+�Ɵ5����Y��O��E���a�g��V��,��~��E��1�}�
���y�DG�ixo@�Y�|� ٷ�O2Ҥ�����'s����6��p`�0�o�3�uNG��ې�'�J���sS{bq����$�P�B��)�t���(���[�N�5���5�Z��0�^�F_� �����P�������hV%5xsmB��^X�{�#'��P,OD˰=ح�a�Z����{!��#�yp0�L!��e�Ǧ_��L&�[�l|�Z���@������;�&?j�#���1ļX�\��}�).G����́��S]���	�%}�\t�sۙH����X>z��l�n���	c�5/Ǫ��	��2�b�9`wу/�O0j���$�!E������Q�-��'��u���b��_�6ٖ9����q噆�����+�1"q>���귃�ᵒ׃m��أ��3�f���Q��,W�Ӽm[�y~�z�*B}��^�p�X݉H>����%��
X��svukʛ>\/Y�?��a��y4M��
@o4������grtU�Mbr�;e�� '�cRL�"Y����O$I��ɵZ�0�e7:��o�"��\�"��%��]/�j2�I����3�ĀWۓ��AG�]ƙ�o�/��Ya,�`@U:��׽U�.*�Y�rH��M���̀b�52�~Y��nĜ����I��n�7��u��9Qa�3�eg���� ���>��6؋����uMX V��PV�N�,|�;Z�߹ݝSx5]WKbi[���s@_{���UH�d|�G���ռ��6�o^�g��_����CS-�E�j���=~��=��ֵ�Fp�C�&��������ѣ`Xx�^�mrw'c�;A����:�kS�
\�<�,E'pOݦ��.��Z/#A�wDr-7L����M��A������a�7�r��8܆�7Ny�Ŋ���
b�ߙ.(7_a����0�����qKyԴ �VP>�6 +��@���Kf-\���� �x[-�`�q���}T>��΃yNg�JV�s]�E���0���Z:H������i[��!��7�'˴�^����*�,;F;8�~P���/�}p�1��ӄؗP�r�9�l�k&O�-r��pD�-ǰ�����t��7,7W��|e�q�9e��ͯ�Yo��7x�3Z�Dp./j���3�45�ר��L
�遈��xRx��������W��<����?�WZ�%%ykyj�h�׽wi^F�mMH�+����=)��e�AF���_tAx�o���(�]�����g�+k�h�ٮ�A��ӿ(bz:|%�Jn�Q��/�\���n�[ *w������{��W�����T4$���?�:�=�r��٬�uEE����Wfc�)n�/T�?@�$<��AY"MY�f�R����u��)�I&�w �{�ej�rD�&$�Ne������>�&�7�9�M�\�T��&�n��F���f9�X+�.��bυ�T�
9ù���M4·,�<��$D�mi%{zR����yUS�:�S����b髵y���G��+c8>��Qݮ
�Ê�:S�JZ�,��2�;�C#�6X"O��$-���hP�(k�.��(��q;m�:�;�V��ʓ�)Y흥nw�)�!�c7W%n���u�W����D�U����{,S�s����̅G��8�e;:��3���C�L;�����s�}R|"&�|��G��bf9Ѯ�ɤ�~��qLyf�nW�\]M��ڄw��s>Ó�n�b	;�H&:��{��Ȉ��/����M� ,	v��N��+�߳���f�$�������A_[�LH�4�J�����c��N���Ybn�@o���=+g�����)�IV-��ǫ�m�㤴�l�w6� <L�B�/S֥�P���:�e#�"5�����͡^���+�8 #�5̩��e��݈��M�����]Uo)%)CV��e�%��hylۚ��ǭ9��]<�B�R\�x@�v��C��J6�X�Zi��_�����O��,�0@�Y�k\�j�x��"*Ę�����!@_գMvT�A�����+�l��$�b�}`�9��r凵$�_,��P�� �)dD�a˝G�X�T�^��c��(`=� ���=��53Di1��'^䝎,�U]W�(ٝ���pDm\Ւ/+��&5	�ڒ��E�&"y�����ر@C��a@3�������Q�?$IC|��Z�� ���JI���m�� '�7cJ���&�)��G{1��[-ݯG�Ү�a�#��,C��|�'�m?/;FQ��`*�̼�A�'{�� <��Gw�GU(_��2��{���ǳ�Z��2���\�L�2�*΃�����,S�G���'���V�.��A��Q���D��0��weS*T�}�����8F��2�Y�ȃ���?�&k�Xo�B�6�3�J_M�e8O�x�z(��VgW{���U"?6n_G��B�����r�ߔ��Y.)�{��Z�������}C�:�w]���S�zkM�;����'5��x��x�$�^���1�m	��|��c��E�Ha�#���@-���^dOhVF�e�y'*p_膦�m�&c�K�n�4ؼWt�Gm3����72�����F(�O�a��`G�F� ��S��r��3�x@���
�Y$@�	��.�z�Hѥ�V]�Sl�oH�bT������������:�����e�3[����u�仈#�8�l��Q��I;�G�7�`��][���.��ni5�{�����̌r3��ϱ�DE�:l�|Ū�S�B̙%N�KTF�|�O��;�(Vܔ�E�X���㵑+i��w7��͙>xq��)���I́{��΅�0�E����`:r�u����v��x
}u����<�9߸iM�ۼ˂�J<.SL����)�W2�B�y� �*�`C?�M�uN!�e�ob�5<�����*�P�-	�f%vf�F
b��(�h1<Ϣr�Y �R��t���h��?�E����I�`>,�nn=�jmD)���p�ZE����KO2}su��Ez��ҕ�;H��=�7џ�L�76j=���{+�\��X�1�U�W�T��O�nx90&�Rѭ��?$���E+��)�E�qv��d�C��(�@��z�����H�e�,��	@X�	X�h[A����2�=#��p[2��×�_��̽T��Q	�K���=R	�! �h��6e��bKn�g9�w`��0Xum�ߑ���<3�Bai[�&gGBҿ
T��A�v���L��D���0q� ��?�X=M�
���E�5��uO�������;�%8��j-^�i�D!l����AΝ�R��l���G��%��e�`�N.�|z�a�J$+T�c ��W��|Mji?��@d�P�M,{�������'l�`��Fw��c,�}�\��3��)�kD6�_��A�z�pC+�~�fC�j��&��~�a9���B��ƒ`W)�GA�ʵ��P��F�����SM:j^�;J1�+  �тc��Pm��=)�,���8|yJ�胊;��_�����.�qX�J+�q��X�%�o�DF&�v�Ͱ�(Ɂ��l�\%xԀ�oL߷�銋����e�%����2���{c� � �J��8�U�vHj �����|�q֢a��*K?�h��Zl]�%KM
�>�b�z��]u�1[�̫=��M�Q5��M@�"r�L)ꏷ���U���Ή.B�r(�'����4�|(��zJk� X�V�b�&iQ��.��s3�������,��*��v(F�>�$t�i
?C<Ǆ�{RĪ���xQD���)O��oO�xӰF����Q��'k:�@sT�����:�J���_�-B4�G������\�za��Et#<15�b褟����s���<��ƮH��͊�\�b�zq�H7x��a^X��8����#H��(�y�������л��ɞS!/s�ӎ�:��\FS�j�rv,)���{�磦�-x� W�y�<1?9J,�z#�~�~r�'���A�=��W��������E>:���珴-�Ld���0�Xi��0�����b��C_jd/�&�z΋lM�5��T�n�es�_0/�z��V���n*�;�4�<�σ�I����}�.�������!�݋D��%,0��B�87���k]�lu^0�o%��V�v��G0���o�~�s8��G��z��l���"Hσ���J���f��g5�-x�Y�X�ML�(\G�<iO,���}�#ϋ����ZI ��\��{�"-i�`C$����tc�8�0��A�Du�;�:h��*_mΥ�V�����[�(���
I�l����<�ՉX��ψ��S�E�zwc��6���si���F�}�qߢ�ʅKpm4�gw@��6�T����bN�/�A��a��(�$jqs��<"�z�1,�*���m���/};���� ��b�ݳ��o�H�RXv�ڣ�1�	�&Pi��f���(�C.D/�$��p�9##�����.��ʆR����S+7�A�4��j��e$G�H����mmc�3���DSY���ݤS��?ęȝ$�}ҷ�cn�v�2I]����TQCn�id:�f���MSw�eΠ�RߚC�s)�g��=��q��i_��?W�!�^�����2�
S{���S)v�!�w�h��%�/v���+���f����E�/�R�
��/*�$��w]z G��НvӉ�e|��W�&�Y�m���=�$6�l�c� �@�~����t��U�K����u��)�|ۀ�N���G>��$Z�����m�.�Y�[��z�I �R�L��]���z���N��g��Ჭ��0כ;)��s�;��r}.�Jk�;�Gc��񱎠J��ŉ���Ǥ�F��'0��-�9�,BRZ���*��e}B}`L��6��e�K>�_վR��Yh�2��)�2����T�t�j�S�P� ����g��Ǣٮ�8����"A�]P Ic����h�^�P�A����B
�	m��$2��{��U��%{r�:b���R���Y*���o�5]XL�|�j��+�/�ۖ��a��R�<
6���ԑ�w J������lG�5-G�`hЎ��+d��n�6��휬�N~��q�F-�{���d�MkwZ��rA��FzOF11��(�I�a=Ц��ab����8���q$���v�zܣ��p�h|��y�f���O��f��I�ѵ�2�By1�u��C۶2DEM�B5g��z�,��g�G/��Q�~Ƞ���e;�R��I�^y�Y���^��|�OuN�-$pL
ճ �s���|�;K�Ʈ���+r;�v��L���L��q�0C�Ha�ۂ�B���p>;��JƁ;����f����_/2�w�zF�BoZ>T�Ia��m���9����@5�N�d���\�pU=&���,[��j4�d����=��������m���cȗ�zܢ�c�_"ɷ�F�b���P�	P����[��J��{.8C�j������iI(JTD�J��7��z 
l"2������%��K��v=4�(��}0��Y�Ǌ�g��j��w���|�[A�L����6;��T��N��-��9W&J3�ft�����?�%]�'B�6���!��eF�@V5p@��_�4�Ӆ��P@6!ʇ�׳�g[Z]��pkk��?3l���:���#���V��c-��.���N��Y���\��`3�*�s���r���3����T+�ɸ�4���.���hC�6�6��ϯb�S���>iDA^�\W�����-���;&P���?}� ��o�iZl��9���H/nJ�Y�	����~h�P�D3������yUC����h��j�IL�f�V1D���2H��'�|�Ix�%T�.��u��+u�+�!�T[ڼ8׸%i8t�:D�Vf�݂-שּׂԫ_b�2��©�mٗD\Pz�x$a0[���b9;q�D�2�v��}��2��ܧ��o���(�MW:�#x}�G/b 	�i8d�� i��A�X%���m�m�"�0��qJ君R�q`��h��ѳ��R�M���t�gD��Z��4M=��AR�j�I,����K����-������X�~,�%~��%c�y��i��60��8B~���75���΁
b>�*,.-�3ǁ�?�a����pa�=5oe�J�s����T�q�|o������؂�kT#h)�SP,�ٶ� Ҫ�e鬹�(��S��4��Ǡ����J�y��J��Q5אH���� Rb:�~@��P|�*�nق��7z�����%�>YU�40�~}?i��1OD&XF�[��m }�Y�8�.�ۑ����/�5QG|�k�˸�-߾�7�~3`�>��9��d�u* �t�J~�"�-m��A��G�Ȑ�e�<�<O�R�栯!��|�X��D�K��rZ!G���Al��/+(KX!�����I�{Qh��b�a����y1vO�A���<`��N��!�ZsT���nNOYn�2U��ha+W��Q��1l1�
��㟉=�9��+���j�dH��+7� !@�m��X+�O�=p\h�pI�;�OM	��f��_��4�bt_jf��4�����PmÍZu��#	FF�h�˪"Y!d���]Uw����48\Iփ%�X�6y]i�z���Y��hj�vH�2�DR*��%��M`]�Ӆ��	6oy.��«*�ǿk�Y-ȵ�3^+�L�� ���w��C����TK�{����D�\�\`�*�ް	���B�A8E�z���7a�������䁲H�6Ky�uT��\��D��8,R�L�:��l1���f9��G�^��6�������8罅o�f��aC�� �}�G1�U#i���Ix�'M!,���9��Z�y׭/؝wW<Z,�V�Kw����G22l,H?���đ�Aʏ|�j=A�������:�i��/����#b~��
��F~�tuQZ.�)��Q�nӅ|�_�p��y�t5��&��WWO�)Y��M'�Mk�k�u�ORU'��G��b*����Հh�y�G��ٳ����t��Xݮ�XAY�Kn���k�t�4a�E��*��i�V���("i`�����&�m;mY3l�&µ �6.׃�$2���^%��[�(��LT~��]���]擩�u�׻Z�;Μ�R
�8�׊#F?����EF���rHYJWJA��Day]S��Y������ӂ�HK��ˡ�h��\��F-�=��T�߭��"�@���{g?�+'�}a�Z"���.3j���8��j�9\�ȑ���*Xv�n��ξ>�j44����!]��a��9X��n�ǎ0뎇6{U���g��GG�w���;
�^X�Ws�<lfF�Z]/��^�ㅵ�/��I+��W�p;м��˽��ð�Ч:��yԌg�`6�%H|D*1�u���x���YS^NL��u ����$ev���ԍ��r�*}}���.�����V�z�e�v�bh�G&	������۵�M��
d���t�k�ao��Z��j�A�	�����Э���(���y'�M���
�G�z���;׳���1�ޖl6��˰��8e^��,kY�R����bH�'�ܾYU!1,��9�t����\ ������3��Z �?��$V��Mz�Z���C�M�:�LjZ�Ѽ;	W�4tߐuh��ɺxYF� SK�@㰼M��0��#8+"���rWQ�l�]��"�J�C���)	�?:��`�PJ�:{#;io�O������Yy{`5�ْ�6�R8:�CGN��KōA; J�K�\����+Zo��LS�����3�`�׶�aȐ�{Z���a�ߛv�t�2E�����8�碰c��L(e]�3V;`-mϰ[�7D��[עl�7wv2:U���Ǻ��x�}x�4	O�N[L������|%-28��,2^[h�7.���V*����;����^W�����[>�"�1��S�X����zP�ɀS�j�(��CIj���N=oY�@AZ��T�Ê3H,2��}���$���[1���|!�o��E�[ٔr\������2�h4����yUořӌ���6v�tA�8�t�Ɔ�g��X>�˒Ӽ���[N˃�)JV3O��:�f���TA2cM�ꎀ|L��	R��)5�F=�݃quR�PP�[8~�9�'E+�#�����S5�� ��I��f��@2���vLq��[T���zvH~Z߿[ʥ��mGt�ϺG%Ý-eP�3�$�WD�*3��>+��I�����0=H!���C:���&�"9�yUGq���)	Y�{�A���Ҫ�ޚ�C%�R��X_$vT�c�0���yJפ��K����"(50�fn+��=y��K'��O8���0X�H�|^���?�R���M�%[`;�)cz�����E���B{�옿��3�<{.��K��9��'4~k��ٿ�e,��Ub	mxXNt�ի�Ȫivw>O-�������E�<���V��i��p�K���R��Ď�'xj����Z��X���\�x�b��x5l�!y^礥���y����~F�>��}�������V2D��!V�u�?�[s�S:���d̉\�Z��膛�p3���C�.m�;�~�y�R{�`rOq)~[ؕ��x��ݝ ��#ޥ��I{��hP:˯{Ȕ�;sn(X1�h�y��p�#&�rdm���?L�+L� �/��?�$�V��-:��},�6M]��)��tˬ�A��gD���K��9Ɩj��bM�J����6��槼�K�ޱ�:���~\�i`�L\�0��D��mg-r��l��pk����2^"h�{!Ee�Nk7����ڠ��g#k�6T�ޖ���&!�z[���?�c�(�h�rg�')�ťbd\�j�V�Έa��@�RR��V�����p��x��m�y�[�������b��.Dm�8<�q[x�/�?�����65�s�g��X�O	���D�����ig��E��������z=c���īb4T�c�-��0Y�#�o�L�(RП�'���3��S�����ór����E�r��\��Gb��d�K�/���!�ș��Y�Y�p]	�;�K��{����o�m��O �H�L;��M����:���)_���eg�ҐZjǊC�&3X����:���߈�X��h���zg�<Q8~��D�^�i�-W@���ч�o���Ci��lh**n�&5>��g��Ux)?U~A��9�+B��eϑ��M�Ҡ��{��~|�v�im	b��Rq-*{������i(���d���.h�������\������/:Ҷ���:�g57�:A�ە���	�A�	%��\є�]I���1�;i,^�7D�	{�F�����IZ�0��/A�����>���@ߣ�iq�)����Ó�d��)��N�"��K%���[1?g�[�z�	��j�S�c�?� 2IR�+��Ro�U3��E��T�4�".��������"q.��� ����'�m*w9�c^�%b�C�JW)����:�,��E���=��Fڧ��:���;����uӱ��PT�r�#)���/�:�z���j��Q��oH�8��3#W'���$�Ԅyb�����(c2������x��7��(� N�旵Δ�v"�?�t`;�t)u�����l��1����&�A@�JB�#��J��k�vY68`��d:�F(��u�~:o�˲Q�x
ɣ����M�)pQ�3.J._�i�\+�|���&���|�^}�|"�=~�`���ǻW>��=ybi�5g1=��5���b��D�J��0�-��Zέ��A_x��jinCo܃O������dQu<�Շf�-K�h�<���P�FT��/�^q�5;�ڴlH�P�����ņ �$~LiK~R����,�Mn��P7>�ű��r���n�H~���1�����p�ĝ�"��+����d�?=0rZ^�\�w0;�̬��<�|S2~�8�(��H��oԴ}k�s�?�1�WB�	!��Ewg�ּ�� '�F�,����Y1�Ѩ�d��9k����͢�u��ӯ2�I�5������^�^A��-<Д�n�a�u>א��8��X-⺖�/���&��:�N|2`Z�gn0�O����_��J]7����O����Wݺ�+T�tI�k�U�0BP�ađ`"P+�{f�H�^қ�5����WR��k�lݭ�xoC �ȴ0�z=J�Ue�>�)P�Q!�,$��/��E��Q2��P�_�6BO�@t�#T�x}�R�p�"����j��r
�Dn������qQq'�2��+(��Ŷ�V��S�"��O��6؂~���"uD|�:�`�V��
��� c�uk�4V>�q:�L�o���2�~�����=:��.����^ð;���܍'�.�`��Y�����TU��5Vl�-4��"��Ǫ�R�)�5ֆ60��(\�yK�ʺ.I':��gr����)�RV2B�|�XھQ��:�Ksr<}{��kJ�}Pދ,� �F���ux�����Ck"�[mY��Ӿ=��
��q	dKe�DVVP5����9���V���6��*����{��!���	b�j��n�����F��j��jϘ��VZR�=C�O���a��	��R�rZ��"���ބ�����]q���I�G^q:vF���ؑ1z�J�f����B0�L� ���"�.b�R��j�cY�`�A�㭼P���4��h=<0�{Ԅ�Oe�8mB������]��h����vw2��^�o��Y�c��ȪxL�����)�3����(�R3*��֣��-IRѢuaц�Q.�q9���I��V�4᧳0�?�#�I�^k�6!��I�3(������L���Ho��h�et�C�7�Q67��dQ�ѣSxϵ��C���n�X�}}a�t�^�4�	ч���H�Mi"�������N@�q�-b��<ڂz媗i��د����>���>���g���3�7���u���y_���J�`��\�.0�L�H��K>��H�'�mD��6��rG]<DUB��󾵪��4O�j�[\�J������M
5�*���f��6�(����My��t��"��CN2챝 �X9B�%���T���lz(g@9��۲�tٺH��¯s�Sȿ������%�̳D��eiM�d^=��|v�U�1F;3Zx_3]k����݂-�E�:h�&�[�����zb�V�iD_�<�a�(|N��M��+��K�;p2���m�S�vε��(�����8vr�y�����i~qc����0�q&��4DG��b��t)'���j�L���n����T׆`ūXrĝ����"	��.� �a�FGo�ݭ��qte5���6r�O���U�6+��2�)k�.}�݇o��&�l#ta�@ Q)QnfV�.���6�A@%�9�p>�����R�wj�@6�:�T�.�ԑ��*=�@g�k�R�$��������W����B��r�ʷ ��z�M�S�6\���n����3�Ey�܉:v�ز@fF�z����X%�y/��TA&��yV�s8Bj�%�;�&gB��:���C�s�ͅ�P�
���xG /`Ԙo}!#+�q%��.�Q���ye���y�[�~q�W�����z�/�)�Ё%r\��d_��C��"x#5񵟈qw��5>����x{夯L<�W^�BnQ��-�c��7���W�c9�IG�ؤh��d��W��r�����T��%EI���4�1V�p�������H�W���a�+D�t^���>�����=~����3���M�~<J��5�����U�VK�%a.?�P��g�ş�UvLu�̔�Ҝ�*�QQ��$\济��Et`5���5?w�%�˴��c{@�x�j#GY7����,TV��!��� �ƈ.�ӓ\W�&�0�茏W�fYꉴDMIϾ z�8�;���XȆ��C��^d��j������Ǩ�v4H���X���|���S�$�U$�1Y&x%4?�s�_�R	���ַ�gqIڽ�ON$e�B~<�i*(;���lL�%#��"F�CBW,,Sls������;��w�5�r�$GÀ��E���,0���y��[�"oI7�t���DA�Y��9I8F�1�*��#�?4D�h�W�-�y^��W���$��L����N�R�L�x,t�q8�GL�̟�z�3�0�����Fl ��E!YQ<��˦=�U�J�W�x��oj �f�c���R��k�.�+�&	s��WȲ^��_�{﫩aZ6Z�Noqyq�YIǂͦ�vJӈ܌P�DR>�7C�yl�R��Ĭ`���S��ؽ�l��^�3�e�K���N�G����G V%�r�L�KH��	 ,w?�������V'�j�HK��C
m�D��u���-8�w����!UL��E�#�c��$�LX�5nm{D�;������\�>ӈ�*_,k{�e��nl5�K��s�1�%� b����O���j���Q�vzǙ>��Qޖ�&�>����u����~�n?j��ءɾ2'���'y�_@I籴;�zT�uXo�b�CG�mk �<�j�ȉ|��m3���$�`zƅ��������ϨC��ɔ�w�U?�4ď�`B�B��(lփB��|e>�l��Q�oìc�䝑Q!��.��F�ؙt����*+����&Z�>�ePб1�"�`���tݭĿD��\�V�e�w��ml7�����������)4�}Д���ۇ�J%�(��?\$+���ğ�c�a}��\�/�.�C��}}���Ѷ�u��o�g/TP���p�7;{����Tr����Y�9�FR@u���\�{&�4���wU�ʈN��(��d���ɇ8��+=�������J��|+�!�pk����F(�����;�6N�
+���ɨ��o�"tXNE�p��:$�n�S��{'��ﾔ�=���?��+VaCcUW��^���I'�C�A7J���m_� ~��vd����Φe��<+!�!��l���Cկl��DÊE��T1mjn��t�`��O�ܳ���a��:�th���}�|�/�'�b ���QwMӨ�	&�p`t�{�f�wo1�M7㧘}������N
��H�D7u�RBi�ڎ*�x?3P�_aA��Rz���S�|��5����P�&����G�I��{�)�P��J��t^鸪���/��i(��k��Tz�S+�h��q��"{Lu�[H�y�i#C�<�b�P �±��Jx���J&U�	:�?����������Q�����U;��o��~lCH$^�#�'s�<���b��Ԛb1�_Q�ۊ�����XD�C
��f��T�=��D�w�����5��r!�?���h�G�I)L�����K������؉ѵ�d5�GS��T˙��5X�[�g��+�e������m����,Ab���1���k�c�X[�ɦ��K��Ie6:��;�ty�����+a� �DC}><̇PFS�0���ʵ#�SQ��e��5�5k��i;$/O��ŷQ⻍�\fN氕��� s+�3b�>%;��F��:qė�3i���A���iM�Ki������:�<�޹/�}�y������ "�X�1�ȢXg@ch�����I�6���n<��":����.���,������\�zu��ǷTs��u�|�erQ��1;�E`硛HC���j�r ���C%��s��4�
���^l]���{��΍���'D(A���^��_��%�BL�e�3]�^���ޠ�Αqak�����;�T��^��qG�eA&������%�gk3g�����)��W-�2!��!�j�����nWdk�5-���E�` ��q��	��2'��5#1�F
�;^��-� ���p�f�ⲩJ3���W���؟jK/�5$z�apr�#
q�9��!�zu̬��l�;�Җ�A�&<n���gS�Ex��<fQ2X/�il��q�?��MnZ����B�^_ j���5Y��V�Y-@����}�&=�������2�]Y!AN�]P`��bhQ-�8����Hq�+k�Ǡф��v�<͘�\ ��Z(qs\�~�#�.ݗ,;�i,��'���WB�l4&�=(�q�����Ҵ���;��*���6z[���H���˞�2����d6iS���g�4��v`�������a�n
�5
�R�W�JxYɐ%-+��Ơi��@���[#~1��?BF��B
ջ[��*T�o�nd�g��-Mo�#.�7aް�"��W�b"�U�S`���ȨG���B~t���TT������eA|�F�-h�CI��s��Ϙ�lN�]�B	��S�����:���U��j�~�Z���˵Y0�C�N�}����ה�m�ȉc-�FRı��!�y��I�
��tH�k�r7�'��Ldn�ouIX��M.�/��Gl�ۂ�c>J��ܘ�c�dJ�~?���ovk��6���T�zq��T��<��pҢV}G��� p��>�M#�XX���Tȥ��Q�-����Q�'�ŝ����	���9�lm2Re��4C,x�Zה���M9��=��l�)�SƂ\Uw�g1(>��A�*��S,Fcd?<� @4�#$�Nx�!���{�4�ll�}�l�$]�F�6�Ԑ5ᩴ<L�E� �a�G	7	�P�#�W^C��Y?�d�:i���j}uV���5װ6Y7�d/�Z�p�6�>��p��!��!qI�f҃�y��^�+���t2d;z/��'���4�n�܎ �����&�����R�)�ޭ9�;52Y�@A �/g�@��џv���:b��Q��n9��Z�=H8��:�D�48h���I��zZ{S�d6r�͢~
�(�16����1-O��Q����*�Ą�gD�� ���b���gRI��3�1���#��t�Pd�7��Z�+cu
>����N���o��'6{��}/���$��t�M��YKZ��1�E:�wڱ���J��q*ul�-��.߲�DD��0Z����J`�*������&�pC��(�v��m�$/Z~z����(K�%�	@6�{`69����]!�?�C7=���g��<lEN~�ӟq{���f��SP%�7�����Em�{d���&��Sxd�]���Y���Z��V��Δ�M��9��`W��L}!�%�������q��kqX'y����68�~��{C�2�
?ߋ E}G�)nl;np�p�%}�
莘������Bj�r�P�� q��ql;"���2�L���HC�����c�����T;~��?ld?1�J�_"�������ߊ�'����]����6�ɥn�P6���iya��� -�k�˳��J�9|�,CN��4�5+���VN"����W�.�o8l�V�f�s�2�Β���|E-��m�^~�;gxJ��k�n�%,�7A�)�4��<�_��쬡��N���x�����%J3�s�v�:ضT�CBQ��M��c���^H�Aw7OdfZ�E�#����Y8"���U�/d`v&d��yto�f������!�Zg�la:�A����}�V%V��V�6U2-���O�!�ٶ؂M�ڊ�x*S6R��K��1��)ќQ&����l�gJT��4?�%\�DtA��WNӮT��o�ʆ�U,J��á$LY����d��t�������x4���+e��a�6V�d��<�K���BJ�+d�����f�Cc�����O҈��q)�c6�I�X���Ƣ(����|��1�S��Mu�.G�mM}�K�NN��N}��s���a�����w��x��Ţ��<���s\���iQ�>pS{ٍ��ס�<���j㌱�eh.��<�p;]��ܟ��?TO�n#�M,ջr{O�E3�s-���t���Zb9�x���Q'��nA�9�"�h�V{_�لW�Z.���*�]}���BX���b���"ǀS��ӯ�P�A�A�@��z$mg������/|�dN�|t��K~�0%�~ ���P	ל�!�fig����`,�i_�Q}/PA�m�5ۼжߕ��.���%��t��W�3�IHe��������ܝ�q��M&�夆�h��d|�ؤ��t\$i����Ks��E��BB�s�-g�Z�f��,��
C�=�`���dY[���0�Ϳ:a�c�
W��]��Y��O�q�M�>OM�����8o�_�ݱ��XS�
İ1�}��>��û_;k"�e7�]�0ON��E��w��\��1��׫�ɰ�I�4|gݪ�x,�F� �^i����Ny��l�nʭ`����.�y�B݄��uF{���C�E�쬬�1�yIi�ƈ�o�hR~�ч;Yx���GP�*t��>����|%��UNҨ����"Hb�00<���D�ֺ^�k��f��:v����O2�#i��e�^����_x�3>� â�e�gx\ۍA~=���釰3a#�x�:	���M
b�:t�,�%��$?w��Uq��'��C㳰���sސ�T�i���W�w�6��?�~붩���4��`/o��>�,�L��_*i�(���C0Z+V�������ӏOL18LO�T��Pq t��x��.����X6�8&h�%?FS��W���a�Ѱ��O����>�y���F�0�	��`+�<�b~�=��-#�lW�fOPHFr���^�Q��.��� b�w>諣߮�di��'A�sDqO)�":����<�e�Q�D�Ke���-J?�`���~��h�;ta��4���O���#��j|��)�k�ͫg	��Ynt��|�W>T�6JD���s©L�u�eCz�S�Z#ƠS�U��L������-��6m��x����H��^s*��� ��[�5Ė"b���m\��y#f�ҿ0�7Yqw�����W��I	6O�玬f6(�����uӛf�+N E��{�	�iG�u��#��C i܆��Z'o��{��c�W�"El|�>�������>v6�.&�������
;Xn�S��ә�<��w����	d.D��S/� �y���7d?��L�y]�&��2���Ԁ���Z5'w����%EU�`�t�u��{t�݋� �Of�F�'}{�K��K{�o�Z�,���^�d(�������.���y�1kB�ȉ�@�gtߝm�k���.>��/0���f�	
�?�Y:��|�n]�]_^�����x�v8"�\l�>�@�
V�������rP�^�
�i��G\0�;%K{9Bn���~`�p/m�cnޯ#ރt�� ��uP�| �H�[h�/�����'Q�n0|�xGL$O�]� W�I�H�9&���z�o���R*n�I�zF+W��l�j=1��e"���6�T��p�����<v��ޓ��=9;�)b��̝ ս`Ul�E���Dİ��N�V�b��)|�>�@�Ի����������$I�/ʑ+ p�� ��R�嫌�VxO��z .9���M���`����ǌe�C�x{�N"�Y�.��b�1���N�bA�\2PgC�+.��u.~u�!!��ؠ�Zz�����B�\�?�?6C�_W���t���ѐDL�;�!z��VZ�Fπ6��0���G�!r�tHit��d���W1��2�$&�w-�Z����,�#M�e��n�3��S ���&ג�����2$��WQ�!C\@[`�o('��|�	���JC�g)��e"qu<�~Iw�;������H��Z��'�lR;�WB|����]��'��O�c*�	�ٲ���)���9'!.�^Eg)��q�5�-ߵ�kP[��� Lxф�Q�WJȅx�<�fҹ��Iِ�%a����'c}ȩo8��O����4$�T����;|��)$rٲ�0�3Kǥ3|08_�1��B��cR��Fx(�_5kAK~Nex=~�u�<�F�iN�z�K�gM���^H��~���a��Kk���Bÿ�]�����@�1�K�h�7�"�0�R�Ue���@���)�(���.�!)���K<q%9�$Z溷�!qŚ0![�M%"�gO�Z;�R��FUO�I͆�+�LS��t�[{�]��a>4��(�."�dB&h�tm�x�F7�97_�Adq{"qF�|%�z.�U7g%3��1���?�c����jz����J��s����CqJ�{2����.6a�ᔧ�#����5y5�g����z�@���N8!��5通>�juс�x����R�\1�}�٨�a��%Ԣ���A�<~�2�=p5�證Y��ڦ�1���K���7dil~V��8��xW6ˋ�&&�."W*f��\�P�a�eqA�6�tq18e �c�|�B�jJо9a!ŭ��FM/��4=�ҥ�|h31�.�\������-�������±@��I�m �D��6eP�Q~P8��E�^)f�/��#�|�6]��lc���4�-��+c�R� �"�Z9k�g��~�Z�=;YT��o�?e��PT�X���	&XV�A�/з-�P��%3nse������|<�׹n�R��g��'�� I{�`!&��e��*m��*�������u�{u�q���j�#���v@w9�r�<�d�{�!�j�!�R$�ק���:���Ry�R.sm���� �Ï�,�ƾ.����vn�(��$�9�V�Y�!�^bt	�6XP��iee}ǮS*I+�1�7o�ܓKZ=$JѴ�ǲ�e��R!L��F�n�g���+rQ��P�r����Ƌ�=~^����9GݾY;�k�渢.�ߍ��%>�`� O��&f�}�T���F��e�5��P�����)M��V̳����a�'��������E�_��"� gͬEÓչ2V�g�c�^���/�B�"[�K�����"���IO�9��a'z�� ��3�Ĵu��y1�K�J!R�9�U�`j��L��\�+�^��1���e���s1�$�(�N(\���%)���z���?\=�N���e���(D9�,��y���ۃ|dWd���F8���3��˘������J��3��+7%4 �H�{���d7��9�f�]&�5c�E��d�X��%R�xe҈�=`��g���^w<2����w9I��aw���"0$�Td#TBtH��D��t�5�OhˎNyd���_a��a��aqe�n��&v^ǝ�j��,ٔ�
<�7o� ��a��N@rʮǛ�E����>�nS�v��ye�=;Q��3-�7&DT!H��\9�/���/�Zl�ZH֘��?ύ'%ځ�c4��q1-�g7�w��0dY�������r%��8���]�B�����j�|	��|�r�ea���ʑ�,}";¦u�Os3ц���"�$�~���7ʅ������ɭ
��F��t�O]=�������]Sp��U�*WJ�D�l���4�|L�-�����-njz@W�e��*��}��h7XFP�?�#GD�Aplj�\�h�&�Q�t�����γ�w	��"�gr�/��t�$hrD�7_D0i�O�������D����Z�0��!��-�sp�}A�)ޭ�]\�/�u���ϻy�K	�5��2��ZG�\� �#C�S��j�[����?��E�/�n�Tv��}n	�(�P�긽;�����Z؋:,z'���@��IT={���8�=�s�7���d�qD�Ȅ>?������@�^��9� �lQj?=��Ѐ��,�u�4g���M�%��˦�}kr�khj��W���g.��*g_�	�<���>��N>��A���?>J���R�4���fZ��`@�E�B�3vJ,dj�_�U�d0ȇ���_�Ys�-rx����H7k�闔�)����c���5竬k�r�i��Rk`��3�W�?o@?��'N�"U45���e#�\���wup a�=H�^��� 1�@��1��Oښ��(~�.����|V{�'���)ju$vh�lZ4��Y#v+�۞��\���q�s_J�x/�����n4a��U�{+�a?� �%��"H���o$�uE#���'�/)#�J8Ϫ�^�2�� ���"$��&�aY)�Q��{��d�X�P�::k�JS��H�؏���Ak.�(G��6���#�$�i| e�� �8��h�0~e�c4R}�6 �xj��oG������6 �V�VLV����i�.!��Ar�����m�U]���1��JO�V�2d�h\�w>�R��M���'g@W����P�H�3��H����Z�����V�#T�<�!�~t����8q?M.}� l�� ����{@N����.OY�K����I�M��sO��
�њ	0�B���T��)bɄ��!�eW%j���Yc�`h(���-by�
&��r�s����/�*w�xVx�چ�rΝy�:v�{:�ן�\ż�9J.y��eٝ�}r�O�����e �ؖ��nT�y��Ղ�\4W�n��0Ť|��a:�-��Y#OFԢE��@][�_�ك˴�ZH�i��z,�8cq�݇VF�ӎ'	:��$}��ԓ-�A�@�ހ���X�>H�IB����W�^U��R[�1֝��?|Sw�c=�LEj�7��;��2�{v(8fϯ�F��'�T�a�T��3sX��s)t����+_��3��{�D.X�u�K�8?����b��� �F4ާ/8AW�v��μ�������e�d K�)�ٴ�8+&a�D	oR���Ia��_�*���aȬ��X�~Xm��+#z��b������~�N����# �:�r�>�p���f��1�r�;��5�;�k����򰸅^[�ǘ�s��|%2HE�D��)0�_¬L�Y��I4Pm,࡬<��+�I!�b,�@a��}n����LY�I@���tJɂ�ܕ;z�TN�x}�8��Y,8�RA���5#:mCT5�w^0���-Oc��)b�<��=��<�]@��SuFi���$�p�c>sqGDf��I�Klꓔ&S\���#ݶ��m8��zB�Fܒ&�d���cLH]^�	�h�A�jM��7��<�B�0奚:��D�´ .������H�1p
�ʸ�[��n�;cM�F/M��� ��<�H����!ڱ|���41 #m��}_jH�^�gd��� ��Z���]�{�R���
���8����q� .�eԎ?�0�LcA�����U�»a0����K���Pԉ�y�� Q�W�f�3D}�G��x���/ؚ�=2W�]e�Φ�O�Ħ���w�)�4*[$B��޿��Yֳ`���#��x�hwݑ���0-��B�p.��$�&٫���h�$��9� ������5|`�ry�ʾ�s�Ai�����Z�bp�_kLD��~����ryg�	*bE�h��SK�2�ًM,��>#�|�,(�b�>�ATߢ'���X�<�����4�\� Lr��؜ha�O}�fFp.D�e���
�J�j��Z�/��#p�ZՍ���Z@��E�"$�������U�ٛu��{NJ�?(8e��'��q�(A��2(} ^��fŲU��.~0L�"���	?��� IF:NgO��c��hN2�΅QU��P���3GhdA�H�l%�P,ͣ�	!œ����
�}a�\<ڞ"U�B7�9I}�$BH��m�/��(\���}��>;���l������U�:���0�e|u�Agm�c}�fW���*�'R�%q]���B�1Z��Yj���{H�9��d��w�G1����=���2�:v��dY����	����m.�����dDJF�Nw��'�y%�ܜ�Aj2k�ɻ�<ꋋ�>�����7�&������C3���P��\�qN��$��������Ǆ��	�Մ�}�.oD"�%7z+���O�׷����\�n��͡��e��VX���Uv���tJ���j��|�w:H�r�:@2�\ʧs�qaN�)yئ}$�
J�Z|d2uv�ΰ3g�Bl���U5��X���Q��a�SbW+׃��Qx�;�5��3�\q�XFxh �nV2#W�Y�p�{%}`Et��������Λ�Z�����ƅs�0N�^�7?�j�r���ʲ=0�WfX��߃��Ϫa�j�f��s��s��v�H�+��ߟ�����Z�A�s�xwgx�o��4a�K�:N[��[oM��[̅c�N�
ݝ�ߋ�ކ��3<��x����L�;���kC�XE�()(����)��$e��CƟ�'��I�Mf�=r��O��`��G	����Frx�
�.�\t�������[��p�����㽈�z5@ �ڨ��a��Xrπ�6�D�v�ợ��z`�#ڽZ����>�X7���bG�%��
`i[���F �h��p����m�2(��;q�J����'��3�NE��'�0h�w��d5٨��{��g����!���u8��桋Sp��gf>�� ���O��[�� ��B��z�kk���ĳG5� S�Y��[F�[���ڰ5C�a�1�;ԏy|G�_�k���܊ꋌ�w�r��ޘ�&IOb;�(C�ߨ]i�f��r2�>��*����)O=�2I�h j�b��w��Z��Ԛ̾�oQG����C��V������r�_��g�,}�X��**6�Z7#o҆�9-3Jv�I_8n��9v>�����2�t;�\p/K�l�T�̏+4�k#�dQ�GXm1��:T��hhEu%Ƃ�([�vp3��&|DjuZE)ӵ��{����9��o#�?�P���XR�
�a���̑l<��9T7[�ڦ:7���M�LM�S�g�.���:���d�VQ#�H��Fvh���r��Y��<M�^Z����U}By���!�'�V�[S��ݓ����t��S-�1�=`GZMo�6����C�����u�ѳ�	:C�~�^#v!˧�.�'#��`:��Aa�� Ƭ �Kߊ��a:��va��Rk��y�=���YA��L�E�{��lQ"�N�*���AdA����YvM4��,�g��7�y�4�E�V9a��^4��f������t�;�����D1�����;�jTp��]i�ΨK+I���e\�� ;��.��ֽ��_�֗���Z��J?ef-l�O�g9�h׼�\v���tL�ӻh�����R���X0�3O�R��W� ��nt��M�E"Q�>��կ�l�ڿ����0�ט�7��7�U�F{B!S1Sd�7�!a]��:�{4�����x�������|	� �}ێ�4�ڣC�F�u+������+�z#��?�?t8n����3�\(l���5F�h��kcTq�&)e�}�X�,�ߓWӿp���&�Z픑�(�o�2�5��`E�q�_@���&F\Q�*9���� ����>@G��.a�o͇��c�S`k�՛���\}�����f�>�ٹ��j�^-�}����ݺ��Ez��ZH�2\йM�0W��7��mvb�X�!t�Ϣt�r���j����6�[���[Kg����׊�_6�����e���G���AK}��O�̓�~��1cZ+� ����/�k��(�h�p��{��1,���l�J=r5H�5�;5 cC����؟-���rXv-"X,{/�����R@Q����v`%� ��l��T~�pƕ���ֆ�*���2):qhm��ˇ��T��H/��-���� ���5��x�ћ�����ԗ�"���y�H���'��Z�`����sw1��2�T�V#�y9Y�T���9)�������֭�*���o����N��?�F0����6�򡄆$1a��@�F���K5T-܆餞����s8^_&:Ҳ�Y�k�_g���@�pW4	��ʫ�c���W���i��K���q����>��i����/FrT�a���Yd�����L�rw��8�m���62Y �,�Qt�V�q��NvO'��� �
ew}�����5	Y{�3% Q�_�V���g�1�˫+�y�֪�Zi]����	?�J�y�s�5�b2��_q�Suu��MF��s۶ǩ�#��:E����a�RVA����}L:Y�󜥉ø��ZM�����C�"�f���e���O|zف���-�EF;�p���eQ� �/ғLȢ2��o�!����P&�Iī��o�1��&�Y_C�4E>�;S�Twm�F�B�_���'�Zcp�=Y�	9{e�E���T�P}���)ԫ��p*���W��x*N���e-C�.�x�`�-��zd)F-���{��=w�!�꫘1m��������y�H��� �6b�j�P ΂rWx�G؍��Y�[������z��ø��.��zj���)]oHo���q�@^j���BD�=j��['w?�~���s<�	ܩ�D<�<=U�92�Ʀ �4��	{�u�x������7.;/��Zx��MD�@.2��͈;��1]/DN<ƙ.B�ىDΘ���Ç4j�^Gd%"��"���>[�L�VRuV:�(Ī�[ ��� �UE���MX��A����]�%3�$+�=S���RIY�Znoa��3hۇׁ�(�)�7�>�O�1�������N ɮD�z�$L�e�E:x�o R��H�f��k�w���@D��X�a�<�!��p��r��r0��?pPP�1�^�!���d&`��� ����$r�B���X��'�k�
�L9�0]��;�˽��P��i:�����x�+t��L�����ʔ��i=h�N�mRD����u� �.�I��K:��bK%P�o4�;!�^<����8~q*�:]�}:{@I��vC�L5��R$��	/��&���q��b׾�%N�6������Q+�E���NI���gt#
�s�������)"/1Xq�5B��+E�߽�BL:�K��|2iM��"��1� �S@�n�6(���3%�Έd#����4�}vz����;��\ď\��-���Լ���NX�'��*uw�qH�x �/��%�;��E�G�#�9���'z�%zG�p.r� ��*���R-�=�a������7;��N%��FR$��dZ\K7̱fe�J�S�����7����D@�z�̤����`$K��V�T�?P��>	���aiB(��u��n��X����~�����_.�1��S\h��F��Fժnr5�c^4�%Ʉi�>�7uz��E��>F�|_ฌ�f�1�+�\�*��J@�쿞�F�&��㌿]����(,��H���(�b�W>ki"p�o�R[�<�>t+�)a&SW�Z:�����@wf7�B�|��^����,��Qa�׾��������*���d�cD�r%Dܸv^Ix�؊�/�jΎ9���H�#	��:�*��('�p=���F���a�E�
v�e����~��u��O9�-�{}�7�}2w$��B�Ԯ�\L��Y��n���fl*�
R�=���4��ڱ����'�}��&K(n��W��>t�Մl��!��`��*�t�L4(�]��L��;�+Z82�H:�� �I��')1D�Π>�F��X.a�r���1��n��%v���.ٵ-���|�DTJ��/�Ua���Uv��#�+[`L�1�\�Ml�(I�B���b��i<��i�*�>�����X�d�l�1�M6��������q��C���V�^�w&af�A���(���D�̲�@wP�!���/TV��XY�wp�O'�`ds�[n��)�XKHz��YK���s�S"���h�r l� �\e���	+�g	����IXS�_kk_u�!�Z�ʵ-ܼ��ǫ�~ƞIӴy;��%�15= v����1���1���`+��>ro����5ړ�V*ӑ�E����%�i/]>=��E��%d���y���p��q�P�S82�>�d��Σ����� "��pQL]Vf���D��R>Q��V�.�^�vud�	b��C>�κ��<��zX����]��30���ʹ�o�AZ��*��#.6�|��W����� ~Ԭh�VB�V=Ou���f�dl��\Y�|����? 뫈�I2C����bw��+���0�+*k�^᧩k�����~����di�|��޳�y��0P�<g��>���짲�e���`�g�0��SƓG���;d��)�>����W��n�)p|��5����io�(?r�.d8���(�!������t���cL�4� �0��%���R� 4�n[�v��x�,��ێH�e�����T�2�ƻw�ku���>�������ZN˚\G0�V�U蛈ǔ����,���<�b+���`�2w�� =���^,�Tp�����������$�2e�!����h]�����Kge;�C�jL~��-<���@�Z΂Q҂�a�i�2��vp����
w�z2�zY�Ι��1�l{�j�K����q~$�Fx�I��	͘*��<2��ͰP�T=�
9���A%��i��G(g_h<�����%ˀŢ%�*��Z+��� u��r"�&��8�F��)�^���i\Rv�W*��u\*�]AAwU�����"�}{ْr�����4��`����i��^c���~e7dA%�0Y'Y.�c� I����tR��oi�L>���)����������X΄��a�r�V������2�����$_�]�؀���9zYB��tx�}�A�G���q<��j͉����	[�{�d�Z�6����"y�@+��x~�|WD��-}�Ł�(<fA┹>���WQf���Ԑ��o�D������I�5���࣐ӘT����T��}���E'���XW�6Ny-�<��Y�Vn�%k���!@#�:,��)��ʤ�3�����m,��$���:���Kġ��+�:�����ȦV�Hݔ��0�JN��(�~R�
g�Ϣ&^Y���f4�xu�顠V�F��&]H�S��=��1���@z���l�&���~��E!�4h���=ɮ�4K��n�;WO݄zYuك��~�IJ~��ay�P�t\c�'Gr~��)�Zkz�T*#��H����M��i�8Ƣ���d���u��/����)���w���b��ٝ꤂�5\�0| �ƚ+��7|�=�ԙ��7ɖBM�B8�W3R��Qb�՛�������m
���!8O��)���J�ru���m�kТ�C���X���[&��t��;#�E ��A_䢿7VT��җ�r��.�
 ʽ�}V3G_�ͯ��G��T�_H��eT����k,������9������O7[b ���n��Ö,}A�������<��H���������<,8;�5�gC�a�"y�zN�����U[�W�ޛ ��5?�5"Un�ξ�9�AdQ7W���p�C&~�9 �(H��ӥ�y��a��޼A&�P�
UC���m�����$_���h�r�Ƒ�⵷��E��eDXlv�2��P$��?Z��8����1}�+D>-������$(h ���<K2)k���+��W`��OA6���������i�y�wd$�s����^"��*W��P�%�U~�B[W,�겲5BIN㢬[R�Q��l�>$�b2�-���±D{_� ��no�s�O�>B��2c�����ɳ�ЗA�'0I�v�[���:��$b��}����P�e����b�&{�w�䑓3M�-DҬ�w�H#L,e��j/Z{�.�j2m��Tr����1��:�#��~�@
��UzVGc�NK�G�kU�-p�ڷ�y�Z��<7~MY�l�%���z������_�"96�5zt>�4�$���9 �h,�}w��f@I���g��V�Eq`�ˣ9�~���*�:;�Ǐ��,�F��7 F����N�.W$c"��d	���i�v�`D�2o(���"(����sJ��@����հ�j�;]p��wR57��$i�|iT�� %)ʼ�5k
�Zm�`�j��J��٨�S]f�݈_O���	+r���;��3S�DE�����	��E	w��HE"X3��@�. �,8�̧}�J�t���~c�k�k:�]ܴ^Z��y��B�;��%;z��[�4^��b.�v�E� '����[�v��g�e��+��,L���o �2�u�&?��"|I�.~�ʧ�W�Ľ����2w�7s��3/����ǈ˵2(A�ՍP� ���=P���>	ɿ(hr#����>
J7�Ɣ��uJ�������6`�t�4���+~��������_��H���Qz[�ߔ*�q+ڰ��EInDj4w��p�K�����-�}��O�
/7���9�h���l�;�� 0ƪ��:�K��5���j,{r�z��c�2���H*�Ga��ɾ�
�����R�<ˇ>�M!g!B(>�,9 k噎�C�T�#aȬ��X��{��a�{�v�m�:[���㟾�ת�c�gKL'�VLS�1��� �8uJ��S���ie֙*�@����9����PU5.}�� �ȴV��|��{�6"R��ca`c�8[��K#_4�-©�50���^�P�PP��nĿr�wAd��� ����!�Ĥ�T۸�]ڷ��_��������g{����	�g�E
�{����0�\��B�[����_���#�J -:쌯�&��$ښJ=h�9������?ǖH��������L�#���>!����e"bh�F��v��^��UE�w܉ ����٧�IQ�SJ@A
 Ã��X����F�叞*�F 4�ߠ�1�P}���ڔ���2;\�/�J+�'fA+�"*:��������w�Y^���L�k;�0:��z��f"���S��LQO�V��PpP�q�7/��͆ 2��h�$�>��z��-�ʟ	���rB��}R@$?*2������OE4�.o�w�c�M�kfk���"Y��jU�����(]-w���t��!���o/�$��r�E{*��P�d}�=D, ���a��g�R��!e��+	 �g� ۫������e�Z/T�O�=�)`�Oه+GxΊιJY����������k��o�W����9YwB�89p�)c��/�z� �ρx��GK$d��+걉�x�S��0:�y%v
g�B�=��E���p�/l�����u�#ʜ5ѱaj,��f�����iFdJ���S+z�Z�E��ֳ���k$W�g�Q��w}ϛ�{T�y��dH\�9킱��dğ�Ic�a炊��#��m��8��Pu8�Y鞟% b�̸���ۂ1l�Pͅ��'�׿��v�ޚ#���g(��<������l�d�B<��[%׹���]:|��"��[��Z6�<Wo��5^\��r����z�k�	��$���Eo�i�tEW�2����Xh�� �`�K[T����Ct[im���L�n���Q��F�u;��	@G;
�Q	�޷��0~F=�6l<y˳����x �u���OFZ�ͽ%$��̰W6XtU�I�?�&lo���I���m�Z�L���z�1��4��o�J�/QLZF�gU�C;���X���9-ӲO��R��|�i����R��c]�i��x�˂OP�:��������/�קNy���ވǎP���loC\��jlrl<�R�G���goG++-�wċs1�^S��O8�����Y썿�l��( �6�����;�� iz�;�!C���g�~i{Z&����q�����j��5��&� ݂<�-6��=��	�d����
�q����;
��>��+�*E�uO���=��G�*�	��7�3����D:�'��ll��au�ƈ��9+*�Y���n��/�D��Yt"�T������KUzKe�19�<ŭ*��B|������[&�+� �@�KĔ��8V A}��K�1U^�HѰ��YV��vݣ���^ X pˈ�R�
k�:�{H�4d�E��*^V� `�#^o�5.�g���y�V���p��U���:��ɯ�u37P(�t}`]� ����|UYd�X&"*m�	N_�˂�pb}�\/�K{�;�?O�c�q:.!�Th��X���v��UW�:�����(����<Y���%�o�fg_���Q����ۿ���};��O���Y���t��*̊YԬq�^��=�>���ʴ�����g�Ү�H����в�n-��5�Duyg1rH"�����Y��82/7�Gf�9ϐ�o{56��}�8q���Z���>�/����<(�&~���tL3�3"u�$��ysFU$cDeG���@���I����5��\7�|�#�:T���|Ӝ�hB�S�~���b-��)�:�;��o���M�M��	i������q���:�!���ݔ�"�^�[�\�չxc������$�$^���@7D������f}��4�5��n ����h��%�(%v����k;="	%���ɠ��AW�	�1{+��<)Q5��X�<�̣|w��:t.�ݮT�y;��~�?4���b<���dru?ߞ癏IJ�:�^���'�=֜���cy�L�_i�	E�|[g�4}��A��𷻛��|�M+�S�O*�Im\��-HO�,�'U�(����C�b�M2n5D�p-���y�
�%B2�j��H�=���ey%�FȨ�!Ƿ1��`4�6&dTv��5��B:�nN8cw~�i��Ȭs�������KL̵��R���1Ĩ5�	 B�f��@iW��nB8)�z�fOl��x�sE�&�*�e
3+�)��'K����. ��B3{��yr�����b�it�{�}�(���+�d�a`�p��	F�C�ta�H
�H�`������)ӨN��W?���O��]��Z��B)r��
"��~?=�5peԔ���<M"��QS'�u?�GQ�����߹�zG
t���k�̿��}+G�t��	׫�&K�^IB��)����xV)�)Z�����sn��o_#�0�>�8Ln����e��������*z��� �	 ��Ǿ��|�� � K�����|ɷB5=�n42�b���,��>�&�@j�vs&��� (l����v'+KA۞�l��_7i�����M������e��8��|�k��&��N���l|?_O�l��P��,k�E�e-�?�H�.������W�s��JQ%�����Dk\<��}�sI�n�D�b�,����5��u�kO/T?�'폈��G�[P�m�'���Y���[7T� ]�p�8��b���<ǀb��-�Q#� g���.��^��1��T�ߵ���1ӌa�?�8�\�|3�Xt�'�h`�d��)�&Wd]I���
K�+*rl;{�*\?��HX	�<;6��Z��7L�|vv��n�@b+�&��S���0���S�g�c%u\0�{0cU�����%�m��S԰�屸��Hq��1��pH`��T%���_��$�M��g�ֻE���>"��W3/�%S/x�<d�̭>�fFS�"�\�_�QLt��O���y'Z5�7�i�.C�+��P�[(���y��:�� ( ,�2VN���m��L,~O�Jϟ_�t�������Y;˗N�$��8趭ӳL9���7'��(p�L{X�������r�jʼ�DU���Z�A
�6�G�TjϷ�*��ܿZ�wk�u��2��HW����GG�o,^�e�ÂA�=�6$\U�q^B	~Y����C�(Z�|Ĵg!�t�[~4�����}���x��NamݡZ�EF۳��M�v����L���\�M����$˙�_�tXvC�%��6�;��gav�C���/-F�  �)�^�(�e���G~�we|{����vCsЛU>��5�W+wkM6*�\X(0���%���f�pX~�ӧ�P��I��R�:2~X�[6e(����'"���r���{$�U�~�N[��Y�?kI�f�mI'�[j�e9�.�L����4L\�[Sݯ5���ӏ��c�WN�,�Ƨ&���'�q^ߝ1@����lQ� 6Dawڃ���9�quRµ�%Yf*dD�qv\�-���Z���(��^- j���op��l�Pη09�'�t�Ӝxn��Wy` ���c�E;|���g���'~]�7������F�%�*���/��w��D0�`7�K��?
L}�u+۾�x�O�d� ������h�`���\�_�ٮ���$�4���f����#'\�o��I�`r����!�7<O&����i'w�#����xEj��R��������cn[�����u�:���Y簣h����CV��Ȫ���K�ɒ<k�� �,�K��4W���f��5�nb��Mg�Y��ACZ/1�-�*,���f\�1?R�)5AlmO0�,M*Fj(��䐰K}�z΁��p��p֕�� 6!TX�:�Bӧ�u����K�X�/]7ri�Pq]U���!�kvQ�%�H�����__Qj�9<H4CB��+�/�gj�|�{�޹x��/�563�7�j@,Υ�����{����7�]�.�^<��oӛ����K����}�e���Z ���&b>����H�ߠk9�a���-O��r��z�s:F1�~Tv�Ty���"��pqW_�6�[�c�%I�Wb?����3����I�R9�@��'�F���u���Mk�%��)7�Lz�r������u6�B��h����y�p��a�mX.���y�^�ȳ�(LL5f��'�5����H�)c:2&V�ejfa�}ɔ�� >�n0۶�ֳ
�8R�T�U�|.[��x.�m�
�}�Q�)?��b�1v���Z�8��&����uI=H�YP��9���%J����t])-,ƫ�ϱl��{��-(� >����g�Ǟ�s��?>5��s/��ƻ{B���z��s�OM�!}+a�f� d�0��Cm��0bJ<���a䯛���'�<t0�,�&�| �Bt2����H ���T����{�*Hu���p���Y�`��Q����_ӗ�±�
4�2��jafí�rHzj΁lǏ�I�D�?�����* ����k΀��̳w�@H���ڄ@�]Q���ɒ5"e�އ(�%=����"?qz���� �����]{T�Y41H҅����z����
,��6�c4k��D��F����f/�^��� ������f�Y��`�h�S�AXn�jC�Ӻݴ�~Gز�/���lE�Ya�����-(�xS��B��#�dƝ��}-�cO_`TX�T��܅�_�؉�F��x�!��1�P~E@:L���z���\�T�:$��_3��	�S ��9\]�a��_cEW�|+W����4�F�|��}eA�jʹ��̓q�0݇�