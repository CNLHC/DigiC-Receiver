��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���8}6l�����^z��=j�jD�����jM�P\6�! >-\�(���1l�W`Z���mKr���4}�H�a/�0MV��-{�*Hq�h��k�3�8?M��v�c����\E����G�+����Z� :� ߖ`C�dVξ��i$4tx��r��υ���"�޵�_5�U��	��N0��՜����>6��!5�UY��^�F`��>���|�L�:FsL6�G�S%��:J�j��q��FU�zbl������_M�S�fqx���pZ��e���h������̸��rDYr�JA}W�]c�I��aڃ������ �T?	۵��E�b��n�Ž�~�#MDp�g� �����ǋ���+[�� c͐CSQf�hP��ڹYƳl󊌘_�S���H̭��>y��r	QDF���9�O�Yx���ZV�I?�+v�޵�%r���(I�g<(�)�!�*1�[�P8Ruk����ccp��۝g�a�|������yB�號v9dͶ)�ay�g�!�8�
o�p�x��m��l����BuS���s�l�+���6o����K�j��-=�У�zʗ���"����Xffs{e=�#�ZֿJ�\����1^.Ǟ��K�'q��.���γ-�9�)�♊�l��:���d���A-(`���ߤ��"���|~��"�]{*�V�P�E����C����"�Z�� �H8B`��W���k�Ѻ� �Q$�~0eMv|c�8�(� �b$:ڀ��R�I�Eq$.��O3�]K����9�ׁ��6ɽ;ַ���� Lq!� �ޏ��-�\ ������kMXR�T釬<ߊ$*{d�ĵ��R��RK��K�Վ�$���<&פ �%2Q�x%@��`�� yb��+��/����l��t��w�U7�����iҜo��0S&)~`� Oܭ�7��n�����Ǽh\+��5�ӿg�*+'M��Qv�O��x����Kc��FO�,l����[�6�^ɍd�q׵e`��lQ�(e�$H�l�k?Y�'d�4�N'�E2�ռ%�V�Q�V#֟ɟ#*�đ�C�.N3I]�Y����:Tx
:�h�u1������Wb�=VG�( >8��י�¯�O.G"��v��������a���~��V�WL����!уi�sB0���n��ع�\�\�(�0�®3*Y6��hU�1 a�$�֔����7��u��,�\�O'�o�C
�T�nfo�p�G��O�;�p��G�|a�e�Ks�wyL�B��]*޳L[U�I �t��7��y�+S����3���h��M}5X��'����aA�W�MA|w�Y��&��l�cUK�qTZ���N�P�T�N��W6>$��׈�N!�ϟV	4��D�V$�t�C���Y#s#���뼕�V�� �*6_wf�j�D�Ex�D�"���!Y�Mg����O��8�j�3��J�Rjv7����؏eI��_���(���.ލ��C��=��l�*���+�U,b���n5���|�2at��l��/�P�'.g2t��)I��H��}:="t��L��|YN�Okƚk0)�97�P��16]���F'jX�Lqd�ď4W���؝~��h�����R"o�����D����h�U7����E�)�	CO'��%��2�o����D2ʝ?�o_U,��@��X4<�WU1�D���J��"uM���C\���&k��c�N�QC|����M��_d�ߊıs�Xm��_��p�ɗ2��4���O��r�͛�s�	Ͳ��}*����3@��f؈������g��&Թ�16	��s�[��:;�T����]��+��x�ǚ���9��7@���]�[7���f��Q!�-^�U挽����i�9D��.@+Y�0T���Y�g:��;�lc<�~���y�cC���Ii��Of�a	�D���K�1gb��D�ʊ��w�M��^���Ti�^����IP������b�*F����Ds��.m{=ٜl�f4�ó�1����Q%}w�a���._ug���w�S���g�4�/t�V��j�ekPF�.�TH�H)�9M�ĥ�>{Po`���6������Cl�z0��p�eH|J�RCu�h��O��5��ވQ�** Q���s�Z5#pnK���Y���H+�8Z$�x����J]r^�	-K�T!�T[$>�����Zy�0���: �uK��q��~YT�b6�K����1�U��FS�}՜���b���8^��VTj�9W'(���? ��r�*N&V����-��D��5f	�^e�ʟ���-�8����?�ۯClق���<F��� �P6m�/X��w�@���n�H���)��Z��J�UJ�<��n�q
-,	©�W��#����$�0{FZ��*��!��7K�G\�{��m#�Sir���"���� ������t�+0Ij2d�K$(0f�� ���8HNS�P{=�J�63���/�qW�K/E�����9x��(���x{�r	JUO��M�9��I��
ƀ�3�O'cW�$*�\���,!�2��0@6M�}7H�ޣ=�t,���*��1�;Ҭe�vȫKJZy&�,�Q�����"�6�&�3qЦɟ6��H,��"Z��砊j�/M��'
��ηM|̀ iTB�CP0���i��rf���(�b��TC2�=D�a/�6��V�lI�@��J����p �l/N�@�����`���3�d��F)���!��x��Xy�Ga��.�9�� �
'v�TY�G6�(�^��_C��|����:1�`�fk���ܛ>�P�������Ҁ��+�����	��L�ϯ��%�R��zň\Ys�ܲhW�y��ة)���b����z�O�NT_S�f>�ՂD8�����r��fXzt�a�NՎ="���>Ե����ڄ�`)��t�46�1ż����y���' 䮜�be�])W��o��L��nڹ}#���oj��ɚ����vY�n�3L�9�q���O�K�ąx$�{��t��ZɢY�47�b3���p�<�2����2Od�mJԲx�b���F�����v�$�GV�[Y��p�7>}�i� o] ds�\摮� ��EΩ ����`;��q�������W�C��G���>��?��gL��vUa��|/���SW��a��[z�I1��pҷ���߰v(��F�K���\�)�J�ˬ���菫�������2d���ؼ�J��[�MF�\r�rmN;�%$1D�⫮`*�S� S@�QO�;n +�@[Y6��T%�0Q�b��q��$"����g}JK���"�2�DW���G��!����O��緈 م4�h�p�GF�8�u$L�R8��-H�+��z`�����������5Z�R�O��
E���(�u���`6�߸ib;�Dc��D���n�/r��}53�ᥢ������f��&�ꋽZ�4�S����4���k��,�o�y�զ��*Q���;;��x/��*�[t���﹍m����&�뮲[ڋӴ�LPiZ���ϋ�qՔ����Q��R)gA9'��!��P��ۻ�u����)>8��ʌ �f�i�����`�<;�!�x�f9����{����E���4>e�@�X��K��>����@���G��$>�j���
*���G�(��q����<T1�	1�dK���&�ؗpw� սz�ݠ-P��fW�t��:��#;�ԑ��c���P�_�P�2FK�b���hV#����i���>.F��'�X�vM���'�m&�%��w�9��iw@-�#���f]3�����OO��o��|�LUg�3]��v����Ql(Kҹ!�n��'y'@E����D̜��y����>o7�r�B]��cyT���ݦ�iE�s��U�ȩ�����J:>{�8#�#�	��.��TB�ы��������pB��*��c��pT���H�[e�2	�3��q!�*�G�ϼRo���|�v��� Sw��\4�p��VE�[	S*�3f3Y�6�؟��ܱ�%9�R��mF���h˺g�����D�'�wvtlPS��Z���<y[W=��Fd�^d��t�b���ZֽgB������Fj�5}������J�O��uw���(m�"�>x��.AL@?�hڮ]����vҟ���!tj6g��ٓ�����5�p��U��R[�U@��
�yo�1ŉ�Z��ff��G*U��`9��j�1e��:��´��M�Mʧ�nȦ2I[��A��l|��OA\�ۋ�Ap��y" �(��e讳,����b� ��3��JH��TʖX F7\�j:���p���N�����bƶԠe嫄�%Ҡ_�,�7����,<%X.a#)��-��\+���zљj��:.�	2��(�~3<�7�u����f=��s�%Af����n�����![����#�tާ�*�AdO����y&�^�'���w0�P?x�<�~z�݈E.���EC��`hecPys���rM�x���17Ͻ��ѯi��y:޴��<E��o�u6.t�Z�ֿ�=��+��R͖�{�J��Q2>�Z�`�=�`��,¬��>�WN蛈��~�Qsଠ�rZ�${襌&�)���>��F��\��r�����f傃'=%�ep�F�gc��%9�u��6���`�ȯ2)����El����`��$@e%�]���<�՜($��/䷟����
X���E3��痜B���kS%ʙȻ8����ևÏ��!�6�Gyĵ�E7�S�<(+7@断i��J77���_]����x>H�/�����5��{J�J���k1���_��+�>߿|���+�j��)�e�H�x�7�ĩ��|de~�*�V��oY���?WE��N�f���������߇g�Ey �?7���5�q�^�̪e\�9%zײ��/��Wy(e��ܚ�����?t�ژ�S2Kɠ�F�>�ʞP����n %��̑��{�X��������X5V�;�bIzlPғ�3S.zp����ӻ�	��Qy���n��!��ʤ�]g�{��0+֑�0�%w�u�>��������wι��o�{��L���<V��z�IZ� /������č�θ�XaӜ��=M�zѿ�L,֨X��ia����M��J���tӄ��ʺ�wCz!BYo����*�Z�	�3_2>���3��u&�k�	x�J�7�QŜ1�)��^�:���)�!�m�_��Jo�6��f|��ۑ}�B�[(�7�+��*��"OC|*u���e�d=ֿ9����b�$��E���N�O}�C׋r��
xT�,�@�|�l� �z�.x/>|pT�l�#Ba���J4o #�࿇�)��<�6��S}E�>�ׇ���7iQ������y.��5�/����b�&kw�m�G͈�++�M�+��l|�x截 ��1�KՅN�;(,v��E�B�'"=���RJUR���[�4����=���0�ͳ�Jq �N`��oѓ�x�'������%gB(�Ԛ��f|�ˣ��1׎ٽbb���kg��VR��lQ,mu�d�����hs�Ъ}P%"��ig�s�ud=��S3t��!� �	���j�X̪���J�Rz���!���,�,^�r�zY.$��������$�pX+?o
��"O����PI����T\� ��8
���;j�82z!:E�U��\8?�r��_��>1܊�U������sT�y�P;�k�L�K��<����B�s�b	���i�G���|ı��:���!G��6��h"~`��ʟ�c�d�ۙ+C��#��U���DV�Ilty0��>�?'�a.me�S�e�9����l�ao���sD<2�P�z��0x��E���}_�u�@'�%����xJ�<�������E�Q��!Խ���Z����؎�y�.� }�Vw���~�Ǆ�8��4��E?�H��q��H�~f���T�� �|Ұ�dʣ���>��	G�͗�7br�V�z^�� ,	X��V.��LA�£����W�_Z��`�\���m�f�m_��nS�Us(Iңv��z^_�y��\�ȗ��� v�����ɱ��mY�i	�X��.cǽ8�52�ɓ�Dh�Ao�lΩ�W��;6���*I�V"�Ä$R��W�v�V~�Kn��9�`�1��W
�n��9Z4�Ü{�f�|M���m�IH휜#�k\�GC���X����iɱI��d��u^FS��قU���ҳn� ���-%Wg=��E�"�#��N�����W���c`��y������NNd�2����rMi�h���m`��9�iH������K��z=���=!�pW"��쮧^�L5o��,�8���gC(�0�`�l����Q�p����<!H�ϝj��L�pgf��L�flx�{�4KL}�4��	9�� �L�I��o_�wݐ����&��}w�`ݯ%�(�7�_�M�� �i��ub�����T���������ŵDFusہ\�����i=!��Jz�8��Y����,W����������K�K�T�C�==��%���@T�I���Ў6�h8����NH�c�J�&Y�����0���V�^$�l$0%Wt0���_6;���|�����m������D��\l��@��xp��f�6�2P����~M\�~�X�Yf��B�Z������Ce�y��?���H��Kj�Y�;�<��$Y�W]N��.�mF7����(mX�K_Bi�e�OEW���^�d���B��Q{d+4�ko�]�&�
��E�1� 4{�ۖ��{]������x2. ��^�È7�՞"�>6�
�p�|�~�x�P����z��Y:�f���V�fO\�)���&�o �ja頇e�:Rv�2F����h��bJAk�Z2��u,��|�v����s6,yi�\�D��9��%�(���K3��XY�=��K�i��~��/i�	��`�z���߈��wC�6���Nr<�u1�}��D�����#������o*u�5�M�68�R]-�S8���a�J9�h��q����Љ�_�����7`~i��zz�<�^¬-��ެ� ���۞�,�
�p�%��z�+�Q<G[��T��~w�MP��6��0�ǋߜ��> ������E6��j�h��w1���0��H���E��z����H�ݎ|\=S(ZDcy�B�Ox�a�ﺏ�W�'R\��,�
�<_�������g�0C�"-/;%.h��A�3�Tt���ͭ@SkdAko)�OVE������f%"�%�\jD�Gr&��$HøCw�	�\�����������0ۄ�5���S�%����>B��8�@�~(vU$F�,T����R,{�Am鏦���X5.�͔��=��O�s��+�����nk~7`�?��,J8�]���͋�a�X���Ԉ���t���Dx�����b&�V����j��ʕq�K�J�b��F~���6L�Ky���{�#���E{2�P ���qB8�qG���2SL�Y���!Bg@�_K%,���u��x?y�`S2�#�I����m�@���_��x쫟'�_�K�IA|N����T;	]�d<H�
;:�T���H�����_0=�;�j6�J��n����HR|��aN�ȧ:隻������x���|>�38BE_ ˳�jE5���Ltd�t �S�C���9@���i�3���I���"�w�������P����>��p(a��&C��W��B�ٺ�et���㌑aI� nU �S}��7��b�3�T����"�|������l�D�G-��~Þ��!�+>kCdx&���n�m
���ee��IhZ��<i�����~�T���g���p<������J�`Js��B9��(��o&�n�� +�W�%� �R<,�6	X�r�8r�ڵ�>�RY$0�I�x��`�B,�z�Z�	$@��;���ϯ��C��������XW���+ �?���o�[Wg�W'�B������s�D�yR��k��!��zkZ���w��q��.E 5b��/��T�R��N	�1p^���x�
�����q҆i�7@B��$/�	�C�S�t��P�jb]pc椽O���Q��-�nw7��q�6u�1B�>Ȅ��~[��P�Cޒ"Qk
T�������X�
��1"��.Mz�:� Le�A��	���܇�b�hH�ul�U+�����?�	�m��8C�M��'3E��]�����i�~�^f�Aꃔ���v/5�-���9��e㥃���ʧȁ;_,���&�C]~�:�g�\�b~dY,	���s�nd�hHxGiх�o5�4M�EP׷�x�ޒ��-�sB��mE{d��,�k5٨r]�r|�L��+�. �a�L��j�C��"�K��m)�$gC��r���*�p�D��b�7gv�K0˺+y.�-�V�W!�yDI�1�����t\},��Ywʭ Ԝ
� ��M�}� ��R�fI�,�r��<(.�=D]Uq���β�.�tR|�۝fgAj4�`�����JBS>�(�9=��|xq�>[ω����[�	���.���![�p�m
>40���B�����y��_Ln�"��r���v��p芓F�#1���0��@��<��xr������~+Ə]��t����灱(��f���X�E�>6ۀ1fq ��.]*�N��_H� �"fIm��C����a��� jW���L��x����`�L.�{2�E�K:�^#Q�.��|H_~l$�:��T���x�m��j�<8g�:���]�&�<'oi
Zĕ%��+%��X6��� ����� ��o�;�"�	Y�����\0�<I4a�`Z�_��{�P�D�;&��1=�ģۈ���������܃V����){NA��k�u'�]�n��$��F���-β� ��@�!CC���\28���}�?���Ԃ�֬ɟ5�LFpw�,^B�D����KMދ�-����Ɍ]ϛ\�@yȬ�q�<�ߢXn"*Y�_%H�n
C���(3�^#��ܻ��� �|4( �J���N����55��#N]i0�޿N]D�,J���gw4��1w�~�C�Qx��e������hy�!��Q��]R�8�'\�9A�A�G��G7��qI�a�5+��jk�l�U��4{ؓ7S�#��3���4�𺝷U~��FLؐ4�J����#6�T�:g�
)s�����*��)���3�V$�"�
�&#��9҈J���\����g��'f2�����.w� �8�����+���O���r�ݏO���#s������>�_����Ѷ]b"���YǕt����O�6{X�8�y�6W�$a�]g�{����ʠDN��N׶腤�z���4U������mW�@i��
-��N�{ar��1�\�,8�����F�i$mͩ𡽺lLC	ؚ�#R[R�^�vx���eʪZWO�ij]��(�����|UtY>���*|����2@ԅ�rf�ʎt�wO{w���Rf8.]�S[û6��� E�"�׏�Rڕ"�:ǽY�X��b����,B�<� fbPO��x�v	q[���F����;B�
�w�)]�5�; #�@q�(����'z��2x�+(G�6+@�.��n�6��>Tg�x)�s��5�\��(���a�����\��+�r���Y�l�wret�=;ʼ^5���0�@�ov;オ�}�E"ʜ!dg��/Ɇ�[p��i��b���p�зKY��$���2��OA�|v��1���GX:,c�0f���$�q"~�ju)	67��f,�.�V;~w+&�n�kE����̺vZ���I�bW�b�CϏ�B�f����
�'I��*��
<�[.i�܁4^$x\M�	����$L)�[���K��n�'I�Q%�*�a�.�t���^O/��+�V�X��Q׭�n#��?���6������Y��rLD^ڦ���D�3��8 o3�Ђ[����u�bÕ,=,�.�땺~��bv�J�ںw�l���`�L��q(Z�0*���K��.]��:���� 
�秂� �J�ϱ��z�����B��`܆�G�0L������p�k�[WL�H�b3�4O��>�s� ��/�b���������H\��(�����-y�'��������P�CYLO����Q��?Ӎ��Tt#~k�����h��9G���|�5z6�R����X���DE=�B�(����ϴ7����t���" 	��
�j��5b�+t%~�DW�֑�骼���^������<��Q
�`H��ԥ��R��8�ݚ��S��,�D-U�¶�|w�(����8��&{-�e���OXM���q��6e������#E͗������{s��ʇa�V��<����5��,�俸4g0��,�"U��kC�y����b��\����+�;��!�{ą�����ɥ�Y�+���b��S[�4�y�泞���{ɣN��7���<�#�~[���N_���:3-L�b�R��L�d0�>�i���U�A�ds=�c�Y�d�/�@t�/��n��F�%w��Q�!e�5zoN�(� �_�i7�[���9�^�Y6�����~����6�#ƈ������Q�Ι����P߳|���4�`���u�5�{�����Z�[�e;�C�Q`������~j�P;�Eq���n��z�#z� �+��]�]'Mw��Q��9��
�u���Dv����@J5;I��Ԩ��&���A����'9ؓ`<�v?�;i���������ƍ��jl��{9�kq�-��_���]�,�7�f搊����%�[d��?*mn�z@��M�h��E�Tj�����j���� qo�Ӑ�	μ�[�j�wu�rbA�������-�%S����G-ָ�^[�ٱZ�_��eA�� \������{to�k�(v�;��~n���b`��m%��s�'�Z<�������'6����*؝�P���X�XT�t(TZ#R���P�đ)�k���({q�D��͡�
�5�p��P�+
��G�u^���g�Ta�m��ꁥ�<BO��a�Y�N\�nA|8�W��X t��E8�d�x�\}�dt5('gL�Ʋ)�G`����_�R'�p<���� ��Z�v�P�d'�d0!?]/�����X�Sn�f��{�:��9)��Jq���p�=���֢3a/��O��F�I�|���<�~�~����+�����8�5f
��m�N Ě����m�|� Z���m���6TC�=.��m�m��}g�T��'��HJ����F"N��
qc���Ec
e�r��1���tt�4�	�0��-+����� V�!��Sg���f���[��#�_`Q"pߑ'��5A/��z���a)vk��n�0yd��v���i�f��t#��r��`C���[o��AHFi�.�t�5E��X1���*�ʷ�����i�lqF�!��AP>Go��_z�(�W���V�N��0�Jc%�Jx(��ikKy�;���1�~�3B���̪��ۈ^Y�V*%8�U��$|�1]\�6.{�VL���r�U� B>�^������`�n:��@��Q����ҌFT}�wkȝ�o$h����'�,5#�v�&m�a��t�	RQ`�NHћv�/�enr����я#Rl�P�N�����}U�'��o݈7%d��QC����H�N��4���+�̔���S֊ﾕ��
;#����b��?Kz�?�1q٭���-ߢ�l���؁�#���o'�>X� ��	mp�;L�?4���4���xy���?3sB�[v�bT�Z���W�6�(����&�S�= `����\'hp�ꍝ5�ɦ����	�hMx��CM.r�ƕ�|([���u��O��Gi&�v��N�<U͒�B']Ν���麓rb�|�b��	C�3fXJ���FȻ�/�=/�~oS�6!.�y�$�V�B�ܛb���B|�G���������::h�nq��ɍ�E�.h�Qx �H�gF���_�P���� �����V�_��'����MÊ�Z�Ñj�if6'����(r��}]�o眆)��YCRtuw��8(�f�y�S��|t ��p$j?��;3���0���-�]?3�k�����mE7����*�Մ͈V/q��N����86W"�}V$	�R'G�cAc�O��z��Nh<;KL������@,�cWr�T�T�Tc��,�L�e�M3�"���
?l0+հ�яb��A��^���n����I��3xT�Q;��f��'(+�,Z�V��{'�ga]�)�C�q3ha/���5@��Ĺ� #�_WH*���%�ʴ���/ҝ�W��{�2����m��-��g�'e��m�Hhi˥S��HV���*��� ƫ�ռ)㠺�ѕVm��/4�?���i���w��o"&��X�6��:���;�u��TUM� �_��Q�A�f����ƞ�����,Z�0�;����s^����Z�YI�ω�G ���w���-��8�� ;�009gǣ-|�l� 4,���TY%���;`>����_֯�SSJ5�w�U�Iﺗ�Bd�Mj���W�6����
�i���PY#}an�C��w�����g.�3�J��4N�����s�3LŉN�i"�~�+��Z_JX`׀L�KF��ފțn���_�ԠHC\T֙�m���[h��u�E2�����k�p�ٞR�FAT��zm����eK6'�
��x���crY�=�-G�;a�������rM��f᫼��(�l�VC��c����m������HS�Y���Z$�("�� �g�I�g��	��>�([���E�t-	�{��5z����<V��5�pe;�Uj�ֲ�e>o�hG���d�P�S�2�<!��m�cjf��d㳉v�a,����m�V�7O�4�%��'�`�ˬ����=�GX{�""*�NG%U��_�`�����y������L�v����3��(A�H��h5zj�v�3�r
���qZM%�*�WE3��:���[_rbQ\\O>�y�"S�^�K��o^֯���*{X�('\V��X/h<ѯ��_:��,�\�\��)ɳ�lWu��s}X��!u+X������Y�۪���"��l)�U�9��1{1i�R=��A�����j������=�s��)�\�J�]с�aSf-���!Åv$��Ż����pH��l���9Q72�giw���@��ௐ��)W�m���a��^M��D��Mj-�ђr�_���RZdz،F��y�AX�hx��ɥ��%g�T$��V��&wp7�Q���Po����T𑿭�D�,�u�|��B�^�����Y��e�������3Mظ���~ϑ������I��1��O�I-^���������x�����T�� �`��v{c�N�3�!s�EE%��Ġ;��4(9rWרc@��6x��	�P�e�+��/�eշpܕĄ������Ҧ��k���T�L�����Y�|�K�&ұ+9��r4�v������y�~7���N}��F�9Q]T�%Vճt:n'@�2��|ױ�%�IG%䇾�%��ɑUK�c�/V���kC:���)�� A^i�3	i$<�~Is�Uб�x���e_�E�-M��N�AՌ�1 HdG��am��W�)�ɋ\fOON�����i��&�~r��d��A7KC�q��	�����ڴb�h���A!SmZu�I��/�F���Zq!u�� �?C@��u���3��@���U�Ѥ���4��T�vH��7Ζi��-@����&)�4�I[���壅�����S�s說���}��Ec��~Ȋ��̾�p��Y%�����J`���yO�o�e�YY��*(<���f�\�p=�O���XL�α}�L�¸Y=���ߚ$<}��ۺ@�[���;Z ��:D���ة{�%4]���B%)=��={o������0��Yq%-#�[�Sή�|�jv[���G��������h��D��ǰׇ'���P..%���k%����|�f#�_a[�;��q�Q�$fY�����szAӫ+���,�7�H���G��lOU���[[0�h��}Ö�V)�����+.�34�]��,%�e �-3i]�Z����B@�������W�IB�����A�M��S�oQ���:~��?�>�^`!D#��];)�i�]��p z�m������pF��Jm��ͯ�wL���.Ϯ��l��g@ ��"��{�O�����B�q32�ox���-(Yv?EE���q�:�[':��7�mp��6��Wd$U�A�����`����?���T[��s���c�#��K4��z�r�Z.��5��7����_�6�#_}m�SR�����w|5WV���u�N���N��-d����*��������Ǳ�H�`��i/I�Ǹ�4e�J���g����(.��ed(��uW�lM���Z���k�}|��r�+.�̮����5|�QVҾ��eP�rÀ#��Z�S1s�1ҩ���Qb�k-smj@v��M��W~]���[��ҡBM��l=��䀓��oh���?{����߿S�)�L&���W��*��T4'����eϮ�9������>�%�1i�R���6%D��>���z�� ��b����6�w�n�v�+�D�tό�p�=d�2\ɉք�p��+�ތ���*Ţ��Tm�N�K���7���+�߄?���?�ph܎ٚCr����`�c�:���w��$�L�y�Ai��7/1�1Eg��N�b����q*a�W�udZU���W�H.�
S��u�_��{�)�X����I9�Nt��=�0{H����l���r�Hw��i�B�E
zԫe
�;��`M5w�����=/.��/V�f���f޳�o6fAW�~����?��)l������,T��)��ݏ[�����뀐��-l[��\s^�d�ԫ3#��HT��@��,�ꬳO8�H�\���{��S�q�����v���t�8H
��4��ɥs�;� ��z�)�Ք�2l��I���f���U:EF�b�6oI����R����y�Q���e�(-_!�t�?����e��Ⱦ�yY���;s��-�$w�]UJ�U �����p����6@��D��oݺj�ĕ!�&=����I��9B�?�S���|��&>���b�V���Vw�R�@~�`�MH,�)D(�A��O����7\�㛿qh���NR2�L̋Fٞ�Cg��N�������b�Y]�cz�oW"nb֌� �5
�YJW��&&��}Wr��D�2��'�T�ݰ� 3�rЉ�lņFA 	ڊ6 ���N��Q�Vq�J�v�ِz֩fdj{>���9
�az��x��E��?�Y�pC!���W��� �1Jι��^�	L
��F���~�
�-�������X) �@h����ޗ5[�%oi[%��#������6*F`�#��X������j���Jj�O@ҋ�Օ8��f`&dhfA@���푴G���vo�P�	�yU��|�7�j z�4�u1d}g(<������CՉQ�7T��������H���49���i��d�ا��*-u�y��I4�o�������<���%�Pt�ɺ+�4�x�.��&	�$������]@�]��s�J;B�N϶>X�t�QqMT�) k⁢�n��_ɳ�k��?G����N���<x�YZ��� b�RĒ����K���2M|�֓�*��G��yV��K�5�R�3��K	kn`:�Nȡm���~���Q.��9�3(hv��7��8|f#�Q,>�/f�[l��2�� ��'j�ڡ)���(&6_tG��E�q�,+�&|�����.�iP��T¡�t�!�e�	GM���B;9?�*��^�D]�f�9��]^�-H�8��L�~��5oq��N�e���Ȃ,�5�I��E�9\O6��M�b�`���3&,B�l�f���֢��6�h�Α`�	�Ȯ�b��H��sNv�+zEq°�}�/��k�5?���X���5�ڶ�֓��Z�O�Av��鬍��� RP�l�b���|[�mL(.�F���\r`{d\,�<��v��ߪ��(�Vz��u
��T��ѹL,��9#UD�ҙG��8���Fz�x��"��>ϊ|e>ӏu�o�A�ꦘ3U�' ��m)r89Ŷ�-'Ǳ��t��h"�F����>�px\NE9��q��N]}�c�E=���3�T� �@�sD����=��	Fv�X>'I(�%�Ėa�S��
�_5#lT���DHFR��a�÷����D�|s�o��Q@�w�{�����ww��<ྂg��%���.�*�,{! �M� ���K"�J8&��װ��+�/k)���-/�`q��G@��,�LB�4�}{D(�cY�i"?�GF{蟤�����ԑ[8���(����k?�p����[�	4����%]�܇X;J���I��Ze�|S������cnj���T�Z:�i���L4�l�划��k(�NH��������r�u�0$6�Q�?��~F �G~��_�xG(�Kf�q��Rɺq�2�:z�ԏ��!$�&�}Vw;���1��1ngA� 5����_ּ�K����� E/�Z���O�f[�9��M,�����3�W��w�n\�D�ݵ��`h7�
���<PQ��s���NT��<`Ec�0ГxH���L�o�v+���B�mcyW/[�Un|��@��:19�P����o5��� ��~���[�9��T"�lj�P.M�� �*/v�y�2
z��~�j+���-(r��}bTj����a�A�>��0"�U��ˬ�d���(��m[�,�0�Q�j�nI?D�bQ%[�1�"|��FsH�i$~���Tp�
��ؑ|(:Z�R�*�8Fc�g	�����a�gSV$�?�l�'4XeN&9o	��I=�Զ(���P;�K��߷Ã]�d�􏨃�8����6���.��bB�؏��q�V�=����K,�t��������E��`X�z��*A�m���EC3��ԛ���Ӂ�>����*2�g>ݳ����g^DN��u��9�����uS8��ŤX��b�AA��I�y�܁گ���c�+/pr�~-�H���}��_�Ҷj7f���O�H/���Up5s>�{<�\� �?��S� ���0�*1��r�#ҟjj���F�O��uQ���BuO��\���������~�hyɹ���� Z"��X{ux�ι�OJRF�0Y0����e�U�c�)

J|'I���@'0g��,�4<� n[���MV5�Ũ���\�oܹ,�"�1�s��h�[��Z`n	�w���G�N�iO%}�ۍd@Cڷo���ǾQ�"Lŗ�Uc���@lw��h-8�w�P,���x���>T��r�
�!_�uAZ.���@ڌ|$m�ϲ�]�����Rۢ���M+��r���x�&c��8*�]���va]An��m%w!�Xҡ�fL۲CHʭ����G� Sm��[���u�K�V�o��x�r[��UjN8~.���w$Zߧ2VC�G��,=K�4\����j_�J�[!�"\�"fb�g�(�4d*�^��t� Eds?'�A=��hKv��9Ʈ�a�����[R�]l���}A��?_����j���,Щ�z�AyS��|�뗌#E&R��o�*?�[
���q�A�r��S�qm+t��`�J��6F='�}�g��k�Ի��^�'�m1�x9�Y���V�����>%u��V���4dU� �nC>b�^���6�#w����[�4V�{���Ŏ���׃gߌ^QR)��� |"S~�eO�0���hXަ$
_�x�7߷���
��g莚̡;�(X���w-�rNבr���E`��Ѯ. _��F������r;Kvyr��(0��X!�_(ą�,E��T�p����p�/�vө����U��ߥ��aY��\��O>e�l��d@��x �)�M�D>���mS�|����Nä�'�J��/Kv�$��<�qf[D\�'"�T hv��ɓ�<lCJ�Ǌ�G�Gc���&܂�(O�<.���Cr�'���.#NXL����B�S��7������{	#�e�VdU=(8����������w'&ε�ۃr؃�Ŝƀ���G��*}�kO;�&�|��a�Ia�N-�}�O	��hE���>h�W��L*��B�T�r�9��zD�4&8ȁ�l���Kv��G`W�q�C5Us�+Cc��1�N�iv�+,��5�9��\Q�PN��z�D7�zq�JkH^( ���A��KC��w�E^=cM�./"�6��M�K͢���p�-��l��y�.��@j�!��A���OoB�BV���uIp#Mwa/v��C���r�[v]����pu�2��>w��F�E���f�<������3�V1�\vZ��;�n�Ĥ}>v;���+�ݫ�6���&[��Z*�3<�.�P�qS�y3c��)���p%ا�����b����V��̀��V��&ܮ�9{0��@ԋN}��]|�Z���S�! ۿ�\��<���Ia�:�bG�yBǳ�ps��^tUB���G�ͪ�EoK���?N
�D�8`B��G`'����z�u^��M���r��Ō-��ń�ӡ���*���B�^������"2<J8����Ϋ����NEy����T�ǾW�A89;SV���Jt�D�,A	X����jbg��yE\rΏ����E뻈h+���E�o��0|	ފG\�é?�yQA|\�Rr��'@����oj��>�F�I�NȜ�_�s{��2ĩЏ�f0;X���W	���[C&����ܐ��|�M(ֹ���a%��K2�Є�=鼱�;GQpio����r�@#�_��[�p�J�`&�&i��Dp@5jj��R�'b$��Y���������`"�z����y�Ct����������� VH"D�ۭ)HQ옠�U�"������.����N(�C[��G�\��EO]k�=�̚h�/c6����<�J7�������D%��mc<�g�X�;Ƥ	~E��1���h�_z4�x��ߔ_U��Q7�T06�}B�����2-����?W�1�9����������<e�s�d�x�J���FS�H�d�.�:"�;SjQ<'���:-:��r8v%o'�t��,7�D:,��"�]�8��ּ� y��+�ͰSs����qJ	؇�x��B�3>���?�<�],`i��v�|����l��W��8s�`����5��2=nw�bq��b��H��Y*q퐒�I����=j3U鶁��2�A��oG O�?sm�S-�B�[�E�%�VC���N�5K�<�����ZX��cJ�_q��lrQ�@���9L��������v�Eq�Ԙ��K�T�rN�w��)����q����Ԅ��Km1���L���W8���]�}Rx��������Q["gw��~h^O���0fu�ȧ�ɔ����C�-܅ɞ�j���S��A��|��y�7ή��qW�I'�-B����Cg^b�ڿ^=���>��)`S-��A��^:�Z#`��P��Gb|��iA@?Idm�#�v/��<_j��a�QHm:�}��6O3�]Qi�*���(Cw����4<W���7���ڹ>�3�d���m]r�w��<�R��]_�sí��n����#��5� � WKǏ���Yڰh&�AH��rOZ#�f����yzӎ�Q�w��'����ƻ$�L���n����6��uc�ΰ����惹��;V2����G�E�U�����X���W������?���I�z%BN8��J
ٹ��fwFϵ7��z�*:��JN��BjP�)v�������p���~������A�zA�z�9�Ǒ<�]�z�. [��QRH�3Za�c��:%�����S�����	V*��@ba���sI5l���L����+��66J�áI$V�TZ���o�j�٣��xT�%�GS�-�*�D�#�i����c�ؾ����u�c|���̌u1�n���3R�*K�Yqtv7_���SG��}��+�M/*��v�����f�� r������(O$����
��}��v���d���u֔:7Ԅz&�~�|'� d<�+�9b=G�<��|4s=>�5��%��e�EC�����i8Ph5 ����|?ҵ�հ���h�^���ü*�EL��q�qhy�ܚY�:�}�wc��X��3D>�w�w�[�+�(�z�}�L/P\��/��0�}�D��Au�a{LBt(��V%�s���Qt�6�at��e{+��c�(��}j[n���X�hA4'cv�t�RC��s��s���f��m-Rb�#��`/,�т�sċ
��t,Y�8���K��M��KH$��8��6�)q>\]Ÿ�����\ :E�L+k4H8>�H�6�(զ��֚a8]oT���g ��z;E�z�/%;�^�`��Ŝ�-��*���
���4�&SX �W�_ۄAi���b�J��.E�N�0�ɶ=S�n�֨� �w�/�p|`�AZ�6D��%ܷ�R�����G��B
�!�+Ń�*~} }t��Mh�N!p��)��� ���^��x��Ψ@T��n	��Z�s����Y��)���8Y�	���.(�A�W2�G����/�YZ����^���s s�C0��� <���~.��n��z4|)��K��u����ʘ�	X��{�;�|<�ձź�ϕ��	�"�9skJC�>!ִ���z��E�R���\����SsX�0� ��K�����糊�D���(˯ϲ�������7a�L�BPj��g�~ 57(d>Q;X��i�7����m�\����n���q\W�1�����I�����FYm'��x�F��j�LHC۩�h�%�^X�{d3���_^U�?6	6�ji��!���<��$�*v`�Ңv��>Ń�J�[��<��p�پ����qk�Q]&<����!�����-���~�tO c���T���^p�_t=�m��(~����AR��#�l��<�U�%��2�03��ZQ�A` Uz���c�CP[���B(�$�d%��Tz��C��$.�(��#T��g���f���a�^xz����S��x�Q�e�+=t����l����L*�S��� ]�e۸����8<F#{����(�
 �H���
�����������H/[/
��H���	�=��Ɨ%��-奒��ߣ�����i8�3�cwz��(+qrG�U>��~��T��D�?A!��y�bun�3 ��tb����e��m����u�$O��N��藈Q���Mm�a���g�L�OA�����*'.��鮡
gLQ��;QO������
��Xu&;TJ�[f�j�	2 zo�C�i����J�!5�"���=�n�d���9���/�-~�W�44�e����G�/�� `�=�U��s �ë��vB���|S��2 ��ݢ�߭��9�FGX�	�b�J�Jy/T��pK�.9C����BqZ�VC5m&p�$CFϝ��sG���2�c�(0�,�B����W)�;"M��%g�"9~ד���ɿ�ήҳ�&S�2�~Fe��tH#t$��L���?�yS��8!��~uto�z�A2�э&Í���fQd6,��/g֏m�Zۏ�H�gW�J'Z���ǡzZt�V/�޶3��4B�K_�&˯�.s?����S�ac�`I��s��	P�o��s�J݆���xrmiB���*����T��x�5b�Z.�0�ɒ]�=�8�e�ѩ߿���q��sK j]\J�k����G�����]R������ߒ��5��³~����	^ڬ]�M3]�<�qٟ�E ���9��Dk�ݤ_�\0,z�843/��Nv�J��](	�Tp6���b���D���lwO��oc�87ԭ�ϒ?Q��\� �����f�\�˱S��ik�A���)�_�J岁�&֥�o��jxMv��	�]�(5�}ܹP6c����	3H�d�N�^�~��'�٧��P�<�#,w �k��]�`vJ�z�- G����ݜp�vI' m�Y� C������̉�me\�:�90�@*{Z3���;�M�X(0p7�f�����x�����	�M�R&г���~ļ�I?K�Q{�8{����JХ��W��&.r�ꅀ��:�)]�&�SP���P��S�?��j}�bm�Z��e�4�H=�!��:��K^�Xk��s0���l_�w�V'�3؉��9�|������,?V����rMkrNo)�{ �	)<yFA��n�& lx���Ң��+��{���j�|c��$�f�m��+F.�8*�3��7�E����6.�����s�*[�F�Q��x��w��J��Y��ϵk�i���?s���(�\�{$��Q�"S���]���<�b�CM>���fњ����Z.� �ݮw�T�N���s��`Cˢc+~.�qm��A�D�m���\�֫"��6_]g�:�D$�E���c��ft�8��Rݙ"��=.��i��K�!�_کь0[���Ak@nF����hI�ѧ����70�!���m(ձQy�8���e2~����,reuf\'�lΪ>s{˛��M�
��HN�&X�EzZ٥�ႍI�N��8ch�yo\A�ieyzƿ'K�&?��V��F�����WQ���8�r:��`u1ӄ����SG��Xt9D�]��[ɕtD$�rYG
�	?��[#	���ˊ|�'%��)Fܥ�>]�hh��]!% <�D���*�R��I�80h*��87[�D~VŠ2w�����a��S���eE�T0��6V��r�=��X"}.��3�E@�v�$	��K��cܣC���@gT��N�vN�誻Dȕ�BBcuMM7u�1se4tY�ԩ:
�V2l��&�\��d�.��/�!xǶI<v#)$��Vh6�b�(�6�m��E�����p���,tQ�1�][�k�Ï��-<���D�,B���,��g��/�&�;M`��eo�ٱ3�E?e>~�P�#���<��f]��Ak#V+��h\5IB�8��@���� `h-�dL���K�������%��c�b'�QҚ����X�{���c�Ņ6ʉ\�x����UR���L�#�H�L2i^��{���>"��� qѻ��t)�>��fD�?J%�ÌiN\pnz��ҝ���qNV ����T���;4]�=p̝�q�-P�^zO��2��}�Qp�=��}�<*�o_�(ʦ%�"��)�ߎ�w5����Q�v�^�P��:�R5�@Q���d�_�V�j�2�Q\��bi��;D�g��(f�"�������a8T�՝J�Cvm�7���ر��"/WxW�y��2�T�R���ѕD{i�ڂ\�-ڽ���qš0M�LNW8x�}S��a��t�EM˨��*b_�z(�}Rq����?�,Km����bٟ����X�ހ�_����
��� �MS9& ��և%(���\����W�n�o�sє����7�V��)�}a4)u8��H�<-P�&�)��9��E�02"Z�S��/P�i ��|�=<��d�ő�
�X��m�9;�=�6�
#��#Cb�3΄��/�oZ�i���?[L�MO�U��N��-��n���*w�	�s��y �q�D�� ����
��v�S<�R�#�+`Z�@çϵ�ܣB�
g��jLϥ)`�^��#�=�?zT�Mmڭ��"0U�(#ܲ(Y:�G��jpu�4��jf��N)�}�{T�l�r3������Ao�ԃ��
�Z ����п���t���ԉ�f<��'�ޭՖ �k�1"�
m
M�nxahxi�K
��j?�&:x���W��|j�JJQs��y�W� �"���a����\���
�_A�����R��]I�F#��_)L��r2�%�ko�;1�-1��;uP��ﹻ���q��N��Q!�Gv�x#�[�vp���w%
r��<*%�m��i��l�~�AT� .�Y]o��<\����Θ(�*׼�n"[x�mnKb�u"���x6E���'��r��߾
Z���8���݃@&Be���teN�O_�������,a�>`�,��S^2�U�'���Y����朻�O�y��w$1��`--�f���4[_|�ٛ�W9�y�`�L���YxM?�@����=<~5j�F�h1w�p������d�gi����~�F���f���(����CX��f��l)���(�@*ų[�O��,p�Y��1����=��7>�J�{��c�&"J�A]��.>D�-�U{����8�:Y�ƿn�=/���: n�|5��=����b)�|��(��=�����\ؑ�x�4��{bAm�:��7��M#n��Xw��x�(c9HW�4����j�X3;���t����AO\3R�l.�i�p�hh��i��i��UH[U�m�.���%t�VP�&�rpH|JBN �c�m��&�àW "���_�c���zn��J�+J��\�;H�9�Ж��Uܠ�	H��Pq3]��.w�y0���]+�|� =SX���R0%7,o����N}�؏��F�7K�ȸ%�D�1��F��>:�0z��i{��X�����G9��������\��;^-�+*hQ��_�Z�_/[�ĳ��
��&v7|,�'��m��.h��S����Ii+�CG)<X3�����k=�<@��N�)}8�Fڍ�VI4P1�l/!��J�eO�i��>F
t�h�" �^��Ч��n��M`��0�D:��<NA� ^g���8��;õ05����Ro�-�7�9��6H�&��v, ���$5H�g±Vq�H�08_0A2�*�O�x��������5���X�2_�iܨ�
Kd"�v�8'�*vmꚸD�v�ɈS���5ڊ0��/�%1��Ӟ[�TA"�P�Mw-�o�.U}��K�3��:��I��JI</P�� ��hK�̙7*j�Ue0�]E�X�(��n���Uv��6���7n&���IG`hV���A8
ʘ�P�R�>����f����=d���V�:�7�a��"�����I�PO�tp�D��=��T/�40��돸�`3�w���&��	�ɵ��|�[�ݰ�*�1cl����}�����lЛ��$���OT�"3~����;z�qA�o����+��gp,e�+it���&^��FBQ@'	�,����HGh����#�ٌ�c]�D�!ɥ&}�|�&+5.b�ߞ�C�I�*q�����좋mrvBkY�{o��:�����˺6	i����U&�G��C�\F�Y%h���ծ��4Ζ���	u�ѝً�k��������jR����,���BaS��br�&ٳP��� C����i���BJK�ܵ��΅�lC�ZW`.��@7���1�����@u���,F���V��֜�Fu����b��N)���t�W�[7v��7� ��j��~t["jP6i�#M�EB�<R�'
|i����m���>�[b��B}��j�ˡ���첒�:R�����O�W�lEkv}^��+o��t���zY�kO)c",����Y��|)�d R��C>�$�Eӈ���q��fpS�[�B�&��$��M��0ɞ�͚{ږ�A�m4=��s3�\:�L�\C��J��^
��ir��������g�@,�/��^���(� v:��a'e@�\�f//&U���v�Ŧ��6R������c���U3�3��Ļ�F�����Tfv��M���Q�ZD�áZ�l�CH�|1�E+�~�S�c��a�M`4!��͘���͈o���+�i��ֺ�dN��KnPT�?��G
�Y��N�b��L��;�C�d���~��v �⺲�Vؗ��T�m�q�f������8lΝ,��X�X!R���\���\�.R�>��ñ����%$3��E�����{ٱ�?�}�H�v��I��O��q��Ы�	q�/��R�<�'kG؃�X��9g	�#���ǥ���_e�"���!�	���V��΋٦v��	��ʍ����|�>B�VV�����K�T�3�d�PYZxXk�x�Lk���)ǎb\�0m���
���g=�OI鎤�Y�Q*�;AA �Ǟ���f�������qh��	����ݪTuN���gH5�H�O-z�g��eSU����o�Ҟ+�|=P�3�R&��K'�J������G�S@�FV�sA}J�}�ƃ�6�����u���D��]�!6}�Q&:s���c�{?.C������?M�k$�җ���r�|ZS�4]F�ΛG��Ȇ��QV���idm�>��Z�AxK�h�:�*p�"�� OӜxt�ZpIp2|�\��d�͠��v�cb>m.6R�����g��&)>Nb�|���$�5,��:)��Z����W�C�Ђ�i��)�
i Ģ�v���erm�غ"���D�D�v滋�=$'�W:ӗI�F#�]3�W;'zުץ���B�� ^�ػ�)FΌ��^Zw����Q;3��+��dH^Ƹ��&����ٻ�R�@�J;�Ĥ��Ӕy*����)H�A[��u�>!��'������{� K�rP�,�nvr��s��k'U�	�>ݞ�Z-�t���:��Z�q���Ķ��L�o�]��]/z�f�F�X4i��k�xH��DPU
�=DS�ـ�.�����Q��s�g�٭���ַ<BkL�ӻ�#��#`XJ7 '7��:AVo��'��?Hpcw��T�R~�`<��
ݼ�NT�R��/�{�lYe&$���O��HЭ�^��ܯX��+CZ�$8D��H��@v�u�2��Dʋ]ru���Vv��q�)\��?�r��Rhc�R-��s�L�y)��(����Ԍ�dg�jƓ ;f�h����r�g���J�|�)lJ��$�ڕ��@v\��V�֓�KDqB7W��6�R��C�Z�i�L�o�N����,RJ�G���6�5?�k[�A*�~�U��d���Vtg�����!~��C��?��E{�{�L�Wn#�Cxe���tߞ?�o�B��B�X4V+�y���R;�u���.�Ν����&�s1Ů,"���.gͣ�j���`kJ*��l\dG�{3����y�׻GQ�u�1�yU�*��ǲU�o�"�R��O����]Ѧ��\�D�<�ŀ$��rUE�ZA�'fj8ABP*�����?�x�5��wa_{�5��5Zs�Y�l����H_�����{p��?$���5����� x4��<�$h����uG��{oe�@�z��A��jޮ�m�����x����h)1u��XTލ̘4N� %��o�khҔ�T�4+�W\�j�a�N�hևˁ�{?{���}��h��?��N��-�f'*{�D�N��t���,�ɣh^>D�1��I�]�B!)V>�ԙ|h�dh��~��?Cq��_>����%�Y �B=�Q�0괳:������^�۫��7������