��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��S??Gl��i�vDM1�<����A��^��j���E�&��Y;�e�m�8�SY"p:�P��.VJ�4���} +x5Hߋ�άN�y׳#ן���i������] 	��@�%���gG��t<C�G��F�N����w��S1�'�)a��Ӊ��`"�Dn�wݼ>�b���E��9��RV��<�+����r`� ��%d�x�M�?�I����YÜ+��^���t��Ņ��;{�ނ��x���{�����F�%)�Aŭ�8�t��_�k���r8B �����͆��ɦL����.~��Q	�uȞv�*i���ϙG�C�-�㈑�U��Zk�y(�F��ݟM��B`�R�1�*lʛ�L�ʘT���Ѥ�u�RQ�$�I����&4u0Tyy�U����w�${FO�'�P�?�ŉ���#��?x��8�۬���������Z����iL�Ҋ	��Re�>�%c$A�`���]��b7����X	ٝ�~�q���w���!���;0�~󜆟�Tj5�$��StZ�%����Z0�3�I�}y�23�@NHzZ�"2l*�͔h�Zu��3���hJ�e6�'W����Mq��� ���^����x�w�|\J��[A���=7Oc��Ae7��6�a)	�:Nͫ>~[��j�T����X��=�����C�;ؔ��y����u�蛏a�j
WgNX��"x��F�����x���d���3�'E)��d�Ւ�>��at,��s��=��-�X�����m�!Hh��i!_��W5 �#n@?�^�̣>m,��
KI�h���̒�Z_]�ɮn�bޚi�S."���b��)���	��
+�]�z��3�8�H/1���+By��s6�`��#�-�t���y�q�L�I[Wz�P՚�g��i�|�!��K˽G��Z�Fа�Y{;3��}�i���?`�a���9��bx>W��}���
3E�\|���!�W�)/��l��/wuxYP �z�]�@(�mwsv�"���*hS�h=Ňge'��4&?�ܨǏ	u�0/8E���G��>O�
��b�]xD V��	�PP/��&���]�_��1�3�gB7����{КZ�-�@�������n�>��J�e�#��v)c��N7�OY� c��Ê�V�,�/����y?��!?�7pt#i�'P�A��MX;���M�l��E���W`���m�}�� Ӱ|E%b.-�)Ɖ>�v�����:��6j�:�%i�E:]~չkC��1�׺�[A��%�A�R�2UG�6�~�쁪7$��zA��t��9y�D�F�j�������V�;=�2 �Ji�f�:�z��oNI�ռ�`��BUh��UZT���#�!*���`�2 5�.+y�����Q���9"�ħ�&�T�͊�$�7��FQblmk~V�"us.u��̙rn��x3 P�[��Xc��H9���Zv`�@�̊|`�l�ǝ?"��}�Z��IS�)�{X)��ܪ �~ZZ"��y�?��W/�`'rR�e~�`\��� �Q�`�x9-�]���� E󎢨����z+�ԃ�J��,��UD�bL�& V�rg����6�Jzdh�nE��6�	Q9=�Ј�u�uj�b&�&�������;i.�\AQ�Ii>(�� +�L�/��z�b·.�@������0�{"�J�xr��=�DV���dų�{L1]:o9�ϻu1�X��<�L�4>�`�/�+κG�y��I 0��D�����FXDO" t C�ӎM"�g,�G�_���\�Շ[�v,��"�%y���H�Z��W�J�1��k<���<�Ĕ�u��cU���v�[�9���j�-x¨��t��g#5:�u�đ��$/Q�7s=iNA�(�L%�Z]E�ۥ�3���_v>l{�R\}�ؕ�#ƀ���}����f�x��3P�/��B�@�B���`{�fP�p��Fs!���HDI�'�E��҇��B��0Dڕ4�&`|����u܌�����y@��(�ݒ����P"Qo�� ��H�W�)B�w,��#��2�'G���xgCu���&͛_��a[���~b4�f�ò���������Ҷ��:�� �QQ02�l�s����n ��;2�wEŘ��=j�<�+����CH�b�r�a��'�U֣8 n]�+d���wME�	���Ke� O�H�O�b�߽�ͤ�P'[ ��O��x���V��!�.P��J|��<����e��O?,��e�/I//�O�0Z;&7�j�D�W��v'��t�p	`�F; m�eҡlc��4��>r�'�v3|�OA�f�!�峌9*$���jԽ�!�N�+�x#h��L�\����l��a�N�+C��M��/9��D!b],xP�ƕ���i�hQ�c�s�Α��-�th�w����
�ԴE������h�<������5�|ar�W��ő��N*eH7j?�ă
�X��zy�m?g|�'��+499h�^��u�L�J@���I5ʴ��OZ���`Α&cr�Fp����<�G������>�7�Lv�r�%���ì�Y����	X�R,������F,����j�}�a@,��2qB^u[n����'��-�}FFؽ{<�_�� ď�*6].��i����P�ܬj���(��d|��j�_��j �X2�PW+e�%`��Ǒą"�ܪ�����ynfg
���T�S�a��E3ŨL��P9���u��:v8�8���4��m�_E)*��رE@@��LY��r���_̿�E��kn�M��C�S�	�H�1+S/��<#ꂻ!6��D���B��{�7�M�-�z�"G]����}�1_<ȯ,Rg��]3�$�4@j��m�G/h#�ʼ�����N�7��{� M�d���_'���1@��͠�j��~�N�0a�)"��b����df�� �NDiʹ�h��vV,y�׼�Q{*lw�x	"����z)POt�㑩��S3@QR���N�5��F�Xc�T��&�o�����_7���#X���3�\T	 s<.����������/S*��_�98������X��v@�y����@�a���:����TJ���U����y�M-�e�������s+(b���%o?cVg�
8zY����s-�jy���pԢO|�;�gX��-޹U$8�5-I�{�M?h��`�yr����Ӝ,��w`���C(���&�s��/5�������s�^+�x�u�B�	,m�O:O|��7�gޜT��:����=�1<ź����TH���{P̜��a� �����Ѯ�'�����f�P��{mļ������z���)|��=���P��u��wz�U1�l1:tK��NR�]M����,F�'�%�n�]<�R+��E) V��~y'֐S�bW.��/g<���8�'b�01$O�U�#�n��L�+xF^��p��%�QR�}�j�;�(�7�����"�ġ��<?)G���h��~ͻ����=�~���60I�3�Ř|���'P��H'µzV6��lgE�)�
�[F"� �h�rwA���7}��᯦ny�OFʩ�Ϗk(AjƼ&0�M*�_�!%�p@T�mJbs����vW�A��z��!g�h��j,�p7[Ga��VD�9g�}�4�V��6+=d~Ɨ~-�T��8i:h04�D��Q�:�c�墩�`��i���!��Q����~�n���~�����1�1�1�<��!������:�/<N�i�lMS20h�r���^f�$�/D=e'�R�;hb8A����X<����+��~3	�R �����	��c}�Fׄ���t�.E/��lvj�69�|@�):�AhR9%������a{8Fp�n�@<�w�i�U���?9�C�,^�չtӗ�vG$�J�^'L���v~���Z^T�H�NL4���l1sW�l�G ��|M��q��9��V�:В����%lp��m���G�;�d��IBQ9�����<G��}|�l�6��M��ṔE����<����hPi�Jl_ذY�jZ��+��e�̅۴ F"(;�<��K�\guO�f?哝Y���F�8V]�ge<E�Q;�ү�!�4v�f���i���R�O�Ζ�b���Y�*_�G�j���D�5���t D�B��ͪF�]fi����K�F��@;�K���XL���F��#B��p�߀��m2�лn^��y'��1�HS����MOI�1��!�y.d~�dO�%�=��W�� ���=�,o�:<��5��H rۑ�qn[����r�D� ���%�젇L�A.��������Bx,9�_���Q�-V�������z&l$!���U�|�1��P����c����%AH_7�$m�q�!���(��D�4���r�
���$��uIr�KP8��K~ԋ.K�!��Gc��A�"�NG*p��yLc|��Ca�C��=�����y}���fƆ�*��WQ{QwǷ"ݼf�.`��T��Ϟ%V�	�������\�R_�s���L��,�J��,��ӊ��o6f�WY�YD�
�����йZ��oĉ�V�@e�o�\BK�`�J�hawisQ��࿏!�T W�wv0;�gCU�3�U�%��U.B����X��M�R��d��E,��$=��J��Y9�p�$���'%X�`�O���J�4��(���na"�;<��ʀ���Kc��vǹ����l�lt}�}F#Yjva���v,�5ˆ4L	�����6n��z%Y�v�}����3�.B�ޭ�l�N�Զ�[8����6-��� �ם+���sIiJL9]�ֱ����_7��/4	J��f���i�<��7��l��)$���c(vz�"��\��� 0S��8l�F�`�D��俴�Nw�"�L6|a������p�>���`^҂�|]�b�����Ѐ.=٫�F���[����(/�7W�.K���/+��=-7�~��M��ּp�9;{m�g���
=;2�bϤRg��GAF�������a��qLyu��.����%����F��$��fX/�,u{�&^dC�j�����Y��W%�e[�G�@������ kc���4��Z���\�4/�N}����ưI��1Q/bX�*QoX�X���!^X�1R��)�e��ʓ�L6���λ��?�p��`mv��H����Q��֮�Wc��i�hM1�ѶW�����-L�Zy+�2^�1��N�E�6/{����"���`B_��K=��CKM�h��2W]�\�D-w����m�2�ˇ��k1�����l~8���7@��q����_�\�C��|d�����f�7�I��c�h�,���j	�*��b{�Dj��׼������0��G-̭�􈮩��A3���K�kl� c�K��%����+�.O_�z�R�֤���	���mc��xъ�7<ܫq13��g�6aD'bA���e^;dkr"������9g%V�U0�V{�9[�B$I�Q�Jr��&܆�|���.�%|��� �b�ɔWq x�ӱ,`oV��I(�p�q6S~L��0en��	�|b��Oa�h����@�I�NY�,�߫Y}�Y(�֋`�_�	�LC��=��W���:s�S�_\��>����! �7�f'b�>�����=Fx�-�Z/����p)H��Ͽk�^�-O|/�1�{��*~�*����-Z��~F�������,�������)�S��Q��bإA�o�j͞s̿��^��m �e�q��V��c9�Ui�|��JU��ǳ���^�(Kv�	"IK}l�5aB����P��f-L�v	w�jƷz�`��@9_�5=�^����gB6�)JU��	��E�ϩ���)���B��wU���XY��Y*p��~��B�ș�o�=���oӹFθs�#��_�\���.�y����8��dm��"%�]��4�� ��^�XmW%�ȬRO�VC��������D	=4����|��>ȏv����W3���M������� +�\D$8U��8���m�"��H�T���|���?1I��(�@��{���A�YDM�+�k�I��
Ռ �˱�j�0�x�=��D�a׳��l	�1��C[{:B2�'TM��QlE�
0��{�3�$�A#I��	��9����x�1�1�[	v��|�IS���ű�'�$H+���:����Z4��*GK��H�*b���lV�)>�h�����U��7�fm�fS�# p-�H������jľON�#����)�yt��ʶ��ˇ�'���ie�J,��x�<��U<��������>�W���ip������N����#$8M�M�o̻���d�4�^�V�q�k��jDV��kW}�ّ�1��. ��ֵ�7t��%�����% �s��kCq��`�>�f�ZHJ�dv�b�!�*{,.&?�u��w�\�����������/�Ti�Ep����E��P�M��]�N��֭_	�.JAF�5�@\|ҭ 3Tk��gqh��s-�Ъ^�9�*�B��m����z*�3�ǒ�K)����s'�=gEo�ټe�w���i�ܥ0U��A�����p��>3��F�4���m�NN��?����5l�h$!��YkqCܐ�r֏���ϡ��II0ˎ����Y�]�I��4v\�p:�!���)������4�^�Doh7��Qٿ��)1��XI0W�m#+yF�T�9��<c4G�,�ALӇ�u�{ZW5��rµ�IeN���cna�O������e<׊�cT��lzYT��Kz���E��F��P�;���x�Ҟ�M��K��a���H�QS�Mr6c��m�1��JZO���b{�Rĳ��{{_/#��*W�h���TY�� 9M�!�F|@d���s](b|�3#�g17����J�\�S��\���#����E�BX0��Q��d�y��1N�$��1�XTv�Zx:�~����t�����E��|zu-4ӄ�M��|4��L� '����A[��<�}H����� �,��%��p�
�h�,+Sd��do�)՛�K��GQb<^����\���Z}��� ~4�.�l9L�0����N��rD9��P+N�r�ltj���6̮#k�Z�0Q�M�fŚ�����J���Y�f�G�Jgߚ-��L�{�z��5��I�2E������,��׹�kyj����H��R$L˥��$ìK/�ΐ�Udb��+kW���V�׆�Ì��/4$2���4)U*1E�f8�rKA��wܒ�X<qx�<dBy�2Y��!��;���o[�^J1����U��tx�'2��H�$�x����y/��hzhn�?} y*Qk�A��T��چnz�Q�^0�6g+���{K_�q]b���<�)ۓ�DR���}��*�^����<�q��=Q&�|*�o�xh���Xj�n6��]j�le�*�N
���?&H�����M'_J���0�;v�A���"7���(ʒ���X������;�E���2l�m~=#R`��|�&�3Wy�T�����l��
��<���mjc�T�"Zp��WD�CGH`&�3�p�ʖ��Ȗ��뇀����N��P��@zeD�{zU�N��k0��R��Z�Ғ,ެ��u�&���S\ռ7�춊7���=�?:�����!�Р��=�Կ��P��sA��% U�Jbg��7��ϳY! ��W]���v�>��m7��� ѹ��W��=ߢ����3����!?
��	Y���US7��H����Ƈ�pɵ���w�������"6*n�В�o\��^w�ڡ�~�����;��R� 'F��i�ãǖ��%�q��7P���Љa��E��m��Ȥ���] V#�1|�؛K�~���׸�O�Kє5��rcU������
�n������ ġ)"���\�개�=gNN����MvZ!1�n���%�h020bQX�WkH�ό�`n~-�Y�Bm.�B;��_ 	��-u"�)�@�󝅤6E�t��w��U��������S���Օ5C��-WZ*6�*ڧrKW� G��F�Έ	Ѱ�����;x�>aI��7�6_E�*9��� 2���҃`���Yb��b��]샺�=�B�6�ʊ��t^W�x��Jo����Yk՗�(�ݎ]�h�!�ig����i�ʋ��v����8�1�a�>p�n�4ݩ�򮲄Akl�B���8V���q�B/CZ�	��삉��O.s�����'�cH4r�sw}�@�_J
\z��}�sHDͧ�iD��K��}2e���ߚ�	|���1�L�{PJρ�̄���be��!6A�
ř����(�K�۾�\��J[��R,�đk��l<.�)CHB�6'~U����R�7fAv	�����P��?Goş��~��z����Tf�yb�m����Ɩ8�G��~	đo�l^�Z�km����m7����,�Zͥe�B���0 ȅ'��;��lCגg~|6^�ђ�������+Ll������i�֑�N<�F