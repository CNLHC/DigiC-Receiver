��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ�����cY�r��j"#�ݻ�|�\_��Ü|N��c�H�4 z!��܌Y���O
�nV����諛�]+aaG�MT�x���A�C`7Ƴ�nϤ�� H�XT�m��%v��e��b�F;��n-3��r�ȧq�.�m�]W)�I��t��,�i�da4-��v�3u:ܦn�,�dk�<�53�^��!}��mR��4� ��uYVɪ
ײ�|\��Qn�� �������M��]�p�Z,꼯�lGV��Pu����2���ފ��^rL�N��dܺYHq���g�3�;�^�i������(7<�I-�ӿN8�����Y>���r�)�=�Z{���T7�:!��؆V��BL��͍�;��*����#��"I1����!U�VSrڧ?�0$���L���$��đ�[����������z�3��:����ۏbQ	ҵ��=q��IN�����E�Ҵ�&='�{���Xv�K1���mf=�RѝP��:+��T@!��i๬�k�B~��������_Hb�t�Ѐ�(�:�ڥ�d6E�s�=��.��	[�y�w�ć�K .�j�Т*�:�Q���31��!���33c��ı�=Bi@��K����[�)����k�R�h)��d���i�
���aO���6G`�Șet8$��B5�#�>��*�C�9�(4!/o�c{���C�
��Q�.��������������.�*���&Y~E����!(��@�J7��6¾��^��uJ@>Y�~����ů�ygaf��RA:#��K���o�R5�	��޸�ꕥݫU�6�L7x�.S�&�ډ���B.���`������T{���FâD�������ow�= �lKxUU�g��E�v~�"��
�} ���#�'uN�u���2lЯ��*��cG���$�d�ƃ���dҷ\VV��9�?>�K+��7��4���U=�1��B���xZ�̱�=�i*LA����{`���+�#����T�c�&���+CT���� �����{&-&6�����AY�r��~�p�/�nw��1��j�/)�c��ӕ�X��yz���A��uJd�Q٩��R�,v^��Y�X�d���Ш2���Cf�T����A��/����ߑ�1�����j���Y6��� v�O�_nX3?"tL��bǂ���4/O���� ��}t�SQ�Q��@A��3�E�����[Ql�����#�<�e*�n��6;��*7��z�K:��e��}b��=��V����5��2���@��\=�!|I���>���A ͪ��W��X������9��������V�)2R��!80:�y/�m�fj�	%�p���3Z
����!�^7�)d�v��7���0Uuc8�Ln�^d�W��-��6��펼i���;�B^S ����[����V�ۉ�{��!��)�B_��tRY1���Ɩ��6���j�ɏ�G�,���zo�/UP��Y��p���wt�]i��
�ib�����c�l\P�]ٍ5�+���UP�i���7{UP�VId-v%ѱeT��!f2�q��(|Hl��ܢ�F�ȳ�.��J��8=&7�6��a�p�z ��yH���@���DՍ��v9򤁑��'�t�mڇTS/�����]p�	���m�G<������,��c-?���ǀBa�˓4lY����n��1jG�ο���o���=+��݇��fh�/�N�H'����0Z���I�����o�/�{Ub�J�0�L�.�o�ҷw�5[��
ĭ/$�:�[�00&%ϐk��z�P�Ctuv��ɐ�I~+�z<?��>�n��o.C��Kn��yl0чc4�˱(�������s�N��s�#+?�;Z8��vt����c*�F�G�vnMʍ�ҙ9��ňV%C5�4-y�q���Ф�|=r�@���DMV�Pу߄�Z�Z������źPa5��lj�� �O����*.��C{4�v9�B��T�7q�4�����F=u�)���t��^���cB���Bf�X���C��6"49ohl�c��u_��A�����$V]"w�4�uZ?NN�؂O;a6KD�ӅP�[�����<�����i83͌@?�}Y4�V�鈠4��?�_�E��*�I�3�du�������k3�y����P����$#�;%+��a`�F����u��2�����m���c�{�ͷ�H�"x���!��Ky��g�yM��"�n��y�0�#��{�����vC�_��r��wIۊ�%���]��i�J?`�S���-Ru�'�4�p@��I���ahzTh� P����e���ں���Ǎ���nAQ��I��W�^e�a���8UTA�ϧք~�Vӣ�YSK���gw��lqeTs*8yQ&&e�-��V<^Z��O�i��x<�i��{	�9d)~5��X��y��
dqa��j���yJU�=��O߹�ǣ1[��O�'T+%�y�'b��K����M%�{q������[�C�/��
d�2M���]��/���H�{�V�Y���	҆m#ѺXe���\%9[E��Zk���Tq���ZV�Jǫ�}0�5�R;�t9���_�I�sq��G�xZ-���`^�����7N��{�2��� �+4�q���i�[�����>W�(�K�e`������]=V"����O��㍲Z���2m\�F����i�2c�17�����4`���.�O����|\�Pq���ؓ<t��`l��Y\�{y��Ǻ�t�s� 2"�9�E��q�_���=YB��>�8*)/���#���u6�b�*��
��a����!Y�G��t�E�Q� 7��O�H ���Ծ�T�����������}R�y} }zԾ�"�T��憐L\�џ[�؈�H�܏t���W����y�e�#�/:�~9�M�ޡH WV�{ ��Ʒ�*s�c�K�<w���Z����}��j�f��;4e\�Cn�(de7Ck>����[���z��4�����M_8ŀtOtkb��y���ȚS����I9
g9�/�%	ԂٜS�B��Ḽ���j6���.3��ڝ-"�'���T��V\5~�O��7�D\��C?�f)U|v�)~<�� <�i�TnZ�õ%�r�7'D`�uF�]N��_��	O���:��r�E�jZrx^"�s����B��|��EF��g����mc��w-.V�ƍq�2�N������3�&6�$DTQ�N��EN�tY��N0|�>ٴ�/ʒ�i�WL�D*N��LjcfA`�|�-A{b8A4����0V��?�3$�WpW�&�#��ѻpY�Y�~�p�ȸHg�������,ŘC�*��VJSV$��m����&�ʛ`y�5׫eŰ�*l��I��{}y����濾y�3S���&`�����3����41��=�%�@G:���T�d��r
�9��Ī��7pL�Q�h�S�����D�0�'<���O�Q�9��>����G��/"uaXӞ�X�B}���T{wX���g�TZ�)ɶC�K���͞L���������"�J�{��3S~��&^	��3��K�\зx^h㯐5��F������'k��I���Ɓh����i�nM�y��.ݙQ����0=����TqwL��O���%i8b�<B��Y���iM剩���R.3P>��h�@���zҽ�M�C��z�h� à��n�
"*0��5/r���ء�)Ա���Ǵ\�@���vYv:�e���<,)�E�ْ������?��M0�"�3�*�k�Y�^��a�~E<�ϕ�܈=L O�4�'z��(#�x�*��F:?�3+���\ J���A��Y�ꛠ�i5�=Qg�C�"�+O������:�/z�M(4��ǅ��}?���v���^ks��UMM��p��-;%`/��oC����YX�b�s3�-�0G�"!��wѢ'�(A�eꙀ���D�-����{,]z�a\VGVH0�d�j�,��ם~� �F�V:@Law5L{�w@���<��2�$���\��1'��(����Y�i}y��� `P���dKO���T�H�r�����>6]n�ikMψ��$�Y�<.�b�`��x?.~̄�B�P�Ƈ^����ya�^�ӯ��Y��$��#�j'�ˏ�i���^�m�z�GO;�y�-���o.���+|o�D�4*�gh 
Yg���\�+l���*Υ���fU%aͼ�2d"����w�@��{ĕJe'�Qf烵R��en3Fl:X�q�myuN+Q�0�r�#����.����%�Q�@�z:e0GߝQ�*;T&
8a�]@_��|�~�͎���Z����P�hԥЉ������.���׏�~�QՍc�Q�6<���0���,�I8�:�%X�.��޴F>}�ܟ��5���Ț�o�݇!�6��a�b��6������0�tH��6�fݵ"�s�bB$ܫ�!<_���+�=�<Z�0.�.��쮎�.vo4����q����3��o8��l~��;~0���	bA{��@�����J-��\א)7!�ߢ�dU
�yq;�qJDp�WWp�0���7�t8�� nɵ��3��*�t�7��U��٢���U�|k�~�w�FR��T���PQ%!�e�ct,_�}FkP+Gr������?���&`�Y����BTA�yqU�ޅ��H9@[�5'��I�\���8i��B��UR�u��]���3�{m��Fn�{�B��2���@��)̚�����x�j���<jO�$A��w�t��	4��}�I�o�D%On��p�tB�h��*��X~�K���l0/�j����G8��9T1�E�0��r� �,U=��b_�����5�I�F���\�F�Ut�g�)��.�Y,Iv��K�)�%V�=�{�b�-O��J�H�m����:6$s�#�'h�O��a���li���vc���1�+V����O�7�2ǩ�'9i?9�?�J�R*�Wr(�^\ظ�mڍ9�j��G=T�y3B�$�ǽ�{}���\��M��h!�N���M�f%��ٚA��i�\Μ�B���~���I>�x�Ö�}����Cs����*�_B[o�yI��<1XZa�F1|�US�鿮:�q�4�۟vKc�-;��,�3L���Gio�,�p ��}w\�n����|�'�R�	MZ� �S��
�bhMO=W\�IF�S[X��s�:�F��t����ȴ5z���P�be�ϐ���%����кzel^8$�)mD(7�v\��`�"�R�R���D�n!��z��h7)2���2g���#�O1u���F��ɥ���>�g�Z�`	�E�F;ń\찭\���ʛ�#�����x����y'�Q��Om�|Ƚ󑯡C�~)��ql�R�q���:�{L_5��Ή��|블�
Ӄʬ�⿢u����1M1"(vU:�pt?��
������:]wb�,4�g�VQ\�`$j��/4K{9���b<̺t�+f�V��@��X��{����y��=�	�D���p��c�3�L���<��x�� �q]�����d,�I}��#ۿ'l!{�C�9�Q�ҧe������ؚ����E�ej\42ڳTu�X~�p0��h���i�D.#W��<�*@��O1��7k����kJW�h�����v[����c��З`h?�KX�]��ݲG�����ڂ블w���Ɏ�(!Ȭ������|���$�]���(�|��w^�]]�
������_Ajy+�����U ���̭	[��*?�H�;I.7Yhr��/fca���kL4���Β�V:s�u�b9w�L�!�d�5@��ɬ�#�W�@@��b���QR�6�Z�c����3��C�2�_R�+J�Ez2�U��i�xh�Pi�^�]�O���:]�]�\�)q��j��"�5b��� �n�U�x���%x"�;�
���`�8sg������������c���U���|H�<��R������[+�T9̣�h�>�|�0�D2�W��&;��(e�5��rA|xB�c�>��j��K����P� =k��nS��y[��/�Jz��;P4m6��Oʭ($���`b͌���[h�d[rZ�@���,_>���1�-��%t��(����o���-��Qk�������x���M�kH V&JX���I�_�=�"gD�T��e^+̒N'���:�D�y�m���:T4���u�ρ��k%2�#Y_�a-���j�;�Ր$~C���� ����MP��|f�j��V��ߜ��盟��[�[��wS�4��њ���xɺ*5ա"�BT_/�%J�zұ�p�~�!�?��.I�����M
�'w�z��75|ZlH㻗E.����j�GB�M���;���������6�]�F=�jEI�:L�;�wd]v
+[�_���>@� ��.M6o�g���K����>'0��3:�TB���ت1�U����/FyB���h���W��0�,O��G��J;�t�&��=��-�\4��V�(����ܐ-��FAA�9�y; "��gŕ�׌�5o���џ2 �B�D\nQ�98�uEs?�V�qE�nA����܇X�HE\��|�&�gp:=�)uɭ^����k$����ȗ�Y�2��b�Y�"r�H������w�� j
Р�Z���0|ӱ�L)"�^�7����"Ґ�^x��ʩD�I���)��d���Cwhw�q�Ҍ|���n�i��S����u{�\��}���£�B��)����*���{���h�e����1�e)Ǵ��c�4����+��܌X����.ʽ4Z�u�-I,�_� ;�gR��l����ܣn/�N֝Ȥ�S-	���qv�o�l�)��G�v�����2�Zۚ�`�7�"��U�ŗ@�Y��l8k�g�,̧���{d�u��"�M$�i�����Zza�w{l�B�	�e\a��c���ސ�G��IV���H?JC�n`MFB�"�#���c��]T/���gs����G`��k���f7����'	4�]��r"gwqJ��.*Υ���@u��yX����B�z����
��|	S���f����E�Csr�����9:�%N@�&�9���/��` �q��o��(z�-�f� ��pE�V��J�h�AȽ������{o">՚����v�~�/�ћx;�����t�v'�?�9�$Y�n_�#-��l��Ch����^�X�$J���K�y�i�p��id3d��7�Z�]�z���|���7#���T ��;';ymZ����g�a��Դ�;�RKiܮx�-QŚ���SU�9�&�f�0��;��NF��9��v�K����6dW�ni�ʲ�o O��p�?���^��(�@����U�����}xv�Wɤ��ȹ�e�$�#Hm��%�/�߮��}l�J��[�Q,�plD'i�Ŏ��@ŏ���YE-pa�,vܴ
��kz��+��'d�@f���?�]B04x�9�6�Cn�^i5���p@]��k�M��X�z
�G�M�'v~��:�Q��{�w��<�%M+G�IU�WT#����;�k��H)�!V[���IN8�a�{F���<Yu��g����D����L���u�-p�+���ae{�T~F�[��Os��s��2Qς`�\�Q'GcöT����,.n�L?�)x��g�.-�0�`�����Fb����1���|^��\��@��D�g-;����	a�t��g��N�nN܃�����crk� %�U_W��