��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���1���"ء����ҩd>��g�cAE�:�VH�
���~U�G���(�P���m-*����ƾB����;"���7���3%�
�@DH[��Pd��ʃ��-д*6���o���&�����%����?׶�s�*���H��F��J&p��3,�n^�f��TTP�����s	wup��R$,7�`�eN�/Ԩ�����K���W~�F}���)Օ�b
`@*�C'���%WNB��\�r,�{���t�v����l!4�T�u~�Nxt�F����*��l���<V��r^<�I�6���bX��k�����dA�Zʁ�(�xJ'��@߭�n�F�[U�qE���T@?pP�A���e�� \u����qӡ��(�?���\MG�a�ٴ�{t�$k�v�
��2�V@��sz0�������vV���O����� o���"@�s��Gkf���*���x�D�W�rO>��wA�}�$f-Im��J5=�X�]fZg�[��h�9A��<�}M��3�eB�F`��F6���I�:�)W��S��l��gh���R���Q����%�=��A|E������iy���T��|Y%A����g9xC#O�U���q��*�DΨ��P�����L[��c�jE�B�ϸ +.?D�;�n�|�d��
Z���̍V�5G4��nf�X�X�e�n�!�T? �9�M̡�����ި?�� 	�|<{d��h�s����+dF.,�9_���Ѧ�le%M�@����PYl�y����@�O�*Wʭ�m�5T@�ݑ]gA^P��
��.�ؓe�<z����27;!��g�D�h}+�*��#z�2��">M�YL����J���%�z�{uc|]2Հ�����qQ�ш��)��ޠ_~N�h�r���O�n\���uc�:f�^V�yA=�Jw�=*2�Q/�����/�k��-����0��n}������4�!�.X�H1�����C{�Am�6 ��q,E9>]/!�#�霵�'4���m��� Q�d�I!t9M�͉����tr$%�	Q��M�}��Z�����D�%��Ts��!3
���CB��T���J���7Y�����@B����&J>S`�z��Ǽ��;�_���DlsH}:G��/��/�� �� �}tf-a����.yr�g���K���T|ٍq�L��L���,�)&��?���5=����_p^6��噸�?���$:�pi��8u��!.7���MKǟ������HRej��CU���J���`���@3~�s��x���'Gm7��D#���"��1}�l�d	t��}#����9�1�������xi�mc�ܶ�b6�`�(~�:J��2����<�9سE��hn�]����k��
��r��U6o֔��Cdm�}g�x��	�iЋA�A4�ά~le��[�ׅ�4��F����m!�W�����PΣ���Fl���F���Od�ꅗ[�'��e�]���e
���N ΂FD��$����/T�VIT������j��r�dCy!ӡ�dujt��Eѭ��M��a;�
�S�	�t)�y�
��t��#��`�r�'T�C�.kֹ��>Ԕqh��)%�����V�w9�r�i��zo�ҍ�U��kI�!E�D�ҷ�Y� k�]����^��x��<d��k�-d�z�$+�]���J� �T�T�q���w9|��^��\u��(V�jI���)q���K>�+�h��ͅ~1�:{��]�be\�3v�3�`mѝ���^Âh{��*��3A�/oEkw��`�.&�f��.��X� �'yM�����TEM�Ux�Tot2$
0��/�{@���:-*�