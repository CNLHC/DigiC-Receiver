��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ����S��@$�'z�0��KX�Ŭ��w�z��h���}�D�`w*��\Fi�;0;@	@&�.�C�9J�N�{��:�.GmP�ڍ�h��?1��D�sm�{�%����۳�2+R��xIU#���l,�4J{��|�gޛ��ʆot*��K��½p
��/c�}�F����;��B����o4O����a٢" �l��ʹ�~�*���L%6�7���x��w��j������̝���V� ]�x�	`���Ut���@����Sw�������a` ����TB���(��μO�0��t)��b0��a���r�����K �@�Uc�����^���R=8}ȃ����	��.�q��-|�=�E�aA�����Lڴ�d-�^٘�ZfJ�z�9,Cy��ȁ�n��u�H h:7�O���d6}�`�f�\�2}��ܶ":S�N,z��ߡ�J[������ў%�l����!�E�v� c�QqP�qQ^(�(�NIx'.昒C*����>�%nzF��t-����=�/�?)�k�}��{O�0'�������0����T�X9��|X�K��jVr7$Q�G\�Ij���7cWó؁o�{֭��)ɗ4?Z�-�@���.�����P,�6^�ޚ�|ć��/�h{��:rr8L�Z t���`�l�ɪ�E4(�L����v�d5HH�s��妖��M��̝�@I����0z�n��ȼ�p\�én�a��u�#;{����v���7�<ˀ�P!�C��^��Qsyr#L�Б���<akJ�������eb����YS�f�]��2Y���%l�S����3 4��3��b�v
$O��,�א�U�ĥ-=�t�/u_BQ���K�q��<'� ��/��=�k�����wŰx�ûw�YB�5��>���{���u���G���z��/��V"��d��rRcV�bi�>�z�u�U�m����1d�4���I����Ӑ�l_#�`�+��k���ê���b���@�@�Xf6���s+���r�z���*�0%d�N��h0I91
�ӖzC�����W�`� �U�P6g�7?׹K
�(��a����=Cѕ���Kٿq�Xf��L�b�o
�i��]{ά��q�$>Ժ�6F��1��L:Y����l���\g��|����	��C�Zf����"@#����i>!
��pcX��ʰ(/�(�X_�E2�Z)D� ,�	!#�IO��o�"$}A��C`P���c�4��������L�mn%O��T67��]%�,����lm�PY�
h�~�_���h&���*Oyc���`�q�?�d	g�9�@��֥l�mr��S��`���1�����;#]N���/dC�ٔ�
C:'��gјð(A��5n�L�>TèW��<b�pN��i���T��%$�f���dr&�:?!8��o��{ck'�Q�w-��ST�ni��ãej'�3 c��U����;���H���%�������%��V��hz����Nj�Z�aj~v\'@�%��w^������Ŕ	��f		�-9	�F����@?a�N�4���$�9�@Z����� �#��'���89�Ɨ"��.w\Ҥu7k�&t+;�$ *f�.ȩ��wß�m=�� � %V�d���I(ܑa°�b^����҇(�>�Z�H���6��FNZ�6LW�N@7-z[�U2�v��(��@d��:�.!��O��*��_2�=X�<�LX��[��ђ��r��ۼ�V�U@����cy�Fz�m�Buf�b��B��ǘ)�]o��9!2w7�V�#؅]��Xub좰��ݤ���?�+�6c9��������r�����˝t@2ںMvI���`����3�C���Ug����[���O��n��n��u>�6�C#��B ��|H��`$z����;�ȶlu��gͺ�x�5�/'�L�mur�3/��s���-�z7'�[ڰ�-迨0��݂$9�g'kS�?�J�P�fyOT7vh_bJ�R��t$)���vA����q�C��*��SS����]�%�h5��d�^@�U���^��������X31�I�-V4�R�`�����$�c~��N�-ڙm�:Y;���$y<~�Z \@RQ�O.&L@���ЉxcT�5*���XOw8Ew��ǖ��w��V��Ԡ���"�Z���9C�w,��?��zd4(igF��?��a�xJ}R�睰H�|%9[q3(zR@�D4z~�N�?j7�%��v
>�"<��[F�4%�֙hr�0�fT����Sr�Ch�K��gܦR�ލ5��LCy�l�IA�$��4�
�i ��+���o����Dgm��9F�[~�|��n�Q,� ��)ފ��dV����F|8�qO	�j���jt�d�ɛ��\�g�|��om�y�5H}�:JN�C|��;EWQ����04x2�m�r�r�c����Z�,`-H�������z$�P�8���G���1�� -M$pL��]PV�3m�P�2I�\��7aTMsl���?�}N��_X�7�d�U2t0�u�-^��R����kac��dO�`��<�	v2^��K��&G��E�h�_BA�=�05@����(3�f Ҷ{�1�5��	M�����ӡ���p�
.*���@W;�&͜��c��6yi����mq8���\g����w:�J�-��w�Հ�����`Ꚉ����"#(�S�^� e������-����Oi(��ᠠ�_�
Ub���+2R��&�\a3f���L�nn0(hV�����o��M�U�Y*_(ՙ\�R:�f��o����yHxc�����K���LB�^n�ZGeқ�ٙ\Җ~jN���kt��
�i�a 𨴂�=~��`MS� ���|��4�X�T��{��\֒�09�yўIUPKɥd�����k�=s,>��]-~*�¯�1����ǹ���h9�o�EJwC��yHO{Z��yo��%z�)N�Nڞ�1��+c�8;%��`4,�m(ڍ���TЪ�!(H5m����?������n!D���}�4���U!�7r�Xq�>�\B�v8��ܜ�"9�q�é�g�R����A��hs-2�M� FP]T�