��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���߫�.��&G��[����zPף1�K؇*���óǋ/��d�?)u�,ov�	�>eaBW$-�'������X���E�A��	�y<�1k�.��4r.�&)6��BjAܭOD���3�=���S;��!� �7�J\�n������0��4��J����v���Im���@���x���\�RWܯ���w"����:��?}�i+�d�W�bm����[�_X��C#Z�;
�C-Cr����J���NQ�V���e�"ι�a
UV��ξ�j�'�K`�&�c�
���45r޸�I���ti��BY�� ��9j6�j/�DJ��4�'O-���]W�Q5��״��%g��ܪ��&���E��ʂPJ=ð揸��h�����_���[{��n
Ee/�x�����x��XxxWL��W�;��k$N?E����^�)������}�7�%�}i�vk-������z9�|�A|�3(�M�d<'��؍�$�y3o�Cxp1���PЙ�q�:�-��r�މ��T�X3�����+j�1��vx%��L��Т��)TLa 3e:l5aCecj�BJ@�Wߍl�T��3����dX�e^�U����VCR�C��2��j6Ox����h��V�R�Y�*c2�$�B�>������i,-�]�%��'E��ə��]�F���R��y�q7�5�K�������6@�ۏ8m�����9Z[d
%W�J���	+������=�eit�f/�SH/���f��#}ѳ�f�T�e�Լ�y�$�{n�8,����O��|�2!���Ip,%Napu�����Ǩ����Ԕ��j�6�7������;�脺�qc�d����KyPf���N"E�.bv�ƯVؾ򭝮��7���׈Q4r8P�%PzQ�����ˁu�?wց�x������A\�������<+�X�^v��6��*�Tp����a�i�����[>�����\K]��rY�¼W��s�h�����h�tC(�6��:E^2��#q���)z���R���
MꞒ�Z��!�������_&墻boT�]����4�j����b�Y]�}�l���"P�³�2ɾ�m#��&�>N�y��޴¾"Z�5�
���D�MXV^��P,����ѯ}������ӌl��s�i9���0�02q�K����1�vj/P7��͵�X�j��N�x�z��|o�z*��?��F�p����龝��N�Ѡ�|�3՘O�G��fT����{���>n&q�)��?Óf�Ӌ4�� �!.�n�i\
L�[_kFG��A�	If���u�n�|�>)�r_]�����Ƹ� 3����F�.В⃜�~��,('��&sPե&F{�'6������ge]���a���L]���M���ߣ�c��ƥN��bYM.��a���C
�7,���.�	��o=>f�������=�z7ay�:K��Cƅ�Z>����D�5}w'T���K��i^^���4�1��W[��r�V�0=
h;�`�ciJ*蜥��Yr��-�LqMe��S�KaK��aA��ё���o�Gz�[�%�CgJG�0"<i��PքCۜ%�:��i^Yx�7�` ω��'���c��k�����\������&Bx¹1t�kRhL���vTD�b��+�:,��%�n���1��kP{7j�EeB��˴y��n�����)t��1笩P�g�6�<y1-uM�K��^'�$��ؚ��&�rPہP:�y�2&���`Il!�Gw�\�gM����"G�,���O~�D��.:�G��<��E�x�g\��&bJ�ѩR�3|a�9�Oz��&S�e��1��
���7����i���ˑ�f;!��>�9~�@x\��Bx�O+�i�Y�����}Q�Ig����^oT��]s��	�S7=|�OP��}M}P���p[K��-��T#5�qtP�|��S��[�@�	���I8�O�j��Cu�6#:%(��ʍ���w��Mc����nF��0t�c�W�rU��r�5����N�Wx�����I��Px{躳��1ڮZ��4�U��aֈ�4U�B�P�5[�@���T�v+�ĺ�.��U
6#�jn-Gd#V�����%T�J��(���yN��K��Fwq���"Ks�!�ұ�C���gE	{P=`b�_Hx@���W<SN���w�C�i��3&^cW��;�@�.lT�r�����+�_���� �Ë���e��J@��֑�d�am���kTN
[6�gG���G1ݱ\qs��t:Կ�$Hf����*�t�Nn�0��\^��@���DΣ��K�vg<�I�	8&�,#�o�YcD[��n��Bc�(�	��mMJr3��l�5Lb�A�"W�G;��/���Ί��}| @'�6;@=Q�#*eX�u�~�X:���(�ۅe�P�e�������~SWܥ͕�⡖z��>z\��?������S����6�_��ט�;|JB����`���gAz� ����������-����^�28����w��^�k��N�p}�W�L�,VJ�v6g" �w��	�^���B�V�3�{��+j\+�KI�T��^Q�t������a�-X�VG�}����,���}V9���)8���:�^�u�������]�PM���x[j�+�8D26Vw�����TxZ�IX��%c��_�A��jd�k�/�dMRjT��N)y�=���?F�
���k6��:�U��ow�|��{l�)sJ�״>]��!��7]<�����)��W!�Ԍ�=�������1o"e�7.�.���+hv���v#&7�Bi'1I�c������6E��r>ȸ�Wl��bDO�qT,?�ɏ�{�_�Vq�#Hxx9̺I�#�4P���/C8�e�?yY#�+bL�j���j������\��g�h�e��L�Q���NO1�>9B�W�hOۅƌ�,p��
���}^�`�Ô�B~5�j����`��~ �A�^A����u@��H�`+I�������Vw���7��+�3�����t��w٘��a�f8@�t��t:@Ľ��u�p5}q�<��q�R�H�Cx�rߓ~'B���!x���ptS)�i�(ⰼ�� �:�9�9a���ֆ�K3�Q�5Ѧ��E��L(�����@���jWy柡����ֈ;��^�)�	�@����i��D������B�zv��l�S�a�!2��.>24]�^���l4���ݤ����޵5 *�(�o�AI����Lʏ��
�4�`�D��"�>(�%-�㿘���}.����^-�+Xe�y�<]z�xF&>0�䈰��K���1*33�F�j�6���ѩy�����]s?��I^k�'|]O�e�f��3��KA�a�bD�D&W0<	sp�����6�Q�5Z(DW��kK�S������Ĩ1f߲��ח#�9\\o�"��N�����͆0r;��JIĴ��j�J��[����߹�B��1*X���E��]$�3a�؋1h���{E�v�乎�����2W��r8o�b���0.���}�'��ܩ[�B���-Ϻ�BHV������$�u�ڤ^㌯k?|���be^.��}@�����?�u�����"��J���x��:e��YE�hp#Z�T�$�b�(��!��+��V�4����@1k�����;\����eK�̃�&!^k��k��k�'����C�)9��4�5̖�B>f'ܵ��!�7�����n-�
��@�T����:�)�x�BW����Fg�?Qp�p�sf,n�jJ��ءK��U}���}�G6��%���Ӊ2ס*�-�?ť;���q���<�L�4�8v�#�����Z��ǟ���Oΐ���\�бLW>�v���~�)ο�Q��gG��jR"P�yP9���rv�v���;�?� jy�g
C�M���%��h����j9)���`�5���}�!q}w%V.���r�r��.Ę���E����!#5�,��g7�%Ven��Ӗ��k}W1����~	����( 	��:zg��);���d*�Ɲ퐝��c�l:��G���2�Ok��^swU��	?�U��gr3������&+84LwÀ#�i��s;�p^>�͠���K��,���,��`%�4�/̲A:�Z	p��J9M�o9L:-Qsy�:#�+���x��2G�@+��� �0̀�C�*$�:�$�Zcmh��;<��<���De��͸~�%�Y_��gq�h�F"�8ë$צ��f���iʧ�����/�<���^�� �}
�z��E�3��w�]QW�w�n�
k6<�0�I�>���)�F�}��v��^��A�ɂ�R�
t<�%�]�R.����k�@
/��5�����o����rq����NR.[���-�w2���?�tj鴀��c�;fYF�H�]�U�mʫl��-�m�:��}���B��(�^w�4RS+c�`���)tsa�
(�;x��˝#���o��/-"�X����� ����XX�x%ՍU uB��=� ��N�b��P��]M4�@Ab����
k��B\��i���)D�c��s�,�9��t�SN�m}}5� �<"(�!�L�:4@�>[,N�����?�*J�� ��(v6�6\ߋ������8h�?���@e��:�;��e�5�Ŗ�MO���ս<��4ہ�B KI�6J�t�k)o�6�<��CX���$z�Y;ZhR�E;�΀����g�䨁S��k}�LkRʐ���wi�p_�7��`��<�Jf���.�
���g3���k0-�^�,.u�^zp��3`�� �v����ޅqH1�ߢ�O���{������DFGP+��~��]ӍTq3�.��pÖ�:�l}�H�.J�D�|�Uf�xA���>�G���=���4��#7j�&�5���m��M�&�%� խ����#��a�l�*��[��0Ǩ�'R��3LY)�m�Z��݋��C?���,�($>�h� ��-C)M�7]!2(�x��[�`KcJ}\g��}譎tt6�l,X)�vQ���$!������V�Ѻ��a_w��tlG�$Ϟ��F�B�L�&�2�\�5� �����²>V?kEF{3(G�{`�����D�0,�[���uvF~_��'	�Gj�-��R��5������������,VRA��n�,d��I��pՕ��������[/�o��+u��E�c�{:ǥ��ٰ���M����k�k�>��(�6@����۫D����u�PdR�����4n~0�m.-����*Ǔ~P������}��n]����.�
�� &���h�j��g��	�4*��C�%_��t�`ڽ�3�:�B�G�����O*sH�V$�j��s;ʹ>�.��I�z�+�/�>:�<�`$��_��O
6�����~��ȼS���h�l����� }�wl�}�u�<�X_��N�����z)��h{Q<S��f�G|{Jf,Pr� F�jEvH�h �.O�
4�bW��i�#��6V9�����J��I��ގ��8C�;O|�}��:0g�K����ґYٗ��5�V#�X�� ��:�,�[ӵ8$,���
���L%#5:�V<efA+fW��0�<i�Ų���To�x[�s��Y����_*����"|ZU8� ������)����0(����=r�?���X�ybQg���s�]�4�k���)7��������֞��[el[0�����j+%���J%�˭�@��7O�����չ�'��g�L���-���V�
7_c��.+�r��k��%<��D�?�����hw5�e)D2�0F��Ea����&g���Fj���P�J�z��=6G�������
��V
��2yb��%��ao�D�~�\�~QA�Y��x���?K��v{a��s"=,ś"E�ƞ<^k�an�^Fm~�$X�������8�3�!wV+��i�b^�4>�Gn���j�f=�ż�cz6h�4M�h�����@ND������IL-H+�}�.��L&Cʂf�δ'��\9���!���ݧW���#m��x��=#���h�ʭ��xu.�a���(�|��ˏ5~��"�h)�{b�Ҭr�����
C�d�,%<
��[xF�CEoR!��p(!�(���q���j �
qN��z,���z����ѣ��=���b��A�&6N�<[��Z�uUa'��\#����݉��~POb��c[|¼E�3��h�S���2s]U�.{$?���:��L�-n�3eF�S�z/�Ak0��Ӳ�ڍ���81�7}^�_�����"ǏDMT����8|�ݕp1,�c��h_�Պ?�/��ݖ*��-��������L� İ#����`$_��o���޹�/���'���u����uv�D���IqC35�֞�f7��f��j@��}Z�T$Ĥ��p�8z�ƓE�l%��&���z�#j[��&�c0�o'{�'o�i��e���y; ��"#1���sܐ�&8�� aι_�H�9Bm&����;wXSE_�������č�=��s`,'�`]xb������i���X?�}t��=���A6��4���@t�z'�?�h�����	$�e�ʚ4���1���]��4���:������'�`z�<����s,3���f@��[�=����p� ��K/	_�!�b�OOȒTH0 ^�}D���n룒gW�����O�oY:V��nC�\t�I�GG���6����t�p��+����Q�����A�u�;�55�{��Xc�B>������[J��5u�DhP[<|�!��QN��5@>m�ZY8$QQ�Y܄�L#�7?WX�o���V�2�6�;]AS�| v���c�#T;�B�W@@O5�	ؖ��	�Rw��P���&}�r<��S.�P���."2?%U�mݸbAZ`�_{�Y�&��s����.����H�6����h�[��kj��/��A�yv�,���U�B3݇]� �-��T�Ik(ߜ�έ���]�ѫ�'²�5�v�O�]�Wը38�T/��^V��O����ҍ ڎ�I�q��}�IU�m�'z@�Cj�,�[�c��2l�1�U���LtV���c%M/(~���*�7݌���7���Z���6o���^vЖ��E������\��ϻ�ZL�)Xv�~>�r��!id�e��s7�'�0�\T�Au����@!R�𤔗f�W��������arUh�E��*����侐�.���bg4�Yf�;)ȳ�5w����Aϕ�TR���P�[۪"'��;�P�DW��S�B��{�Hǟ#���L��P� ����vbb��j���2�-����g�*�]Hg��X��"��E?3�8W;�u��n���,����MA��8�2��Qx꒯w[fi�/2GN�J��uk;��b�C[�-�~�&i�U��h�a \�8�;����qr01��b�7)@��}�><����A��!�cyZ5�$���}�܅�|i�sSw�Gk�&p�T��*M%F��f��V�rT!A�6q�߯�g�`F�%E0ﵛO�ܾ��ηL�����#�^������h�+�w�X��e�e:
�i�
�f���w`���/����۳�cW�Fx�8h`�+�R�K&3(/����3E${�#��1�kK�����,���?4���",ⵌa�?��q�F�YT�)�k�����ǿ�FΩ�Gz	߽gІ9����8�R.�C"�%�"��H��w�I�N�b��(W���Q��R���^U�m,�w%b3�VB/��(w¬���t�l/�oɆ˴{9
�/9�v�hy���a�vfJe�'�'<(*J:`e��\#nE��)�Ў^ d<������>��y�y��Ʂ�3��0���n��>z��.0�H�Yz����X�a�ġ�C٨XEd�KUqJ�m���5 J��	�Y�8�x[�m ��q�|�E[M)]��c�b%�`�J'Î"(�R��a�0]A��*�Ru��U���@�p��ඔ��;��Y��K�	z$B�2���
Vb�&���z��q��n���dw�y������z�r�x_Q��Eq�=Z�/�'�P��0�r:J�~
VhN�q6,]��ɂ�r��/�����(�GR���̵�TOd\_��j*���p��rs�^�7��=+��~����yإ2#���6e��'ǋ�;K��<�Ђ-�[Llb��}LfSk�-��~��]pF��1�P�Y���#�]����e�`:Ꮉ�2a8�@����D�# ǡ0�P��M�@�?���`�8+S�%���c�OS.D7x9���E�"r���\��J�Q1�~?�T�����Lڟ�Hd���3�lic}N=�[oQ�
����'��|C�V�Й���Xǐ�Ӽ�#-��)�q�p����D��|�kj╔�!�uq)s^��,�kD�z)$S�o3��a.о@;JڶX8���:#�C�^@�.��X�}.���F���EE2��3̜�� �aQk���u:���Eu�<h2�a�ڳߢV}�����P��XD�֢BO�{:�r4����|�H��t��0���w��9<5>ו��A�PF���kSV�׷&�.U�ئ$s�O~�8�o����'�u��M���k�\�U�2���0��q���;�����(nI`Vi�!ͪsÆ���%�B���O,�p.z��}��qIJ�YL��&���(�c$<�=B.1=�U�H�5�V�@�E�	ΓI�O�vM	�,����&BBr�g��gUYg�^¶�t�&���&z���[|"��7�~�P �	���:���C�n�Nw�r�~�~`c�D�bat�I�Å��gǠw��ʜ"���W'�O�V�m!�8I%�~]5�lYx' ��3��e�{̛��3K��Q�������A�ZTi&_B�u�}�n�&��*��R�#��py2(/�B%�?�+���gu�e7)SӥhE��{�>e��of��r