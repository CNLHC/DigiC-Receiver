��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M������O���R�$�lIlqֿT����N�B���Wg��i�ٝ#ei-�#�D�ዣ�I��n��Ώ!Hg7��@����!�`IHiF�JR����`��<I���v��n}�^�@|��3�4����K1�)���Vq�
V��������'�0࿥�>Ȼ���x�2CH�u+}�h���I�h���:1�>��οL���.��UQ���]k׋��"�s��+��q�.�ׁ��̣��Ѫ"�m��C��.�6�;�qa���Ħ_4��;����������9��X�  p�:������ՎE�yņ�KƧk�n\4&�^
�&d5%t'��O��=P:��V��LN/a�������um?���:o�O�v�@��&�)y	�C�y��[�	Bk��f��\E:���<����PX#of�E��Z�� �h�T�<����Yu�&�x8��g�V��bJ�z���Z�{�&��2�;����"H��Si[Tyӌ�p�����*�=��G��ڶ���h�	��!}=�V^
Y5X�)	�A�8*zO^��)����m��,(7~�B�(�D�,*bn��x����#"��,����!2(K�v���ߍM��)aI�IГ�G�g~�P=��dMA����"j�?��)&�䆾-=e��m��K��0�U�.�7���CN�	G�Y���w�K~8�т�A�]�R�t9��|~l�d�_i�E���->��J8mB�C�ߡz�B�6�N���G�$��nW���v�Ԇ�DN)�(�@ٛ�3����i��-�s���KL4�1�
����OO_�8i/�����g�ζ���������ݎ*�$��@9�<�ac�H:F�]Mļ����b �i
a��-9��	6��Za%�*s�G}5}k�t�K�z�5äz���PT�<�a���{mb�w�M��C�Ȱ�8\�O�$���H�8^.����>JPD'\��j�a
�#i"V'g��L�t��	=�����r��.��cV�@u��)��Y��nH u\5N0����49j�
mg<Z���D@�}�uvo�в��[�zڊ7z<nq#I��j����������?W�d��rfGR�̄(�g	�fQj*��PYZc��Ըc~@�~���r�N����'��xPe��:�;�a7�qWg��e��AZ�K�@LarY����!�cڻ<�����B�ʟG����z�w���^�G�-@��;DtP���c�j<���C�x�0���\N�>��IJ̦�����LǸ��±݆�=��f@=r꧄�Ӱ�ƚR �d��;�_�IZ�1����~	�Ȳ�N�.������!��]p+GЈBr��ǔ<���k�0m�JU2���s��P
.j;��~���R՜)����-?�����N�
�� &��3{X�ɠ
/+z���샳9�X5n@\����aeu���繿�PI�?��R1!��uRtLd��>Y�J��l��<*C}(D�r�UC8��sƆz�1��W�O?E3��Ɨ'��x,�畴�Ɂ�~�o��	8�1st�5_�����"���&8jz�,7��Y�lK*ߧ_����y�z0OV�%q�a-��"Hȳ`�^EEN�J��}��Bw����)�)l��\uN�8����[/�ӧi�;��{Y��i�W+t��šW�ܬ����+�,a��c���Q��W�����{h��!�>e�lc��
%��B�^9�{-�����/��u=ر�t+;�kT����29,"Y�����q��\ `�Z��l��Y��1�qC������]�V�J��������l�^�G�A�=���ڄ�|�8�yw 	!*�W�l�`����Z�ٛ,7,�P�5�18��E���Z\ҏs^Yu~�cz4�
7���	��!&
��^���)l��<�=5����8B����^���}E3X�����O���S�� E��N�"Q��FK��y?<��+�t��[�-�6f�l���,���i��G�X�r���쇲�A�����kM��ރn_Fh��I�λ�@i�p�4rVu+R<גV���O�m��b��:��"hTe��gkhDl���.C(y-�MT7ԯC�9��(�Ē��@����0��%�X���L]�lM����-X�V<ikah��K(մ�X4Qݦ�kh�`��	!d��m��	V[�+�#�E���Q��D5�&����e��_F	�0}d#���ED{�"��DB?4�s&�0������0zJs��y�)�ڭMd;T������2�Ԭ���%$\o�Z��K�z����h6~~��ϸe�T���f\u����Z�*}=[�D��R�¡�;s�&+���=�Q���E�������4,�]&��p���)!v<���!_���5�5�^>0OxܩP���膶Y�M������h���+��k�Ӛ���������y>x�KRe����.?��G��^��>�e�鬨{U��徭�gF~����8zW�;f�+���vI�s2�ֶ3ۧ2���߅�'.�	�(Os�R��� ��w��I��M��Zuc�gI��2��Ж�/�����?��-H������Wh�^�Mf�n�f��fO%�QSi`�۴(���ۏE7�',/��Z�X�~�v��"F�0
�o8c�l5 ��ܮ+H_X�Q~r�ʢ*��0�)K�5�������m�\�P'�����Ú9� �W�������2N��p�����\�(uC������K�v��A$��b� B4}�n���p�KJ�	`���m��+ύkԒ��{W���z������yз�{N�{ޕp�l�)�>kL����R�1b��;A�J�I����i��V�,��eo��FeF����@�q��k�H�q�׌�M��w��.6���/V�#5�ZjP[��A=T��lA��Z�%9�n�'8Y/�ٸߟ蜅SI0���17���)��up���q�R�N
��u,d=����v�\�$OPS�DԢq�I�O ��oƮ���&�tޛ����P����ɍ�^r�S)� ��/���W��ݍpy�������"��Q%g}�%<&��#f�ߧ��������ނ%cxa	
�\���/���E���{�*��,�Or����_�YO*�x�'&��*��`m��f��=��{�t.�9#����d
��Iˇ���� u�@L�3��`���u�.��<3��mz"(}�)ᤙ��*,�Ϳ�iÿx'�|���L�]�]c����e���j~���%�Q	p��QK�;�u��	���ğY̓c��:�;¦��<��wsB.��I� FE݁a8a�Sm_'�[���2W��0�ìw�m�K�C���6����x��~�5�ƒ'퐆��%cj�[Y������ߏMDW����%�10A$E� @�V�,�����v��,D�b��}A�(cq���
`�4h���($QV=?�7�s��x�������f���f*V8f����l:����HF7`�QM'�u�t;�k��ܜ6�i�SW�R�`��/�g�|�v�m��zOTB�\ �	81�ټ�~x�̅ܗ�)�1��G�Ϯ�w=l!�9�.4�L��3�ZZ
���Xq߬�ۂ�T>�'��P로Y!����,�h��׆��Ap5���>������)9ZHk�&�?`�	@�{1�%�"�ǔL��C����`4,Tt��+|��>	�ȷ��b�����(��������(��խ�+T��$�B���RUu'0,6gt��/�ڭ��5-��#�I����Sg4�R��9���p�����2b�s蹷K�
��um�A��+���9�ے[W
�=���T�ZFbd�%v�]�uq��9����/�t���%|��!;��]���}yi��G�׌C2��~Z��^y���������P�y��	�?C9!M�]B�0���V������yb��g�����0���H�� 2��PJ{4�H�?M��n�Y�lV9w��Gm����mޜ`ǋڬ�f�6>���	>#~�jҴ3צ��E��������K���IJw>���3�J����H�<�=�ò|�O�9���F��^��oB W� ��.y�Ci�Rd��U�J
wl�Ɯ��l~6��Z5���� �,&kU2���q�AqlV/����-d��&l�^���R�ǩե�t,ֈE���"��������'b�il�/*�d�&d������Kf�u����i�_ĸ�"����-e����v1#���|��6�C��Yu$��Yz	~P�QW���f�����ՙ�6���w/Lϫ��j5������U(|�y%�{�O�=�՟�|�&.up�U���׃t��5�ϫ��_�ڻ��Yҕ '&�N��{m������9�>R��-�u� ���)yh�"HWC�����b��2G%�2JZ��F�#��|�_MY�u�R�G���2�y�p�q��fiv�R�g��~f�%�s=�Rx�7&�H�\��2<�AIRi0,�)��C!55]ź��@9B���u�{י��a��H�n�f�\Br��V�ȗw�
��������ಲ{�}�a��o���e�?2�P+r��~�����,��ؠ��JcS\jlL�ƍ����g�X�;I03׫��Zy�?a��� P�Z���Eнhr���7��"���=���PP�1��PR߼g(Yo���EGl��� �x�z��4{�H]�P�z;����ݬJ[xݮ��@\e�dy	�c>���8,�T�ߙ苋YXd0p䗄���7�!Kٍ�d���N�o>G��;Q�)��ddy���k�n&ZϘ��ҹ(!h]S~��H_T�\��L�L��y"Mj�&{Xjz�G(h�g�x�TP
����Zd# ��KnҞ���~����Z��Q� �^ZZ`���O����g����G�-Цc�HҢ��ϥf�{��3ú'KJ�H*��T���N�Р��T1r�<���j$������Cm���#�k!<4w�v�?���,�h�N�3�R�+v�p�Z ?�C-X��m��ӗ��\I�OPe`d�?ǽ�站8W�ʺ���i�
��zl��L��z��O��O[$���~�H؉�GqYQU�ltԷ
c?%�b����"�Wr��Y���NRfݛ��2P�g�w����w����q[7�*���P��@��_�ɈN�F�4*��)f/Ѕ�0�^������n�A"ʣ��kQ�{߿=iv�����o��	JR���f��'�l0l�Gn�aW/�����t #˧�@=2�)j/kԭ��B������"��5o߂Q���Q��Q���!�e�;�ͯLY��IU#�	р1N`�{��󰋀�Ԃ6s._����[^��J�>���q���etM�U""�F��\�mHc�I&� {��#Z"D ��L��w]�V�:,�&������~�� �f�*Y$6ؕo�=4��Lƞ�i_s+�0��<̈́i��]Q/-��������S5@2*$�Ꞿ��-W�kW7��|�P�į&�H�yXޣ<[K�;d�V-�L'a?�\��rN'��3�c�y���r2_�A�l���@e�:@������*j6�@:f�ٰ��-��2�5��1�B��kY���,�]�(c��Is	"�X����^8b""9o�q_4��K�C�#8��b�Y�D��?�S�*V�v���F��3+0i�~��,�^QMH\���^�G�dF��zQ�+��p|*mu4�d��Q�a���Z]��T_QR�X�Fpt�ߡ��쵪C��Ҫ�er�-("<\�W���Ǡ��GZ:�HA#�Ï��0Bcd�U���#��r?g��"�!��Je֣ʝ�F�f�N��W�����C�����&_�}ь�粹��@�:���l��Y�-��
�Z�(!�]I���&$�Z꘯���A��^�Fk-@
_��h&s��Z���'���+��a��;��;)s��8%�
��f-W�>	Ĩ1�G��un��'7�k'�B��s1F��G���
^74X�Y_��C%3_v��~Z�<~�W���[̞�VJ�g�9)3�����P��D��G�K��[ /��=��"�!Y�>g�H�~�Xn��<�\�n��SuO5�F���C�c�q)���۵;����^����nH�Lh5%�g9��!p8���h����C�7f�r�[�=�H�1Z���9��F��ޥ_���(j���Dr6�QXvԵ�+��k�<�$�Y���-��m"���_�B�c ��w���C���B�D�ՙ�_v�Xzs�5� �����ѽ{���
��I���z��ڍ��{b�Dp�q$J;��#��D�3�G��7Q�F(P-��<Zx7�I3¥����Fz+@I��2U�Ĩ4�߯�0�^C%T��)+Ǻ,͌m5�w��F�A##�*M� lp����j��ny̗q罶3A�ĒZa��"[�ê�J	u�uTC3�ԝ�F_�R`���~	)��u������6h��7U��[����_);(6���Y�#�8RzOS�3n��?�7q���R��wG�q�m��/?=7�Ze�ƚ�\��5�@1�z�8�+;S-��$0ƶ��� P��vO�g��o��|�)�U��Ǒ�yB���F�����@��"��,��<�W�����f+͓�uL���S�`�R*2�3	|�0��������nMJ2 �c]
BPA� �]$��ٞ+W,�H�!���qs�k�["'���z��Q� ~ T�����3#�:��HqjmQ�`�<��[�ġĠ��㴃r�)�e�/+���m��9�ڬ�>��K	hȗ۽V������������X�-"|���2+�0�ޖI�Β��WxK�/xH#\+D�j��Hn_c���u#�y7p�	}��r B&�i�p�6R��h]#�u�f�����'Ro�j�C�J�I����vϻ��*�MC�}����
*.t<���(önym�*w �ؒڙ���>j�wel��y��/�����V֌�U��؀��डRGDb,^���i�B�0�r��ޠB�;�߃N��:2Q=��L%w0�0���yٮ
��((��]�g+�Ca�z�ax���=�t�&!�l�_�[i��o��k��L��G�xo+A��e��kf�ʔ~���!�SIyʉ��<�J+���� )�H:�z3/6�l���<���Vp� �+(��v�����jS�����.;;��~��V��2�?��}�4 p�j	1���;���Dgv�30��hIq��%�¼���sZ�G�Y�^a�ƸoX��/{��$�Ԣ%��6h��ݙ{�&�&��]lz�=�ioG{��I9w�I�G��W�`r���}�%>p�Vq��m�@���r���0I_I �<�"m~��r~v�
� � d�=U@�Z�V����DҖ��\�>n���n/���4B
FDm_�$п"�/��S���h�+)8c�D�+�_6k��l�&G��ԲX|�h�WY[oe凔:�����B�!;.�9h	k�Q����E�1�^l����'DhL�g$�Ӣ���<���l��u6`L�l{�-���d���Je)�1���
_'�c-7�V)�G��FQ�AP+�m�Vׯ�2N�ŀ��u��cB�5��
@���^��$ࣽ��gM��l��5��Drt:��^�9�XfYQ��F(����"F��.��׋���̇��[�WquW��CX�D��"c>��8��1�2D7 Et�Y������W�·h�RI�ut|��q�0<�I��N+�d��3u*M�n�yv7z�E}��c"e�1:�x�͈=�ܞ�|��j�c/�L��A��ÿ����*n�ResX8�g�n�U���auE6@e���K۶9�f�g���9E��S���ڈ��i��.~�o�e�nM�+<ܦvn��[_(%�S�X�1���V���V�8]�&�3�i�
u�aAw��\~����JZe,J�q2H�"���q0P}����]o5���w�,r�c>����A�^z:�����B�k\#�b�������W�>�� �h"sS����+�4.��eُ9������OU�2�
�}93�LDCGB2e�G� ��\�zv�
�=�7���Aë~��
��H��P�m�/j������@�	��M+�?�	3�?��� PMO�Z�ծ�����#Y��#������C�6�c;�mtK<�	�2�e>�J�jp�[X͠��A�4Od�G(���E!�����!��ʓ�.�#�i��O�!�}�d���%���F��%4�	${���ҩYze{kU�@Ӌ��S�b0ya�(�˕&X�[�U��C`j+S��*�zHdD
P�|�{��S����&��\|Xr4�R�[K��<�����~&C�I@�V��2y��gx'Df�_�������7�u�[�008��%.�O�����5�{RDD1m�E����v���{�m�'��L{�;`Nz��,��h�j��3�/��ڱ+��n����}"���ܽ�g(��ij�lJ4�(h�?��}0����%h ����(����A�.�]�Z�˥���w
�Jx���q��c���������c�<���&����ί����4�	{X��Y�\�M�P��k;\-�A�/p6�f�����\�����[s^���FB�9U��f2!�Kt�v����kq��{�++	$27��Eܞm̠�J��Kqz_�U�M�g��Oud ����*���I���p��!$٬<����k�}�/���ŊPSc�B���K��YHc�X{�ś�#;-祗�pe��`Ly/26&���?8��ͽk��������0A��h�ں<3jIJ��-y���0�A�qfy�h�;5X"��mA�0}�y1��Y��/7�	��k�y�G�D���/��NW&^�Ȃfױ˭+6�iyV+w�oz��d���yIJP��( _�B��!I��C���l$�6�A�ߐ�����>^W���'E�3o��d�)X
��ѭT��3Ҵ�:]Hs���S��؋.���UBi��H�/�ߤ:�����c��s���M���T	Г�qD:!��o�����kJH���$����;}�R��zB(;�鷧A$�}�9��?�e�a�6��;e����N.$,]�2��^�d�� �Y�:���N�0	�]�χ�)�u� d�g��'UJPV�Q��+җP�B�?�䁆���ލnS[��ի15灎7X�Ζ�,>j���Bz��ā�gWw3��z��N`�\?n���䬏��@��޾�F>�<>9�0�Y� �E�n{�L7���If|=ڗrt~�Qj{'�
��F�����$�1"��ai��3*��I�8`{�P�r�Q|�snye��p�@��������J� ��#�kQ"X�쌈����&���\	�j�1�b���k0&����N9��Yz)=
ҽ�@��źYzc�x <�w�h�k�&���h}^��l�s�P�1���I
�/��Ee_��^Ih�~#{����b�������^mbz���7#�h��_�a�}l�����.�-��pn�(�g�Ix.�GE�~<�j�YzRYC'33������]�M(�3�Xk�
��b���� ����������y�Hq�(�l9��8��!�K��c��>��@����ɂ�� ��AE�lF���܉�+����ご$���њ��ă4YP���F��RY�B���[�Rb��f��4{�A��_�<K�~(\��2��H�U1���Fk���T�M��M"9P՝j1�ToVӤ�Zp��[��^6�6�3��ed�p��Nٲ�� v��
\���+R�SYYҥܦ<2�j��/����R��"݉b�͂��d�
G��4���ϣ�OiBe��-Y��ÓɌ^ʰ7�ŭ'�/�&.��B1P�1�8��P+L;n6�!nz*p��t�߇_?S�������}e_C~� �&e����E��C�����/��ωl͔U�^k!;�>R~.�T5�6�n�D���g�g::V�9��y{�gg����������^zZ!M���8B��ꓱ�jx'e�N!����"�I-�Z��3S���i�~.d���		~ߚ��H��y7�2�싚�g`L�c�ت��y$�O�
M4w0��W'�?�*��4D����@����d>~�fx�~㳿�:Cy�7�)�5��k&U4Dϵ�1OKS{જ��B�bI�+w���Pr.w�������h.�`���?"�͹%>�f8�Ȫ����� FC������h����X�G:I�0ZL�۶D2�_���#���D�ږw��/������r�nJu�$�-�L���<oI��h����d��u�عb����C[�<���R1h���ukq}�7&h锲�D+p�t���jH��F�����G)���o'O`v|W�v���'h��p���=�C���i-�&Z�9�1+砤�)l����j�2f��h�0C� VԾ�ۓtD�]1�{��[A�z�3��}�	2d�M��/��J�,?5�Z�
W�ߔ	��7���@¯�OD5@J#�m'|�]�xSGSE�-�|��!]�$rFi0�L/��@�1�������l:{���NG�����Q$^��-2h耍�6&����Ǳ���Ewx�Km��d`���9��}����ĚC���hdZ8zw�	�$�Bb�
/ff?��B+EE�%+͗�{Z}�
 �#�����}tdM������-�#X�21c�X�9�|�C��4�tQ[`��b��-T�o�B���%h�l5{`���mJs�*��9F��F��	�Ԗc8wף�H�< �5C������'���?�c=���0�"���4��/j���S-�f�L��j
_�b�hzRP��^�Dj��n*�_+��O Q�����S�SC_�{&�{�vl<h�lT@J������Pb8�*����9[Å�)YC�T���ʑR��>H�ED�a.�_��SF��E'mC���jgJ6~���)��F�r�B��s>wW�ґ�f�?��<�%=ږ��mP��HB8�;���,��cǱ���R%W���[2@�<�M�7|����Wg)�԰ͭ��b����QХ��Vw%��^��V�`n?��Q���4cJ�=�mV�N�ĮD��>��Sp�~ |�����Gΰ���|�q�.���3� �Fp�0s6���<�ć����2�>>^-u6}(��xιY�a�"�Z��{�B�{�,��%�w��E�c8���%�!�h����I��oV�2Ou��׭A�;fk:%W>��B&���U�^U�S���I:D�����pQK��.R����Z`�W?M�E�6|�YuL�k���UJQ�k�@��ľBΛ�G��,]*	Bv}_��hB`�B�B>�h���O{�����d�)<M�8���xK�!e��i]��ʮ�n�\��C> c�	�xv+t�>-K�7�&�g���je�n�p�����eq��g �"���6�C���=���-�l��k�p��iu��'ft?\�)<j�Gk鸢�󋒬zg!�,*_/|��oW�N{��3�	�6Dp�
/pƀf�A�$Ⱦ:��89���@6�@@�)_�~A���t>aZ���o��	��#�5;���d�2�:ϵ���ɕ���Ya]�7���y�� ~9�`����,�u1�{,�����HR��:�������F�Q^�Ϩ>��h���❒\4+q)+k��+��qNiH�z��$��p�':+�3/�1�k?7�5k+��Rc��7�HVZ@iv:T���u��sa�I���8&�ү1�W��,w����Ê������>��
�DŁ�dޗц��/,����\�D4���Y,OO��J��y�\����͚L�]ۑ̚+j�?��|(�ϦX�Tq�)�������@v�/=(�2@��wG{)��^R{R��j�69Q\D�d�{ܵ��8�yh�&{$f���3փ��0�N�8��^VC��a.����|6��u�}\�Wܛ���5�V��+�����U1�~���۷ܜ��
