��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]�1ҩ�r#��9���������ƍ[��h����%�N�
T��M�T���'��ZR��o�v��I���A��?!j`�ـ/�u�"���~�R��j�ژ4��1�+Kz���,%���1���-I�fA�;`������_U,��cm�7n J^fb`���m�>|�=:��fB07��W`T:��b��'R;�t)�� ��z�ܟ%�(�׉�Z��F_�r���<��n�,=ƫ�#:$�V�X�v&7�-��<�rI�g�+Y��~a@�ޞ����Iu�ǽ�Z3t=�_�0��]f|?|7|C ��2Vzć@���꿬�K����a�lN(6�P��p���qF��\���!´�3�t��K���Ba�Ӣ7ـ�����,>�I&x��o�
�-�+�~�G;������C�^�.x��OND�S�lJ��W���ks��e&C��`�#9\Yј^���T0WJ�p��%|p�
�1R������U�-�.{�1��\�ڤ��ߐ�m^U�Ը�
;I��W��^���5˿E3{��8O:����:�8����}S�����S_�n�\��$��IJkc�Ҕ
������oV�$z5E=8��.�����zT�WX^j�>����X�H0���#���	\���R('��E�V�YVVv_����P�5l(rB���i9O����*���.#l.I�R�l�I����7OT.�~td<��;[?T,�=̀l���t�f������Ԩ����8��>H�����/hbQ~o��������LԽ}T�9�� ���x�Hh3 ���n��#�,���P�mv�l�-�WU�ř�>B����
~G��r����˙1��O���B�J[\��	�f�P����{	��d����G5*�/������ڈ�V���a���7��i@�h����F�+����Prv���Q�(�����.���2�J����g��!_/Ě��Y�6O�E-2�􄕲)�9]Pc�ݫdg����7���>J�A�b��x~k�l�R�Z�����}���S:�z|e��ܼ-���Seìj��:L���f�DB�r�@#�-:�֒�@MK�@���b�R���Z�'5h��
�e�J�G4=(����{�^]�q�H�r�F	���?Bb\��B�OY�Y��j0J��'%Тnm�D�����F��}�����ԁx�܊��9yw��Q�������$�#_(�������I�����=�/^�"l�HT���L�}�]���Aa겶|Z��GzAq��f��DV��uH��[Jݿ�U�2I���1_}N��;�[�g$��M��]��x �]�S�BҔ����*�:�s���!���\��U���n$�e�ӉQ6(��)�ɧ�U��bZ�n#�壅�H,BC�&���x�Ϻ:1���`��	��{_�Yފ�;�m9��>&`���d�_>9��[����O�q�_F̏c¶�5�o�}�
Xn͔�6:^#り��(s$���>�i�}�-X�6�mdk�:[��4��Q�W�p�Y�o�]��R^Uj+�/�]p6+���ٮ,��A��7���3��X�ĚI�����~Fk8E=`�xB�C�'���+����J8���>TQ&F�P	�(�t��^7�h	l/��,��p9�����ʚ0l�K<��=�UE�?^�>�����\�8<U���ڏ� �T��d%��E\��I��j�з��esڥȩ(y��!�O<�2���Ӝ{��=q�+��x�������ل�EO�{�)��F�����s���؛���Zvj&�k��<ȭ���H�ʸ�Vu�H�_����?����P\��sY|ɂ�zL�TeHS����CJ͕9Sz�F5�q�|b���37�e� �����aI����!�����:G��cr��ڡ;���W��̘S�ݚ�|�9x��ІBd�GYzJhs��N
�:�s��r�
G�6>A����؆7j*�3�r�F�Z?"�=�-q� r���^���{�o�E�����?��ر�o��5��'W�KC���[�$�Z'�6T�\���b?n�z\��f�"�Z�Ql�!�Pxĕq�DnS^�U�9	G�LOl�۔�Ń ���Ղ��GZO��ͯ�/տ�n퍚�=3�iʅ��3P��|k������;�Ooo�;n�V�ZeFS�����'""��� -���"~����D&�����+�	ʂ�|;����U��)��9K��g�UNGj7��\�=NU	ӈL'^��)���B����)��ы*i��,�X�S+8���	z���G�0nFI�`X��I��e�G�������,����,��.���KzQ���/��[75<��# I��J�?׿�@f^���5��㰖�� ���6�L�mf��>t��G��b�����*9'2�����n+[F9#,�Щ(��b(r�f����1�A�5,�S���v7j��	���c����[�:$�{�=`�W�F����s)���SŰ)ړ0���6f�_���+	u�uO�n�H-�[$�]^Ȋk����B(Q�C ���d	ہс9�l�o�a���������Vg�"��&|	 ���/{ݣ����ƛ��9x�(dB�4��j��m<e�mҾ�8�S
�^6R��Jp����4W#��Y����h
��P�O����)�D�YC���Z:�5�%'���iF�s��i�����G�Y
x�0M�a�E�v��4��ta`��p�C<��}�~���tz�h%=~���2&��~��(7��
J���G��>[�GH^5y��L�ރ�gzkO�7����I�Z���n|��<�oΟ)ȳ�տၦ��-|���b3�5�c��(�QFG�C�Bnߨ����
X��2��pN�ք.O����Y�Kx�:��)��Zǳn2�����ѻz�H�V��Pd�%���;F~��~�������<&�&�J���c��c;�!��:�Okb�V��DUR �ۏ߆���e�����Ln�V�%1���in/ĲG����n�k��iK�L�hwj&�tK{�� �� ����Ì}�~�1*��e���u~Fo���xm"A�-w��zlEp�{��^����J�����8a|����RZ0�T���0�
���Br�&F=/AM��['�n�6�9=�E�
��oG,�u�A"��m�M:�1E®�@"��l=$}Y������P��Gf=ii��}HXb�p�A�'r���&�Cɩ��ʟ^{�]�]��6 :���1���E��~p�8H���L_���z�a��b�8�OZ����7� �	H�tMpg$#�J��ñ+���S.&|�=���	�}��=[ q��&>�U&�9��mO������摝�?�⹍���6U<�&�)����ߔ�:�o�`�\uO�����/" ���*Ed��r ��h���o�`l�.��?�B,3n���1-l��%g�䣘v�i�����ᡲ��-άaf����d��Z/�� ����n(,�P�Sӷ���ѷ��x�2O�׹���4�Ug7��D�S��BV"���?e��GJ��T!��弢5�s�4�g���*$gG�*�8R��XjvQ'_x��J�z������Ҥ%I��o���Ə�rd@�����ܓ�e��w�/ ����>��z�vTq&jLΩ���]W�PZ����������j`���n�W��&�I�ԢG��^kP�Ο���e��4%Ӂ�3y�O�"���<�	;�n ^X`���4�Kh�iF���}���M>�M�˒���a1�Yp�g��2`�r��މ���̍��j/�,I;@P9qԠ2��m��j�����L�'��<��;�6�8R�=��3���bb[�כ� c�C��>���*�n]�����Ę*p%��H��o{���6.������x�#Ïo����G����em�z(U��?Z�hNL���R�F�m�Af��g�e����4��	a��r{�!��~��=Lv浙�7���/��q���|��L@d�݈�SA�����_�}�E�-��j]�Qa�,��2s�vg-�
mUd����.,6��٠��0��ujkJqQ+�{��k��#�9��D"1��̟,zSY/�EuE��Q��˒&$䂤�=��9p�d(a��-�5����5>dO0GZ�iA"e��G�+̊��Df<u�������M��w�!i�
ۈ����Wr�_�-�B�i}�m>�����\��d*��vv���6�����hJ|�h9�Ȩ�fW.E�K�wdE�����/;U+�ywi��da�$��t�&���
�X/�2�^DZ�!�υ^s��H5 �9G5g1�f�;�N7g��k���B���o͍��81#|(:*n�o��j
K i�i`Ks�9��&ꄯ<�oIX=3��C� ��a����t�9H8QY�#4}a����ê���6�Bb����L�#����K�/r-�.��Ƿ+�W���2���B芎(_�8�1�6h3mȝ稜>�k��b�����!Z;t���2VmG#�<�����Vw]s��&X ��s\ve�G+�W��1hF3����"��+�{p�j�đ��Wů3��&<�~Z����S�j�\�`���}��0�4�S�5�[d=Ab�L�%G�����
.2��g��
#�n��\S(.#�4�N�˒�膗��j�U�v�> ��lp>مMPZU�G	�	�j���J��_�2�`����&�i5?�z��k�"������#���EE:�͵�]G��|��mdJ{v/�����x�==�Z�������Гg�P��˯1������9򸵻� �[R�;_�Ė;,��Iٙj���5o��.��__{����f��ݱ~r?��� �#mt|��^Ӷ+�@G����l�Pl��ᚨ�c�K8�eĖ����g��ژ6`�����V)���Zt㭀1���H4���Xz�Gf2��,b��!w��*�#��/h��(�FŸ�c�~�]��N;N�'�դے���L��p��M	[�L£g�Rn1~~���a��r��T0)4����4�4nȟ
�K�����ф�~$4�3;ZK
'�1�$��X?����4Y#��gq�e�fU���6F�R"%�U�%=Yx�gKjQK <JV���3���P���~/I#�T=;T���g��4y<�5�䅱�Iq�-9Iq]�4�6$'�5��#�ꡄ�T���䘻���(�P�����L�1Y	�hMxzȅ#6��
�8tHf�vԵn�VG��ȆC��
�Wo��Q����ѥW�GM~�U�P�d[�9{P���v���
Ы�'RԜPĦ$l�;�a�C|��ΐ�o��↤�8�,.�mm��-�Uo��8l$�w����\4��F�����ƐT�B������_������{�&�v���"�o�"G«�������lX%+�?�7q�,WUR�j�g��RXJ�8\{��W�}�,�Έ�
�б�_���\/J����%j�t�lY����š���$����`����N-���E#
0ԤI[;��2�NH1�}Q�X6�<3��7~��5�٥�z&(�[����~���پ�Aη�L��J=