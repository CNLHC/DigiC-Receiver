��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o��s4��<�	�ʡ
ISE�ᭀW�]ǀ�h�a�Bc1��D�_Be�mP�jH_E����9NU�����TC]1o^�����N�	�$��U�(H~3ܺ-tϋ�q��&��ݝ���o��d�~�{o'7�t_;���:)ل�l�%��S���"�B�(��.��������px���5��a�՘�c���֭�푽��Pd"�E��Su)��Fn�>'q��c��T���<c=:Aj f�Y��M�gl��"ߪ�ڿ�I﷭Z�*|����nȮ��i₢8�z���[�r���D��D�MR.�Z��^*�+}�.0�<_�� [-��.K�<-�EL?P4aKSX�,��s�J�[�^�@'I������:�����W��T'7�:��2�nXJP���^�r� I�czP�'�@}��R���YA=|w^�(���tH|����s]����L���(�LuGX�9n-��a$������t4���?+��ܬ3���l�(�ז��	pa9v|C������{����J��a�36��9�62��,�lPi������y�Afs��L���RO�
�"��T����|�KDH�����k�2n&�|B;�4�JǢ���lZ���"e�T����w�g	�[mf�#�#I�Y��=�y���7R������E�tE��g���*��I5eQ����cIp����F�؟``R̀Wa�6��`|��B��
@|b����%���p�4A�ŪJƤ:s�@���D��4�9�j�Fm�FdyNG^�80_Z��٫�xW�¥�#�c�q!��̯qQ��w4�SƎ�꺏`���"O�X��rP�Z�c 3�F�|�����R�s��z��{�̕����,����&����O���r�d����&�������_�3�*o�j8�!��-�E8ٜvg�?|\})ŧ��]5H+��B�/:w}�D�b����'���[<���P>�H{�:o�cA>.
]�|���n��f��+��~�M������0d��\�q��[%����Ȧ��6t=�lX��#��z&c�����7����s�Q*��J!������2�?2��=�VR�@�b+$:�~� 0��S�w�b�:�%�Xb��V�;��ky��~4���g0&��K�>�������x҂`n�o_�-H)��%$7��%��Xⓓ�q��}�d�mV�_��6͵(�]�������n�t��D��P[�B�qZ��G�����wR���UwvW���1=�B�˂/Q��(c#�k�z�����;�5uDh�y�b������%�]��vzj\�C2J��b����AE����ּ�Э��Y1+_o�;�T���ã~��V�!`y��j�����v?P��=<i�n�����}\�s����@�ŧ�|kx�_\�?I5����P�g��D��8ul'��U������mXO�26��q]:�Vn]b��-F�#�v�a��1�h��0�iH*l��0=���m��nx���R*`�!3x��~|��T$v�teI1l��V5u(����
�ϜMd��cYG�j��kv��'�ewD�;��7�z�A���#�p�sJ�H֨��bSX8�E&�Ta�cz�I�O����U�� ¨��*���m@���麝�a���'��
���#�eC�'�b��=�(w���q#.t�X�m�Ļ��;]�wBk&aoLwf �nio^��g<�ax(��0w���ں�s8_R8e���,Fk:j�a
��p�v��m�M�>q֜����q}�i����XO��%��̐��M��-���-������[yPL�yH'�r��9�2Ӟ�m=��Œ����	�3����Km� C�b���d��4U<=MtY���oZQz&]_R��)��UO��E�RK>��h8�P+B[9��2�g$fU�?`�&��4�h58���9��^�_��O�"���
x۹?�X��3`�ΠeU��b���0�y�~�TS:���M�Dlf{��q]#���� �ח����[�E��?�e� �j�R*O���7<���ߢ�_�7�mQn�0����Lx�hQ��xr��H�y<I5��I�*+BI�~Uϐ�O{V^o��R����@_��e�Ux�����\��	�A��_U�p���1۾ XI��ש�"F��B1��2F�h���٬������G���駾�Mj<	ʓp���-�Q�9gH��jf�C�`Q
	��J���<7-�IN��������zO:�m!&$g[6�^ ��lL
�/�$a%�.<�A���$-��Qf�ޘZ:���@"|�)��N��Ƞ+�������y��µ[��-+�a��Ε�Ȝ�f&��F� ��8ui�\��ܻ��x���� l��2l����H�T�L<���B��gc׸�M.�>��)�/��
D��B� �$����r�j
z^uWC31����(��$7`�XA$���gHiC�+O�t�����V���&`*�9���db�g�\d⪖f�.A��l��CoݭK ��@U'�nn�O�G"�>j鮝�We���, ����WiQ<�:��n\[	IE"�v�<Jn�_y-Pb�~�t|�!t��Skg���#�j���|���y�-�\F%�	*"�饨�o�3�˾�^=Z9�(`�8P�<3Y@�ZZ�*���L!�I�HK3o����í1�x)|A�o�T� 	:���R=-�B�B��4��o����o]�7�1+x�I�N��ko���Hh�w����mʴPHP�:�u��H��!��!ӷ���CCP�;�vc�jT�P�u=�S��'�^(����=�����$�E�3�	륈���|[�1��	�=m���e�iy�k��J��BP!fP1G�f�tu���D��8�ϋ���,w�L"���Υ�	��\��NǢO8��h��h:����o���{�z~�y�k}��M'�Jo�=5�>s����@Ԯ��.� /KqN_K��_�4;9�m��Vtmu�[��M#)r'ih �B}�L4@��[�Ɗ�^�Y�UU.�� ��I��C�,��45���|p ;�ꓒy�����9��g���nқ��s��>� bz���!�hI����oj�b}�#��I;	�Xmt�ӽk+��A��<J[G�����ϫ�{=m����I(�G���QS��(EH�IU��GzV����Ep8{ڬ�g�C��g�/Eۤˉj���0�W}z�"��1�\p��~����>� Ba8P:h������#6\����Uٷ�z^`� 'T�xF�YG�4-Ȃ	8Q�~E�&�Ba�l��;{�y��'�ZE(]�&"^UL�ڟwN�ǮO9����|��T_�CO�F�Mn�9�T��Wʀ�uJ�|�(�z���l�������$^��Y�me�ѫ�-�X@�/�1�tJxRY�h�]�ڤ{�w)�z���up����
a���[`K�J`��R!pbaE>f.�Bx�.��=PL�@!�:���Yk֮|j�
�
|ƨ&�y�� U��P�˛ ��8��-��Z �w��ҍeR��;ĵB��>P֗���Phk�3Ӕ،+�/�	�����ȅ~$�o��k��lP;��9�?k�������UT�K�W]UB��b#ۥ_(H�c�/���(~��!�k�-:�3g3l�4$+�T�S�D�gT����Gf��¢�-��Ro�TaÞ��'�>�o�@�ۋX�\����#��S�\��ބ̟�9Y7�靺?��T�ԡ. e`N�tn����Z��b��OK�0�"�d�<.��Q>�Ԥƹ�P_f$8
k蟱I���}�,��͐�O܃x�h��#P]W`9K�\5���c�]��,i=y>2u��!H��>�5��M)�!��$>t��WR^`{U����d�!pk�#������:| pӈ��*�,�{%��X�������kJ#W�-�K&Ò7����Q�j��z��K��p�=�񸳐߬~1Y����伳`k!Y�xv�7��C|n~c&�e���b_r�4?��RT���`j�Q����J��U�q�ߒ�|0��gO�oM%��UP�M+R\�W�%"����&�JS�ʏ"��� �RU1�5��"�B�B���,�BA�w�u�`�ȅ�[K��+v��&�]I���ٳ\*�,c��f���帚&�u�'ؚ��sv[��������߿Lg)Ez񮄿���K��+;1�[���V>�#�G�!T������jU��zU��U֋?\�a�A+
�iO���on��=y:�L�䯊�M���@���$��>��G��A���|Ϻ:�j���	o���j��au���YĒ�u�L�r���?����ϳ�Cs���T&�f��h��)��y�]'���,Me'�D�REB��hS4�#��'`=�� �L|��=J)QGh�P��b����Ӱ#�x�f��j�/ZT�฼4�����@�4p�B��%��y�4���`�E{P�N5c[��O�OK�6�����C����Us�k@��T�C�������kok�R+�Nz�~���\����=|�;�#�M?�u�����&K����k�5�磌0Tn�O �3G����0�@
{����� !mF�6���ٗ�wd��B����	��Xϑ�ջMY�<&��R\`G��d�jQ�W��nl˿<����L�ʂ���ר�[b�M�
��z�M��.m��d���Hs*(��L-��]"Os{>���6������Bb��b�!?y�;B�+�9N	R�	t����R��~��u}�R-�#ɴX ���;n]n
��8EImRsv���D������֕(��=b��Ew���������[�O�,�|�0f:,�#�z���f�S��u�2�ڸ=����h�9�"����q��(z�a�%tC������|�X/u�Λ}h�S��;h�8aM�R� ~�����=3��e L�KsseI����\T���$�H���4��Lζ���>�M#� f"4��h`ơ[Y�}����ԓ'�x:���Ӓ���bW�5\ú��}k*��4ɪ������3P4�!���d���aQ�r������+%�O8�Øzӭ|=����})�����6��?�#� �2�0! ����}���-������ɟEV��B�s�Bu������EV��c�D��J/����ZB��zM5������\��x.N�U��ͼH���S��~�wuE�9H���
�RoLD���@��Oiؿ���sU�9�G��Oc��}��]�	r�҅�����J�,��lJ�������Yj��QE�Ƨ������ܹ�D[���t��i��Y����"� t��\�u�f�2�������r��K+e�ۖ���2k�b��@�APP}.;�V�F_p[	��dꚙ.b\�?�e���^�LH s��P�"����������)�=2\�.��߭q�c��q�cEb'���$�x�i�����x�3�01��֡`9����㢏������-��F��֨���7JV[����&TB@x�?".z�c[C�6���@�g
��!���˕�Ck����qg�]��*�M���wt�ڇ�������>gՋ���Z� ��)U���@%"� �!&(�\��j���8�*��8�.��!��{Ń�^d�!˂@�ۦJ�X�c��F}GH��ϥ֡�6�$�j��G"��#J�m��q�k�sb>>��6ih��ƽ�v�ʹZ`*:�N�P���΅�<B���J,w76����Pj�z���hD�ʿ`�02�k�S���Nҥ`���~{1�`����K�.�������ڍߣ�)���= 2'��Ӵޢ( �

�ssr�Ի*�`vg�����VS?6ݺ��sS��Y}����w�!�ӫ{'�q��������&m��d���`℟�*�2}a+&P�|�����v8�O�з/P^*9�C�^/շ}�cJie������Se�S�D�	'���*�<^O0~�ɡ5NZl��xj���=joa%�_��zLuP���_��*���`�Z���:�sK[���UI�����)��G��ۜQ{��[���g#l�w��a��l�6��!���D5����;t�Sd~�����f���#����&���ov�58P�� d~mx52�EkN?L�[!�#��G ���}���L�1 ��1���fla<��|�B49	���)���M��e�|�g�)�	���U`���^6�=I����+�E�N��m3U�|�k.�p����=�iǽ�X�,�A:2*�y�Z���3��:�����o�tu��:��ɔ$y�3y��Ⱥ"����UcĂ�Ex4�$��aNjL��f�eO�݂㛂��¬U�uA��C�tQM�J�������g�G8��,�[]��Ԛc��;E�}ų�f$���}��a%iЊ�[���n����Oˑ����L��]�K3�#�)0�(Qs1@��@����#�l@.�L��x��y`���|^S��h���F�|v��n������,X�4Q�j�f���N1`�/��q�Y�n0^�"�~wX�F����ќz��.�X�S!��R�����,�=���Ff��t
=n��-���2���W��x��+^��?�%����i�A�^4�:n���'�d���{,�q��Aj`R��q������5�2ks�gv��Gʽ�Z)�S�d�8|7ڣ�Sa[\��=��a ��^��f(��	�T���Zc��8qy���T��P'݀#�=�BDK1�`xT�7����	�l��s�b}ݬ]�Ak1��J�|����8*Q_�&�K^�x��X��ypP��T�Q�7n��Bz�P�Q�r��>��>,n�;���$h�1�����0t@\�������] �k�g?���T��S�a<��)�R�5<ĭ�Bu�/�״��b�]���#X�y&S�5���+��D
f����;"1=���g$�^������g8q����$rZuKÙ�����l%I�ė��\"�G,���;ˑ�ղ��pf���|KGz�NG7��i�N*#m/3c����A].%4��l��|�,�IZ�����Ta�J�hP��PGދ@�j�����ڿѤrJ����ѳ���=�N�%{D�=d^���v�T��uC�r;�b6�������Qp��'���5F��?ǭoh����#T�C������<�D�F�rc��6$̐#l�q�X�*P@suv>�9� �����������(���n��ơ~�H��� �^�W���n��j��Yp�q�O�:�=��C%�h�X����KBC7�q��n�{�m��'�̸�ݖ_挤;����]`�}rx�|�1�� y�ޢ�-�O���f^�,�Dd�B�1�K��H	π1���gsf��H��G���Ua�q���H�:�~]�����L�H�@�i�,Ʀ��������, ��M�q�d.$�����R�\Ce����v���狒��p���=K�W_kU��<Uqդ�:��AV"�$���7+b����<T�2�fg��R9pbWհ�d�n����:��`֊ݤ"��/��؄s��$Р��p0~a����䴳���{�o��[0��*�XQn�n �3�h��QP��%��M5�oQ,��*r^q_#2�]t1è"l�ǌ�D�`g������؆޲O���@�A�xp�Wdٌi-Vq�ç�$f/bv��B�9)?����ԁ1��I�겴���Ƹ䐉���N6u\Ј��^�[,�����y5���I8��c3�p~)�F��7� R��X�򨋈��x+��erL!�%K��˹?�d
�p��Cj���p�V�L�=���/��T���OܚBk�AQ�`�����!������C��ξ��I1�ԫZ�j�F�|}G�`'�Q9"�m��q?�H��SM�֤XA��t���&��,��G`_Y���N�ǀ�Q�� XN����U'��I��X#����΁I�����e!��2�s�L3�����z�y*>�d��1�*����ZP'�٭��B@�=�XZ�t��~h9�؇<f%�H��qV노����űe�D�5��F�Չmx+��;SFs��?�G7/��Ҹ�.֯��+��9����$HYޔ\�e�e%t#y�{�Y�Q��,�K����`MU���k�*��B���
� ���ѻ:�@ ğLU^�p"�Գ�K9���j�2c^CN��g�4wMއ�D���� �����k��E� �s��oUQ���P� ҳ����Q!ji��2l�z�+�����(�Ye�=�|�,�w�#C'�v�ٮ�K�K����u֖�t�g�]�9O�3�l�M����6ya��_JI.���j N����7�:jI�B��߈�-CY�s���t��" tx���H�S[#��9I��J\�}��9����N���g8��Vv��v<���)0�����BR%���D�O=LL�F����Ïʫ,(�(�r�������hub�w�K��J�V�C�"]J�9j�@�;�ELX:�`+�$���r=x�ލѤ�LX�5w���^�`�!�A�����zo!�X��V���	B�	��k]_�4oɁ'~� ��(���I���n� ��V����o���a�RH�_͞�9Uj�kZ�2�zxG���
Y[�͡Qj��Ƽ�*���rބ�V�����zy��Dw�� i��"DC����]u7"@�h�Mr�g��/��<�z2y��\d�∎޾�m��s�d�������3`�+�K�;� ��k5�wa4Qi�8j������ܠp2��vА�(\��. ��|Y(��Hw)�1g�J�s�.sE����*�/�^ź��+�����i�b��Oւ���0�i����M-%m�3����U[�x�c��(/s��ҝ�`�۫�>bB���_��f�X��Z�W�X��_QT��6��UV��	��J;kv��*�x�pEs���SA��M�M��g��D4����~�1�� �^�$�+�ԉ�30!������;��7�;�6��t���G����l�B�1�M��M/�E9�{-s�pl�D8r�>���7M� ��Z{��Z��:K�G���o�#tX(�l���
��6�HY��ۂ򏝪L����3,������RLsf>3�r*���B�X�����������@��2��Kk{\��qN�y������^�U�&�ۅcɄU����(�ø鉡�<��).�`���AQD�q�L,5�&}�!�G2
@�}�,���E(�P��Z �[b"�@H92L�^�r�@ ����(��R� �c�4���M`/ĬnFH�ɣE��*�
�K�;����5���j#�qR3�q�3�����|l��eQ��� ޣ��h�8t���A��͑Cډ$�����z0q��|]W����� ��^����h��Ϟ������d63P�H���$�mt���辝y��$�{�$�zC�(�V_㴸���8��?.ay>"�}�R��{'��f*'g���pVyZ�\IElY���F���\쥒�@Ok�N.�b貱˭�L�bt�`�ϓF��u���O\���l�`l����6��&ym-sz�%.݌=�Bq��b�z���6߾ �v_NV8�o���)���q�I~��j���{_Uw�(p\w���J��m%x�p�͜�T���V�h���Y�;�H�'�]����Pqs�ss:�4��^�����	���3��B����A�]1\�������O�l����I64m4%Iq
y��s��2��1%V�0���`�i=�=�����[��z���#�_�t�o��K!)ˍ�'�Ucv�(�3[*WW[OV~�C�.�=�{w��
