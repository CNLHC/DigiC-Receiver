��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���į�?d�tU�0Ѡ\}��XC��X���@hš���}�:�b��ֈ
CvĜ���T~�%�FXhgP�T�2㫅\��33������&ꬾ{)뫍��@��V4����riY%����L����֣�p�'g��ٛ�s3�t� M�W7�u��HDa�����8�"�w:��&eg�(�>�T}��X �bV���+tN�G���nl�,$��7�5���M=�w�*���s����<��jb����)��v�$��(��$��"6�°�3�,%�>���N��6�a��{1)�	�?�Gg����ެ���J�ol����M�\O��(d�4�)/A}�-iŒ���F^^��g���~���m@�&����F�ꛜ3kc?k8���X��&� ��`hzx�Zt:r֨0c���!N��:�u>4?w/�Ӯt����y�%�������D�kT�\�053�w[�)�����\�S���SD�VIS�A,�����:���kw��O�i�r.�]w�pz���{;щY��]�0���H����:84#�H�/�G�XM#�N*��kOy�.� R�B�����LD�E2�䓹&fĩ0��69G�6�jeCn���Ǒo�C/u(�<t�7�;��S� ue��e8�ϲ���ԼU+�9m�+H��Q�S�\�F��l3-��K�@v�S^�RpD�V����a���/�������"M��o_h(������cP�[`k-��1��[e�4��Z�����4�F�{%Z�s�@krv
P'���]����WO�w�߰	���W�w�/hC��YX����Cr��my<���8Ζ��wȯ&��˸͔��M{�60=r��M\����#b'��7�ė�F�V1Q}��i������w�9�V�OcF%��G�_ @z��"%/�,L$+I��	�g�R�"���P;��R8� ��^4���aj<�u�O���pdU��X���}���1�%��a1�2 *��	ݔ���OP��[���P��Iͯ�QVM�o��6mJR�,��@͗j�j�.��1���8��2�f}�O��CQ��4n�	�����FL_�!W�
�&��gN(��(�7^^�M6f%4>�����|��B,�m
}�E�����?�i�^K���JX�/��Q��5���bS���jU��q-��`eF�S�7�#jsd߾s �#j����xm�A��k,oʢ9��K��_ph��&q��\�#ը:)e��)3�L���x/���*}�8����J���I��Q��p�U{�ʨ��M�}4t����	\��1���1���>/n���Z��K��h���{x���E�P�D�\�hu@K��d~��*�(����� �[����dJ�tRB���*ۓ�Y�R�`Fa#���U�w]�p*$��/�Ő�i�px'V|���95�Z��H��s�@ �9�gM��Wgb`��HD�X3/�b�763�@��r���Z��_��al�*�]3�� �)9��S��e�,���S�
��$h�w��˛�)���7�C��wh�Y�N&R��L�l��xQ�ݔ�tlS��t#���:�l	0"	��z𓑗s��2� �x��n͙p�8{�}�e�zy;�� �U6�x<�_����VXE�����Ұ�xި��tbIW�����'g������7�p����N�/T-�S�P�KQ<��e��=b���۬�L����nɒ[&�[u�B�7���#�P/��`{v��ƅ����s��U:;�2����_<5h��������F���҂U��>ɩH�2��]Z��/AG�Bt$N���<��vZ�wl+����i�׶N�7Sk��{O����w��^�ɃׅF��H~���&�A�A6����u#!RAd9&,��c�f0<�QF�{3�b�s�D�,=�佇D(L��,�xf�rA�O���{p�*����.g:�OAf3q6{�tqb
y��e�R��X��a���F�.f�&kr���Z;�E��_�s��d/�> �-�g�%��N�A�ZH4�dLZ�f_��kF{6��i��Y�.#e��@�c�v�o��z��0��{-��d�,C� U)�II~�(\��JP}=�*t$GZ";�Ϳ�C���&�b���2�$�ƭ�}��ga�YÕ)��������|&�&L����w�\�)5QXc�p�mūq��Z����:Y�t�1w\NH[�����Xڴ6���w(3汑��dok%B��*c���"��p�������q��$%���(��r����ZiU[����vڡ9ek���X���r6s`ٻfѴ��y�׫x���_��M������Y����J���+8&,�0�����>J�&�i�=N�:Gl��k����``_wc([!���b��b�<W8	�'�v������_ó.�"k�$r�n�y�pyF��ǲ	�(�tu=F�_{"aNC1ȏ�'D�
ՙ�K����pL�Vͧ]i���YHK5F�H������5D>Y��kVb����lbY��*I�|���-�&\�N��c&�s�"�)�_��L��B�p{��g�õi�'��%X�Q����G��pQ7��� l�qd��Uگ�SD�i�	>��ڰ����j4�!�Ѩ2��l��ܔ�Aq�"�J���|����C~�8��]�
�q*g1�"�{�������FT
�G�#*�5���Y�h9ď�3k����L!��|n١���fɌ�2%#�SQ8W��k�)�'��"ٕc��۪�Lv!�/{>�~u�l�C�%���i�M	'�HT[���=ɒF+�b��o�\e K�у-����6!d瑕6V��v�U��B�31����3��w[�a��P�v2�	Q�:�XP����$̉'�l���+C��7;������Zz��o��k��y���:�@ �2I�,��_߸qj�n��ѡ��T�۳����u{���t�#�C�����!�2��<�Cf�B���R�"���n�����ɛT��?M�A�95���L����=g���!�K���vaS�e����|��~�@h��WS<��b�M�.�	4��G�e�]���K^2�RS3�R(�3|��*�/ʳ���h�&�f=�2��� ��p�EX��I�o	�w�C�Iz��P�����Nq�ѫ&4���IZ�Z�%��Me�Q!:jb@{�Aс�~\K�/�ǩ��N��{>ġ� *�yӌ���qE+bw�=�6j.G��h�^x�wQ� )[O�դ���;)�rf�<:�n��߀:���!����y����B�u��/c�zu�39 K.A�to{�?NMW��6b8��U�4𙰒�J셁��D1��I!U�k��8ME9V_��b۟S:��Ӣy{Zc{��ui��h��_ٗ��]l�/"�� ^^Ec�V����_~�C��ߖ5R=��ς7�	�;��̞������X��}�}q�W���W�ĸ��'���z�~y���yM@}�囓)�v�0%��$Oaq6AЪ�?؊7=�Ӗ���o�-Y�ؿ}��}�����˴���F�w`���6����Gv�����W�V�8�߳�VH4����܌�p
+l� �=6(�j�R�y|�/x=��}̿� �o��L�I�f�!�]+g���(�M��\�z���6��t�x��s�9�Z�g�db<%6R:/J�߷����-^�Nq8<�u�,�,K��j�o!cj~��xGu��2܊+o~b$�1O�7 ǌ<+�˟
��V��f�/�F�p���A�#��r�|�q$�ZXJ��%�I�qw���ܐr���)��f�y��%(�Ol%w�t��ڟ�I9?AJ���:9�����Cwt�����=��8��Jd��̠�zJ���s)m��K�3s	xw���[v=�NO��)O��F�c�.H���V��)�hf�K�#���Z�Ê�lh!��9�zOQ��uH��ķ-xQET̴f�l����-޿l�٭S�b���
�#S�����o�{$!���.o��g�ϓ���&�{F��]v�C��6������%6B�//'A��d�R��"��v�{?�f��6�.#0�sS�oteS� �$ �a����jO�B�]����؊�a﵊��n�俎?���+b�^�492�����^�)jt3�W���-����{��vt�L�g�[߶���h�fU��F�^hU�l�)�=<�Y�/R�1XT\�ahG��qk}̸F�<z��������&��{�rPn�g��ɝ4�T�M���j׀u�5� s���E$���^�TüI�}R%��'R_�w�7$����Ƽ0{�\{8SBv�fv!kJ-�� ]��ݜR�A�da��|aK~��q	���|�au���!m�gy<��<���s{>�i�.�2���	Ն�����(j�Y�/0��O��Gf�"O����.j/��&��>��C �1g+�D�oI���e�4z�5c�$;m$��LOTmH�������jPM\������� �4ܖy��W����C^{",�j�d���r�׶[m`�/��g�KS��:u��+�v|�~��^`��q�_z�����(W������d�C�1�?�� ���7�R�Z�4�x=�>������U������c��o��[��HdO��{���a��`���!Bi�c"�uU�j0hL���?i��(�������{��5��6Q��@�<V�'3�A���f��n�o>*2�E}��V{l��fw��L?*���vs|j��m.T_��|چ�����7��Nwh�ݠ.Cۤ$2��&�P��j0G�kMz�u��S�z)"���v-���^�-/^��0q���B��PalTĠ.>�����k=�*�	���s�zg�^_0� ���{(�P�B���,��[(s�+���z[�z���~l�*�/w=_F��{مP�����/G_��P����.��{�ҷa�e����i#@�D�����Dv$H���+T��3* {�PkD��^�pl�� Z��S�)6�[�Xq1���d�rYV���;�U�^���-�~�&�9{O�)D�W���ab��LǢקA?aR/y�`y�J:�I���m���׫{#�M�����1@��Cy��N�Vx�*�ʒ����y[n�BV���r8���GX9�ߢ�"w�e�Te��ʀ�F���>� �?Q�Ӭ �� G�ꛊ��r!�/+�Q��|s�.B$�坵��<|nd��b�|��`�T�U���N'�~��W����O	���2�&?_������pG�+�a��Y��g����ìO����Q�)M'��H���A�a��V����A���槆�M�3)\��D��a�c��B�X¨z�� ��hK)�D9 �S���/L�B;���{IȘ�2�I�	N��~��s~�*����G{dX�L��q�,V���k�du04o�N4C�G*��?-�|�4	t!:)Z�w��w�|
��P�]{�ߡ`���������k:��5���"@�o�.c�TIv�xֶ}�^5i샏<Nƍ��8�2�cu&��4�惁�����T���Gn�q�y��ŕ3ú���i����ǐ��g�𥎯�]�¢zm߷�K��`�\y݋=у�|�M�&��5{�:0�,{D�)J��_��k��C^m�Q�zݵ�C�XU=_A�� d��2S1Z�.��օ^V�ۍ랖`�K&c��E��ۂ|��=Ϧ���̨��.a�{.�'��WH��Q5W�#y�C)�����pe�����iw������v�D�11 �mu�fV΃=D"�}�E�|qò��Cݕ�6�b�%6�{?�#xVA<9�*���RՏ!��s�������^�d�u\�����`"M	�52p{y4��H��=U�*;X�~ó��^�'!}%<�q��qBm��D��u9�$i��h�I���c����ʡY�M=���\��;�R�Bl�I�EM#�|�l4g��`L�q�Y�O��/K�षt�%�
3�������.~GL�y!8��{�es�j��>��[K+G�%=�W/�c�WgV�=���e���X�8�Hĩ ���	�XZf6$>R�X��z���"�{X`�T;�+,7F+�ڐht�k;�ظU.ȕ1�
 �B����#��'���8�@��lݝ'\k�cumȂ���ftO��=y#vd�h�_5�����Q�����Ւ�k�D�����Q�~�K���7�������G��4�2�<���K����?B�Gn�%��Y�׋z��/�������bb�j�0��f^_ b͎�fFEN���m MT5^QM�>m�v~�$�G*osd�|}ے��=(�����`������@�}�y-���}5��(s��$��bO�S𱴱<,>�L���I���Ӱ�G�m����Mҙ'�2�-�+]+M���'m�V'��x2'��ك��ϸJn�k�Zߦ��*vS��\M.k�/�P��g�x���G����-�Ā\���l��?��W���x�+$e"j.�Y�K�Tc���,�fn%�"~��Ȣ��):k۠�zL������jm���|�CLV,�]�բ�!Z��ra�=��@�&�SKM���ZR�M�a:(�x-�׆>A_�c��]�,tKK	I�܍]�=�*���a��Ĵ`�y��7+x������K��[U�$L6�����N��M�T��%��+��(Y�K�M���-H��Ke�J�n2Ec��)�>]���a���@� �W�g7�J.�m,�m{ �l�k1l�����	 ���i���
y���ҵ�5�q���,N�b��aQ7�[ ��M ��G|lq����d2��� ��bi�v�����P���-&َ��YC��n7#�+��asZ,��6x6^k����D�;��&��Œ��I�@��V��:t������,��Y&șRB*��S��ָ�n���d�Qq�(��XTNz��)Sʁ�S�k��L�08LU:LAP�ݼ�i�h'��"�M�����h۩��JK"�񇾑�w*�6տ6ѓ�юX�t��?��O�I��P��xT�kP�<�l�p(�f�d!W��x�"��q,��6�HL�A�b[�X$u��gl�$Hc����9�3nq�gv� <r�+�$!�M�8T��K�1ߛ�qlр���OH,'�?�`��O	����
O��E�X.Dy/d<V૸�ko����s��T����<�n����,��)�D�Hu-͗���I��C0�N�4B|-�7����)����9b��$�������l��	:�۩�l��8��(�lq��z�ߘ�A��o|��)x#(ݿT��]7�?�F��������i����]z��Rt�|�ɝ*�*�(�*��%@�����,�O|}]�fP�Y;�H4X�7ٗ�/�~���q�@V����xk�
ی�dK���5���`��9`pz�/�����$��� lO��;{����KL�7#j:��������e}�8�Jz�਋�G��]* �Rm>:��Z#����h ���[����]�u�/IZ�=�x�v�^��N0B/�Ե�(��	����~�?lC��K�+t�Z��Ά��mL4�x#��y"H;n1a������R�k>��U^��q�0��L>�/7�[88<{
1�0#ߴI��:F�Ĺ*W�놩3�q ��1��`�H)2�(��e̀ߺ����Y�R�y��*�~�lC�0:�e�0)RaS����W�o��'TD�!�F�~�9�0��s;�(����Ҩ��R�]|�����{3o�'pTǱ�»�K�� �,&IB��֘S7V��R����+OjxשP}����y���v�h��w��b䁼�o�V�aۍ�H�TȮ=��Wӯ"��.y[6����^c<�8������B1.��>�rG��G�ۿ�/�t	c�!=i�5�$��^���wF��X�_l}�z���D��<�[��BٝeώD�O�8�Q�,D�_%�I�u��VE��=�L�Q�mLd<�٣u:n��C�
T�ׁN
��C�V�KRSq1e�e�]HW�*�)Kv��2Vp3/TJ�Cd��:����Yn_Ze]�u�o ��c�;��)�ݠ���(�=}n�Ye��J�բ�򩱟�*�����g!�*?��j��!��@���R�x7�ӫ�D���j���ﹸ�1"(�T�����!\��k��)�쟥:���H?���(�C�ֿ��QT6�^�����M��h�/CFa7r&��Mq�n�����!1�f�js��T�e�7F��˞"~m�MY�ms���F#=Oؘ%R��T�"�U�׹H�57�9��>�0�
cP�%���f>�n?��5����i�A�l[b�u�zL=������v^�𱑃8lk�TL�5�36���3U>˹�<W���h�z�~rO��̬�ߵ��G�/ ��� !��v�{����	���&��n�[�v�!�	�r��'='xv 6�Kiv�V�#P����kme�e����I�a��gl�È���&GM}�HX^�~6h����L��\�!~DVc��	ӽRex�����9�����v��5�M�Ԩ�
������Tpf6Br��<��:1b�!��i�;�� 0�{0gf~Ie��[�+��M'��'x���K@i3'��0E��
st�#E���|������NJ��G��<fOVZ0gu/صQ�A�%�vB�]>���r̄Y�L-� �;���+��3쏱�Ef�V,���:\Ņ�Rͥ�K�N��QȚ�����C�P,$0�_c7Z�ַ��J�Q|!��yoG
�xvWF#4	�W���T˦��χ}�Q�B��b�!7��<��/X_��z�i4J��Xԙ�%�u������yJ�R8y���L�R��_�|ǖ���@�ק.�R����D��\r���sX\�{��K��iy=3��.�v�tݓ\g[��#H����HQv{p��k���'��/�#2�R5Ȧ�� �(qD���u,���b��D�@Ƿ�lnLżD������Z9�&.���oe��E���U��t	�ͼ�R����3c���<�yy!���O�v��a�"PM����c�2��lz>��l��@ԅ�/@���:�M8UyI'^7��l�|TLd������L���a�E�u�>}�=�|��o��΂򾫕p����x���*t�Y�t��6��C�0�w������U�i$Zarݭ���ȇ�Ќ�&D�.���;��o?�r�+�/>�&R<h�`7T-�~�աO/d���PJ����e�o�G����}�?�:�sv�n������jB2��T�u�'W��p+ �8E�z䇃��~����X��=������ wy�F�Y��rbT!Y~�[��Ϡ���P�>�����I��	�]ƌŮ��&}���b����=�����s�?P��eQR�WU����a��Z�H �C�X�Ҵ��M�L���qS�:]n5�&�|�E��~khզ`gN��ֶ++��p:F�:�Z@
1��a��g�ֱ?�����-�U� 9�����׽2��3!�2���<S�����ĭM��)�H1�IT^=0凓Y��O�Wq�ޢ@%A!���*�)��c���١K�T�J( ��ȏn�%c~�m�}�~_d9ik4�X�T�R�/����I�N��^_z뼢ۘz{ld��a����J��tP��C8�Zy.�[x�Y����:��˞�����Ʈp��X��GD�$�uv�Ǟ�Տ�14�g��;v0���Xc�4��Y?3�5�b����+����pTeX��!���&�_2�D�YA�|�x��2v�y}�db���W����~H�{4u���I���*rk��HJB����)��U���?J��kJ���N��~N p��2 P!����� ������i{�6�jY���9�qoj����OKVv���fhOQ��ҷd�Y��
�TTJ�>�,�� 8+��z�Jp�.GSȲ���氝.�f�d�=yG���0Z�/>=;��������*�#A�h����E8��x�rCYbb�S�+�n[��:<P2�p����S�ؚѫ�	W�n9������8���׋,�,�K�?�#B���;`��L����s	MHm��+�qEb����_���5�KHk��P; m�������yHkm�**r���jgφ������W+��2��Kzzm�3	��{�=|/���u'�k5��&h�����Eҩ٥����n�����4��Ց��������Z�+<�R3�߼R��Ua��nW"u��4�TY�>�c9�D�R=����m�����Ī�m>r�Dl�[��;��]Ln];�-M�Rh�b�e�t��꣺���M�F�R��]fvi���C� g
�J��f^�b:�#��q����U{��T���K_�m�+/�^���%�꿠>��Y���^ât�K%�r��ג0�v>Yt�~ڋD�Cø�6���W�eG��{�bq.���ɦj�z�D<�����H5ccf t��|���]0x�7��BYNe��1�E]�'��D"���G�sW��v�z��z�ү�D����a�	5�Y 00U͗��L�:��q*��u��5����2/f�ֲ�%)��Y��䯋�z52��~�4>�/Epxb/���ׇ�P}x�l׬�n���ѻak0��cwE�(%G5�=���D�D6 :�@�c٨k�v>�l+D���^�,�Tp��h4�Ue��L��=N�HXA��|��>���m�j�Bٓ�*��3�&��T��}��)��S��T3��#(�H�~ޠ�g*M��|����`A��+4R�^�'v�
Ў�	t�h���>v{�5��R�[W�lj�+I�##l�`��R��q�Z`���﷾�琊 �K���*��ȧ����B�Ϳ}�j�XXe���!"ف�E�9�m��Qr��?DuVс���Գ�$���Fd�1B7�^��um��_�M@�ނ��Z�a���7������!��hi!j[9�K��v�yX<�1���z"�_%
�RT��ڇHEE��e��hy��4��|���F�wO�z�.w���Xǹ3F&���G��m3�C��$js�U}���,�Y��UV�{��#�]wD�d.Q@l���8�C]�D�>W�H0B"�c��y ����V��K�S�$���z�u[J�J�QjQ"����Q붦Bhƶ~�/6�ra7<T�R:=��[-�O"5Bt�k�	ĭ��kq�&O�[A�B���jV���|!	���IŰ��(k;��`'�_`?���&4��{"�
�3TV#��s��h=��i�8��9�[C-G!���ŏ�˸�W��u���6�Ieg1"R\�1��-9VR墸��(��Y�<�'o3�#w��<�8tR��:}	S��"Eˣp<r���τ��8��h+�o�����]�٠� �#����z!��}EJ>�NC�'��@�H�^Bg�d�a<Ӄs�|��Z�����ȢӑN��=��+�8��t��c�=��,ξaQ/՗^���.P-�B��V4 t�R3��\�U��fN�!��7d�@�#}��7�ݓ 8JX㒾��o�oq?�l���p� 9��\f�������q�߆Z���\�� �5���AS�v�m�W�h�
Kg�a��x%L�x�\uT����1�=L�~�l�߀�z��r�+D����	n3��o���d�(�a`����Qu����gC�S�-���<�O��E%��C��ST1o���\g�GNi�$�M��`�v�:aRP����@��H%�_�B[c4�9g
[ClĄ����7��:�-����%��
:$�MV��&�3�4�eh��n�jF:�^Мρ���4$�2Ƈ/���E[�>�'��5�at3���,���7��D�i#�6�s.��2Ã$x��ʙt{�Z��Wؕ<6��'(p��Eǜ��C�Y��`� SgaF�l��}�����|!����s�z4:��l�^P��cNr0;��h/1 �]�z`�]�@z9�jl�|�����o�a(�H��)r��+�H��T��ꌤ<ˆ!ѫ00�X`޾.ׂ1��S���+N�y���^ҧcP�1y#:�;�$�����J�%�w�⭁V����9��z���F���e�L�(6H��� &�Թ_j�G��`F�֏�������Sא���%``��� ����m��N�Cl���4�3���W�_���l}���R	������R)Ty������'K�� ~?;�+�7�D�m˘�z�	'�f���DY��C�G��;[��~��m�y�~p�d~x�"��+��l�G��I�	�y��j���}���k���᲎�`��N��[3Lۤ�BT�����@������������-CU3$}�j�k�_9_��M�|�����Ȥվ��v�-Ϊ�u��<2� 
9��'�x� ���dEBF���;/S�B���Y^ù�'۟�:IO�T?���[%��4{ �N��F'N��'Y��� ��̿h�pI��N��	\�߽���ٹ�eç�]鏤j��uB�<p�|�f����ޞ�@ok�_�t�)[#(jk��4g5�sd�~������i[xAF���"	���C�)
��i�d���o�.� 7��K�9w�7#�f,�����(��L{gE�H����Z�ũhY�S5��w��1���Y_�?����>�,b��/�T��%��˂�j�O��G�M{��v����H�Ɖ�S�od��k!6��h��aɩñ�anxr���r����r��6#�{���b^�[:+�N(&R�^}#�ɚ����x8�Dā5�QtTP��@ ��o��,v��A���\�:{p�2s��c�	ٳ�Jy���<1p�@�m�?� 3C���X<����R���39�����Ѓ�u@��AE���vM̫շD�[9�߾���+zv\���&U�]�kJ��3�>:�ZXX{t-g�x
<�MA��gU��"@&9i,��	�
��qH��m���y�����.�_�צ3�/6}[0��ق4P�ɸ�ne 5���;q!�f��`pk��/�=X'��
A�`�ԩ��a�(��-�
����`����?i�g��H��ik6(�����Pt�䍱�l��ej|��ݫp�u��o���DR��|�Εh쿰�6 �k�����#ڍl�=5�QP���'�k3UʗS}!�����moo�3j��Υ���u����ŗViN�_�,92|2���%��]�L�<�d�Ի�r52%�l�Ћ�"�2D�5�|Ro�Z�sE�.�#7�����Ԧ��h�m�������[��O�O�������Ύ*UT�[��kC�-��L���#���3(g:$�{�h!v岦	�!�B�T�����B�؟?*���R����Bdd�ڮ��װ\�(�5ޛ�'d�?��oc��i0��AYA��e�T����P���u,	�-�#��*hG�Ԗ%ҨIm�3#4��u�{-�t:�ۨ|�N�C��H_��DBM
��-�>q�z�#�9�](��w��:Z*��Y��IQ�OAUI�D�(#�aB����;�
�%�����5�D��`�NP]ك7�t��	�N�!�(F� ��C�Fs��Z�g"ӃC�7Ut�)�3���
2���Ui�}~ҙ��}WmG��˨6;�ԘȥSu���\���8�!D'���q��y]&�w*b+r�3m����T�Õ�y���
ڜ�	�͍��E�����i�rm��������u�v�8F�n�-s{p\g�`����� ��g�xY��5W˃8X�;@S؞��j+Ud�"�Z]�3K!īp�<R|�����Go�9�Y[�ɤ/	�J=u��d�A�0q���g��ɔ�Q�¨����e�=�[��\@IQ	[�5#���$��˱22��K��]�#B��0�_܈�%��2)~�F��0�ٓ,�ǠNn�^��F|�0Vd"ș�譲�%�zn�@�Ť��
w2���|N��QZ$�����sd�Km2�S���JM�F�3�c3������R�����mdP���ѯ~u�XLgrg��9�	y�J���?,w��j�d�j�	�)�=�8m�sh�o��290�	�7��g|tt�O�&�v|&h�"���8�N�"�g��ຳpV1\�>#������b�)�rsZ�H� ��7���4F���pQ,��
��^	����/��w�����&�9��C��y�~�c󤽐���[�L��i$���#��r�MJ�������J��&>x�}`�x���w�Z�2�!س�%�Kr�)�>�o;p+_�vN~�,a��H�He�:��/_{a�'Y�� �
(������}���9TDN3�
V ��B����ｋ�e������T�{�c�/�-��ko��u��X	ҧ������{��{H�p��A9�b���e��8�`[RZ�^r���+�x�u�j ��͔��x>�sTk}�XW�I:�uڙ2%��[��u��i�ޱ�V ��OA)0�L
��M�:ƻMaTy�T�lu�9��V�#bRegض*����R_A	qڡ����TI���J��*��K/�>v�;LU�����>��[�h1�(��k/*�0��8�Wq*{��C}PʚB���U��8��c#�رSN�/H��!�Tv�57����^
@��#�<��O���83$�ꥲi�E������s�ҹ�/)�졋�^�.�.ZV��@2OV��G0�|A?��&<_�y�o��!�/��~��v�������,�eK�L�1��[�����e�|���Kl��v�ؔ͊J Y� ��g��M�X��xܱrJ��hA��b1��7,��r�[�����P)��ȡ^vʋ5�=޻Tݜ9�G17U�O�s�޶��R� ���W�]��������n���̻�CDP/����;p��P��D�,U}��TBv��\��U�RP����8iW��R,{��nD�QiW�����O���8_����&�P��<8��e�����u_~��a���,�D�|a�>[(%e���KcXMo�}5(�m$��7sS�sT�)$K�4�zs�y����6�QZ�<�ш���n�1Ѝ�1r�:pd��?#@����g���!�^��J�E��,0��N� Ha���w���p�H
�	'ӇD4h��梌�}�tt���&� 
���1C�%-�5�K  .��,Ф`��,S'�k^t�2-Ŋ��F��m�����{��2J6�G��%�#1�������%2����pٟ���y�J�8f� ~	$o.��o�g`2�`	n�8����3@�0>l�yQcWKk啀�R��#����0�,ّ�jo��F�}G���k�T��4�$zk��p�Ui慡@�\�P���������[Gz@�6GܦmC�`���tz�XL��p�ft�
�8j���/�{Pc	 `22�{.��r,A�R�"Ad��`��L]�x�[+�,�^�Z���W�p9��n�ސ��F�f{�&��] nL"�|V�$���&�\h���qӴ˳��k�i�N����
P�;��r'�z���JM�Ȱ:UNIm`��PBt�Z��+�x7雨��j�m!L�#(�sW���D��7�B*j#R������pd�>�p���3 ��`��2¹D���~<� ������u�d�p�7����bP� ;y�1G�����m�8���$K�/��������W�9���	2Y�^?���)D��
��w�c�� �iD]?0��!9\/��Z'��YU��cq����@ �T�=Z�n��6�_�'r�X�
J�� C�x�N�5��	8)�����r��DyJ6h��ɔ�&>e�������q��rw��T������+����j������^��^�e&��s,�W
�{] m�gs�?`J��(¢n� k�݊�f�j,Z
+�9_ͅP�����ѥ*}��⿁_��O�КԘ��[��-X{ƃ�Aӷ0#	v�=A���M��f�k�!�ꇴ�EuNc|Q�2&��^���|�Xt�"	���T��޹0	�ׂ�C"Q�]v�yk͂Õ7��&�m����#��^����d�5eV��>ߐ́K��{@;�J[��d����ca/%���?Ne+��b�D��V����P�h�n�H�����~��E	xƵ��O���o
�=�|�.I�|����V���X��6b�k;Fp�Њ�p.�ιz�!�|d�Et���4�<f����ȋ��&&�*q<�{Y�i����D@� r��f=�u��J!{�lCU��g.A}�����~@{vś�ia��y��\�-���ʶ���\��t@�8$Xx���x���Y�pȔ �Dߢa�MD� ��}�PuDܥ�'���cǋ��M����o�y���H�>���D�g�3�8�_�f�m\�`
Ŀ�֩�'t�
5/��'ӊEj /5�n��F,��e'3��`l�'0�Z�q%��n���L�'~�ڇ���+k\�.W�l��u4$����	t�B�f�/�ї��v{��|apf��v6�N2əQ��t�?�X?S6t�(�ޜK:�E��1x�2H_ϝ�o��Isg�wڠ��f�$��V��T� �)�BQ�$71E
��p�p@e�9�ZG� ^�����H9�,�c��Q�+ �"W�%�Ѷ����m�lu���6݋�ύ��Vm�f�%V(���|�ȁ A
I�-��O�����$��y홹g�j��Fq�\2�آ$Y�b+�e���D�����b�t%˃M�%��#d��BCs�?s\�*4dhGHl���+
��F�{�]a�a���!�؃�j7q�KkC.~�/2P��<׈J]��$m3$iP;Q�I}1@K_�����/tƭ�m�錋Ԋ{Ս�c|G�c�H��u��㚟�C\n�����P�=�/�:� ��60m���ӑā��߱^��5(��1�MSi7^岊W���F�'m���/<Q8ą�3Xd�',3���8V��f��w��u��&����=0�`���؂5֟ -7v�����m��F�����ͅ��Gn7<9�`�Y�cq��4���I���u�l��|1��myT����%*�G�؈2*8����� �0���bt�����Ϊ��.r;��rd]S�q��M�4�)� ��M�;B��WM�+S%m=(�8�&rH�@0�3�bq������4g�!�SL�dy;3��ѹ_f�t^ z��#!Ԣ@�p��E�*w:�++ME�x����Q�n^�C������y�uWgM������/R/�P��w��.�)H�^�K&H���+��ki?b�����>?���(�7Z�S�o?�{Nx��~:	-�k���k���]�2%L��!b�ݙG��hy�yHxSGB���0z@e���A
�'7Wx2��i��1hw����-�0��=��y^�7�|��kkO�1uٯ�ɫ�+iaX�J6 ��<��᷶Iw�Ze�F�8���s~��Ϳ���A�a���.C�)���,����B��[z��A�����c����RJ���9�¼BQ;���E���&9F�:<�"Q�.Vp���I�iT�}�o��u��n�77E0��Q�d�)2g�~id�T�c��� b3�a@������
�S��~��@s,i��QTYS����)y�����L�/�c�C秐'{7B�·0z<b������ϣt2�8L����f1T_}8�b�@�Gk�[�X����Ju���+%�����՞�,�R�<�R�*�cV���4�{�2���i�S@�]U�,�����U�}����jcuf,��f�z1EZ��rP�y�)����V7Ǹ".���5�4N��}Or�U��A�U&����P�te�|Dٜ��r\'�$��6l��4NՈJf�-��g��QAڹgq�֓$�TRf貴ơB�����db-��Ʀ� '�nQ
��Hᵶ.7V�82`*��}vv�)����y��+�H|||ﵘ�P� �]h�PF�w��۔�A���<�Q��C��U�i=�򀓥�S�cp��ߨ�p4I�ֺ�MN0��c�O1pz?�	�Dg��#�v���v0D}U�� p\FS�0�`F��x��G&���x�J��^hG���D��l��#\\p��ɠi�t�o�խ��(}�.�Aw�p���D��7	��:�O,I�-0=c��ϧJe���@O������n�2Ti4Ꞟ&2�Od�I䌅i��Q=�qA�]M�O�5+��S�-�� �gA���X�&��ү����%�E�?�`3u���U���JI b[<��?��<�i��^��/E
���'��Q��o��-"��7�'E�a�@v�/���%i����lEx��ų�1w�!��A��R�94���2�x[�_�� �����Ɂ���ZzqOs�mAE��7�F:=�T����ۙ��B��g@�˦�h�F�%���V�e�`R����uڌ(H�E)!J�q��3t�ע��M��h�ϻ)b����Μ���q��CK	��6eh@�����?q��śX7ӕV�®�ann7^�~�0�8R4��^�T)?K�6{��꼹V�j��E�?E��P������ߨ��*���(~+��t� q��WD?*+��Dr�a���*�M9��omqq�$_hJ���O�Ŵ�>�1�g���D���H���ʴMĉ��C,�ym���r������'����nҒb������<]��4� \ku�����*�l�|��P��\w�(�����<�v�LGL�CJL�Qv࣑q)n�V	x1Kf�t�dY�<���?6� jϴt�݁��emI� ���� ��@/Ys��̈́��*(��N��\�3�����4\��H?~Ⲕ�5'�e�u�8��+[��V	Y��3l1]�,�Q�I,�4
�	!���?*،t/�d͙�?�:7N2ƫ�,�D�?&G�� ��i����NNگr�Ym="�%�\(��ޝ�ǃH�y���x9���L��c.˰��q�~�$�ٹ#����]y�w�r֙y������ڮ�YN���Pς��*a?�k�>X�� )���Grƒ�
�p��ʘ���&����L������� ,K�Ϩ�����
\�-��5u�VCGh�$q�.d���V���ک���IԄ\��<��)Q�ӆ��f��e��S.i˖�b��9��g���o�]\4��97�ُZ"�'�Of=�X^dV&�s7��.9��e0V���ꇍv����w��ƻ�OQ�W��A��������b��Rp���Y�%��u	��u%ClZ�RQ��EH�N}��ݼ�^ %@���>
k�-�����|��p�:�@0���;2=��+'P�
���H�y����� �%��B��9>��lt6V��s��[�olWLm�=X���f�ݑ�!>�/�^M���ς�b��pH�͙�cL��%�����P��LE�ʳ��q�/�bs>{��ft�lL����;���q�������[1�;�I]2�����V�!�~�gg�a�r4Ә�t��/�+e����\E�=J1���RQe� �����*�
���3(:�	P6������T��%8N['F�^�"ޥ,�ҟgc!��i�JO��ɔ�y��r��5Տ�ą�ɴ�B��g��R�'1�p|�GQ>d݀d	�L,C�@-���ܩ����9%d���܎�.3��D�f0�.^������$�wtnP���ol�����Y�)��*� U�3�[@Y�{���yم@{b��g�!ׁ��
���L���(�&���5�����d�������G�>�{ǦWhkUE? T���V?�-4ұ��mz8~e@���������i"���sd��áXˮ��n�O��jީIE�Z��>�=%�@�xu�lPz|�E���j4q��?�؛�"���ۃZ-|�É�I�J�4A�����3g<��.�J�%*Uj7�g�b���IX�)^��e^��(X��Q<�W��%&D���b��������m�@�������l���A�G��A�F]ul'��&��s�C�Â��:�87����J<rE
#�B��bv>���v©��<��Hx4�� ��@�M����
Tʙ��Ѧ�	��h��,6�z�щ�w�jb�u��$2�Z[�@�P����������f��M�CEL����0e�I,�K���_��Ws1��G)a�a �BOǱq��*��e,#���	+��U�(8��.��Fe��	�������20y�/H�����SxQ)֔�c�uޗ�b�雥���3}�ڞ��(h;��@�q=\.�t(z�8��#�f�u��pk"�{8a,w�S3&,<sl�C�I�y��QQ6/d��� �l�wk�^�o5��B2�T���������i�Ȟt{�h��%Ս8�ךt�)���w���1�4g�������\M�jdB5��s �)7s����E'�ܱ=�
eoS�17��3�y����V=�ƴ�e�)����n�ɮ���T���bx�ڴTtX�g R�m`(zj�d�N�_nYk�L�mm{���ĥe���U� ����H
�b~o]�v�<vD��fL�XM󰜕�}�ġ�@�ǎ,�l�l�o.�E�]�J���HV�z���<#�x����z����J�Ltid�>o�X
S�9�K�����"���<�-����������L��$�%ۋ�Z�4��T�vY��	V�eg�ؒK�D���V����N�p"�P����5�/(yr����(�fJ����k�^��'�ԱY����&�n�-��5B�ߌ	<&�8h����D4W�Ыg��qo�������Q�);�Q.��;��^p9�;����\���w��x��:�c��^ ��3k��O�T����$�����Lm`O}e�mڹ��}9��%I�o�q�G��Ŝ���"3��}>wb�1Yک���8��J�g;F��"�ꆋ{�{u��I�}@�"�jV~�sG�Ha�t�"U��#A���E����%���%ޯ\�˗�}�?��Z�s�����yQ�\��E���&aVe�	�_=AU���FK"`��\v�5��(���
�-a�I�� M^X�����4��z_�0n�LmH>�\۳c���x'_���<2�r�G�t	�׀%O�I(�&�k-'a��MQ�[O2e%`�7v�P���nӻ�v������/B0�d��/��o�loqʤ㖖������ÐI ٛ�
iC	��9�H_����v�69;��0({�D��mG��ЉHQ�WN�s8b�'Qnг�T�J�$"D|���L��":�PLq&�ų���B�!,�Љ�ҁ����Ë�V
d&��B�1sK2F��y�������I�RQm�۟бb�O�O����Q]�L���K��%��(;�8A����	�hE�����gJ&eح�k�@�V���$?/|����&�S�.BFI��=���9�i��1��q���Ge��ja��tZ��'�׮�}<n�hx�7V�[�.τ�0�ux	�m�g��D���c���r���:�����L&�m!�cG�R�i���j��2�D@iN�DR�; ��	d��b���4���s�c�!1��Ɩ�woC�ѐo��K&��lqJ��0l��� ��%I�Z."��ITޣ���vTl!/i�yI��Z��܇Lx8U�>��5;I�S�kl�S wu����A-�6vm�	!TL����j֬������D�0�m>��mi�H�q�	żR�h��}%�j挒ǌ�Y_	��٤��Rv�?�úl)���5��D�n�
��������&��~NDh�>;J���e8|�[  ����J@���n�3�3�5�zD~�����L�k�S���s�B7����*���1��t��
�v@I&���Ҫ�\8�^���R���8��.avS�ґT�����,U����[����Vx⁹7E:��G���U�fB���eE�m�a�}�)�'ˠ���x-b�����rpN�������a7{��	9hv��7�w��B��c�ҁ"0n�	o�^�X��S�o�:[7?�}99�v*�v�a���;��J��T�}�Yތﾼ��{:��%�M��<� ����3
qX�iL�i���P����M�e�B��2�s%���㑥��)&�d+lOxۺU����P�ɣ��{��r7��Y`�S?��F��)�<�W݇�y�Y�3�Lq}���I]ex'8�U�����0@@�>V�́��9�9��Nq�p茴�%"Db�gl��ߢ�.f^�U&�%��1�7���	ܟD���Sj,�>'��_JtѬ%��@J��v˾���=����x��U�&4��QCFԱ���T��9� �±]f��������8�vm"�rWO�d��k�eD�E�W�x��c��w��O���_Ș�J"��ҵ?�%ܖF	ɑ&���wXD���r�r��#�s��x�z�TLx�O����ID��%���RÒD�(��$� L�s6��m�����tV����
��hg}|�N?�[�VQ欰�H;��{~�E'��6��?��[�`��^�hv���J?�f
[�,���! 7�E1�eҜ(A�
�����=w&��~ �r\E�@�5�V 9�K@gA~ɟ��#�vkj"��n1 ��G%(@J�Dd�];Q�<���H���5���Ӕ��P�J }R$k��S��Z�b��.�.}�}�����W��u�Snf��-��:���`�{�ӛ"H���\W���;@Š�(���P�]�{�G8��ZC�{��1��~��\$���L�8iv���Ii�۸�Z�)Cf�q�l���)�큐�j�qڄJU�^��lË�6�AC�S��%�u �XZ���D��\����ۈ"���5�����{����Y�6��K����b޵Hk��v����n�*̳ܵ�f�wX/Q�����{	I���]�NkU���ȁ&��q6l��B8��I����RBm�K:����XR�A�Jq�-W;"?B��^0�'���&�����F/�<�kE�%O�^�ރgx��m#_��m���B���}7E,k�,c̪6n�#Ͻ#����Yd��@Q�f�3�x����|�d��\�Xc,��b;�6S�����,W����5�~fE�M7�$���ֆ�Fc��A4r��d�}��]Og��Y�z ��.E������1�;^o��<;�2_������o�m�>P���-�� �pu���C��w/������hݬ����Ps��c����d)e��_X�Ը�f�M���8��|�V��t|B�TS����
n�vv�	d����>�*�Ϥ�:m��Kx�S3�}����LQ�d�i����*�y<ߡd��x�'�t��D����ӛ��~1o�i
�Y聚\
��m��9ǗԱ���H��+۩�[�^v�G����la�A?�E�M��4������]� 2a��+�n;�� 2i{���d�Ep��~�� oő]�c��A�Þ�r�O��V��i��'���~����a�#����~3Ϝ�L��t`?��)����	�򒎸�Jns�k��M �͐',D��¡ 2�g�B�mj��R�%LL&�G�f�Xq�C��nGura��ԗj2;ci�r�l�g�`lT^���hB-A1w�������-΂�t$�0��&�%��{�����r@�L���HQ@%��T�����pI�[�����V��������̔����N��5�ql�s��`����Z�i���@i��$|D�=逨�O��
q|q��P����V��V(^z��	kNsO*OB����A��a��%�*�8�^�}�,�}�ă� 9_ĠA��k4�v@�B�Ae)�eL��'!SE���z,�y�Έ-�h;�jD����D��!�q�q��=]��lz��M�T�P�+Ȳ�?7�Ri5�o�j^6g�5B���<Z{�5��;�C���2J�`?��h�)M.�-J'/D���U�a����>e��Ό��:=6^��4"��ӿ���U�c�F�(�$2���m-{ü��A	)G��!mAue�z����ʜ���5����Eېf�o��z�U�N;�N�r�/[6�ޅcԽ�Ր7M�c��}�.��O�34���ի����ұ���B(��9e0����}��K����.�f���
�1ӑ;dzo�t4x܎!v���k��cy�;�-������Ӣ9��)CR�=��F��������bw{�q�A�s�>Z"]˽�*��b4�tJ�	;ns�am�V���>ͮ8�L{��p�zIDy9*h�{����bd�`иO�ϒ�|쵄#q�R�J�k��n��xwo�i5���ʲcq0��-`z��?��!�^��C_V���DP���8ش!xJU�gn�,�zadeJ�Z2�S����@l�yګ.`�'��'�uө���_l����2^8�Rn� ���ݨb4��w�ٮ�1�5�^M*/��a<Z8��S����qNL�� ��௢�J�1�乏܇4�|��?�M娙��A~:1:��{�	���,Pp��@��x�Fح�Z4�K���~�p�LI�<p�o�'��ӄ&I��H�:��>�b�����-,LWy��[�Z����F�;�ŗ�=�ɇ�42�ы��k�]0< �����i� y��;��j,+c�N��#>�e%U>�G�Sc��?`���ܰ��?Hg]W�0��������Y�쪏�I�]]�dе�:&	�";����Úu�� ���@�+�L��~4:I�x��=^����H�߻qAQ�o70���W�� jw\�}�	��L���cQ��|(E���e4�[;����n�m�tz4a�U�%��OÅKUz#a��-��r��#�s��7v�Kź��]����W+8-�_(0��u�$�����yv�T�_{2��X&? +^F����o����L�"���� `�����k�|�+R�Qձ�]Zx��Õ������߭y6�B�r�����N(�e=�_��Q�o�'or�*���[<��ļ��?`ʣ$�H\��o�O!uu��>ݾ1�ƻ��/J�1VKQMB�iE�RM������Z�e��%6-C:\$x��9�c�{��i���L����%��_i_$6���H~�X���4jT$�^�-��>m��;/��c%Z�_6J�X[�r`3�i���_P����-cK�Ǜ�{�+�V{�;�i�Y���c!H�f�Iۤbk�-�ȭm�Zv���8��:��ꩳB �kP��WO��H�!4VQ� ��V=DJ�f5V��l}H�x�J�Ҳ�e���VM!x�$����ŷ�W�K�K��v�	dp�D�R4bUt{�y����S����)-s�A����6�?�z��ߒ|Vל�.�𱃁�f��3���Bj���ثvx�[���:P)8'ܑv3..}9�[������2��=w��,���t!���W��X��Da筒Q�9�7�/��I��U���u)�9h���q�͟9��\����-��l
巗2kѼ��(�wze_��~{]��d� o�7���1����(���H#r��.9�7��FI�PX}�>&y#�%��x�&��~2��2����(��i�@��Ȍ�)��-�t�d�T.�E�ȿj�p";�.=�g�ؒx�d�w����_n`���lOn s]�R`�9�Y3���+���3��FL&/���rTR!���WK�=��n�2�+��V.��������8����,4�?KQ������6��ĲaID��)���5 L�!}��g�	�1d��da��N���=x�h��� ��L��wp6���Œ��&��Yd�v�J�I~ ��j �=��O��"���mOܕZ��9[)Zt���=���G�kVc����<�V��談k�?�S�Ԫ�J[�u~q�e�Nn�oYl8r�aڅ�T��.r����0.�!G�i������bT�S�Wx%R��E�[ż!�����L�*��*���� Kf&rbHF�l��Y\�(8��Ls񕛤�Ը�$�zjǇl;�#��mo?�{:2 � �&T�~�뽪XءY���J�2�w	`=]S�W�����)_z��'4���Z����~���m^"� ^vo�?gɲ�[a����`
[�9yv���ص���r����&>_'6>��ˣ���5ʓ�GA��;����;��9X>6��}Q QXY���ZU_;���Sg��.5C�Q&ޱ~�l
���˚m]Ҧu��0�}�V&bn�=IU�̣ ����Wq����B���<>��RW���)��V$�]��އ&S及.�����f�<���FȚE`���F�=�������v����R$N����}
Vj�2�}�����CF�R��ë�PK|�K��t����8"7	��jRC���:z�jgz��e��-#�3-�c��Kz�e�'���\�E��_�G��wL����=+S���cl���zH��Mpu��d�D������FՍ�V�5A���I�aW�q����|��=�mʹt�Q�1�V���{m/P�u-qLڑ�-��3	؂7?�@�N��uE� ��+5�s&ʪN9�<�Ϊ�`#v�T",�>grN��G#���#��e�%~/H�5;�+H���W���
�g6�A��Hm���o_�+�~�l4���\^�{L���E�M7��8�g���׏C7�E�8AY t���C(���4Iݦ&d��8h�\s�q�G���^:4�2�>N�\���gS��N�a��Į�33T1P"u��WO�=QZ3�%�k��z�u	b	��pKnG��g�{�9�=���k ���@��nt�g���T��I�|��v�4�s����#O���|��[s��IdH��(� OA�r0�\ke903�ވ?Y�D�u�Yz�.�t���5�9q�h'1���	A�[P5�4���H�u�gPq��P��6�åP5�9A�.�^ߘ�\�M1���D�܄k�w�FTĲ�����3�F2�t����{	>�_��}&�E�ңB<4�~�f"���>g*�i�� �ӝS��kZ,�����.�~�u�*ې8x���~d^'j�q��Ud�"'Gv��ۣ-T�E�b���Q齊��������:�L[��ͥ�G����:1�� H�Պ"�Jbֻ�먹R��Ɏ���*	I�T�E+=��
��'�{�f�jnF�Ȭ�,�HTp.�\5&u
�o���U�Q��N"����Ⱥdfc�z�<Hg�ڜhe�SA`���7��3��,�����M\o��TG�?����;�;�Z��+���#:�,������pp��I�X�I� ���#]����φ9�'���%���9'�:�bE�ᦓ}��>�ȹf�g�"�@u�5,����Y�s5�c��s�)�k徿��3ɥ�`6��XM��W4WBњnC��G�/c����:%�P.��	@�A%��z�T1��Yn��|f��b����Ś�2D��	�(����w�'�5��\�H+��S:�1����� |�Y���a远x��#���kp��?�PM��[��#�|��%�X�QV3�S�{2�0N��kp��n>C���<%cv�󿫗���1B��k.�2��2��b�I�Ta�7�c�ݍ1VK�aM���?~V�R��Gv\00� -�)b+v���oL|̪XXb1��@�)Q�A���c��7�����5o���i��K�{5eA�ʓ�6B�Pٶ��\�g\�kw=��.��'��٤���Ku�I��0�y��q��Ej@�L�qh�N��F�ҕ��-�-���}졿olm�=�����s���_�p!� �j9���[Y����K{�4�HNG��6B�8NVɛۺ3���B��#�-/��S�¤6p=�lN!�N�Eb�
�+������������Ф,�f �Ba80�5;��G�dԨ�f�@�a��������(f(2<�殨Q��B5X�f���<'̬9#�,��\�zБ�,q��
N��iW��X�M[�k�k���l������pz�Ǐx����`��a9����lG	2�\�4�$�`���sզDݥ�
|3�2+�_&���
�W�g�_��&cl9�D��8��A0E�^�}�PR�H��6N�{���*x�*��{�=�2�q���P'��]�z�k]�r�
�,������U!^H���ܯz��ʭܾ4�:����@��5��C�ټ}ɝȣ�<�-<fe�}�L�G^�T�D��ER��!�lT�=��L!m���)�p帛&���kL��:����q�#s\}x�|�6 '�q���{C����Ro�y�W�[�vZrk=A!�$�k!ư�T�C9���� FO�F��v��:��x����;�k�S�2on7���Tw�������!�LE�Ґ2*'���zȝ�Ǉ�����&O&��lߑ� X�]��^�v ��x�� ���=0S�������6����h��Fޫl��33L�����ݫĪ7�]�Y��K�0�S~­Y�	����N�ZJ��^ޣc��_J"6���-Rx����w<�����3/B������.�9�����0W��l���JIG)�U�3��ؾ�{$��=LPԍ����R�e���^�W)d�?75��� \S�LP	�����k��>*QP�I4���Ή��jJ������q$����Q�ݙ�O(m�K�khǟs�x��������:��a%d
�Ư}�#���L�x���'�%P�x� ���ݣ�[��ِ���1�E�F����!;>(�=jVƘ���{��j���MU"Xc,����i��϶��H����Q�Ji��钎�l�n�����`;�3(S��M�a1�������r-V�:t,���	�
���^oo�5�6=9�Z�=�%�E��?��6�%�z==�A@:�ļ 0��nImk��\�ٚM�{UO8��ZLAP��&�Ħ�c~"+�
��daF��ާd�c��(���gZ5�c��C��TjL�p�}[{�_,W*�|&'������@C9�{��Ꭺ��,i�rd\H'��W�����Z�����]�5�6�?{~�] ��3�X�M��Eas^
��J�(�覴C7+�^�Z`f �O{�vU	L�8Y�#iz��P>_f�u�*6�X�wDIv�Pǘ@����ʉQϮc���`���$���OEJ�#��_��BO���L���՟7�*��O�K^��[��`��.���	�ҳ�~��T�3>f��o�%i�TZM̠jC��]4~Bv
��'>�ir1C���慩���S�W�60��+4H,��bXd+ۜ�5wL9qN�1+ExӾ���#</���v�5�02�85�2�6Z����bteT��#a	`~�wf�4�,dQb��p���WM�-3�I�z�T[RE��F�z*-��TLV�7�y�<H1�?ɚy2~�N���T#��Z}j���qza�{/#�ӥ##l��+�9i��y~k%�Α�_�-�v�>�a��K�1F�{/
�u\�{ڭZO/��~v{x�Rn㠱|���B��\��C�:��Ҡ�ĵ7��i�O��[l��B,�$D!�	�~����a�����7��Z�[k,�d�+l��n����Sߍ�#0������k�����U��-�X�͝硭���`Hj#�pwRU� ��N�����$$ ۰9Gb_x;�Q~*)h{���S���w4�,1�%�p{NQ���� ����iE��#�k��:�Ǻ>����P�' �ʅK̳�ZS`/3إ05��)m�m��T%�ϴw��={��_mq6Z���*����>BDGׄ�JB�:��י[����^cV��\v|��hj�O[rӒvVA��p�j����������E��`�"�x8H�m#�>���l�t��Y/��`��ƫ3��گ� �Bv<��q�4׏K�p��&2LX�@0��d1�$6+s⬱h�L����m����SR�F,��P��[�k�����t[�M�QЋ�{b��,��M RxX;XU[��6&K�UK$�`�آM���SH���H�mn��L�01�+c�&gwD%q�q�MH��:�YzĠ��F ��/�B�L\h��}�
�Ħ/d�ܛY���,?oja�?5s<�B�t	�x���o�9t=Y������[ܔ+V�:�k)�k�����~h�������p��Yқ���"��l�-����m�~�n�F�V�x`���~C�2n4ok��O���&~�.>E��d���h��Yi��-h�q+E(j��e�3��s<�9ZV��W����L����؎�t���$��W�n5|e1���S�ta����s9������}�1�.e�2�yq���,�}�T�n���G��:���h�@��z3pK\��2A���@{6�m\T�A+v�������¦��2��@�[�;��H�:�J]����]-h/�Y���|b�[���ub2T�g�M�&�i�Fϡ����P]$� h˺~�M@L�]�B�����vOֳ�o�|p �8FZ�$/�����Ϲ��IC9�%�5��a�����%�<�*�	�צ߅���hx�^�MHn�G4,����mZ$�6�	2�^-7ǃ�J����$�&lTt8%�5@�n!�S�i�N�4��Yn���e����}ȹ��H��m~:��"������pT�L�)�̌�S��ݤ/�Hei�>Z.�*:_vW8"=S��}'D��u.ST�j���{����s�3�(���-�J��P8f)�m�� ���3Q�����3;EM2LT*V�R�R�&0�ocuѼܤH�6�hK��8a��o���t��(z���"�Ѐ�ZA�:qh��c[�ϑ�<�[��c�@}߽��Z���B�~�E��tK�K�P����W
T�:�������a�1�)�ޗ}���J�O�<%�.
�kt��kf��dj�����j9��V���)��L��N�A� �N;��K�r����kv�X:��q�^�t>�}� D�"�E6o���6�Z�Q� ��f&��'���S	{��U��'8p���51z�+%K��u��,kN���I��92�.,�ڥ��O>"<e=���M_�u�Ŝi���RXՁ=u,��D�N��k�t�XQ{��A��L���_O8.M��ʔu�ԉ�D�O���U!������z����i���� %bjhB�Cx*�`�jU�.�Ҡ����NAN&�H �E��x���ge����P�)�{_�����bڡm�-D%F�hs��pu{�.�����x���l�:�w�������+��ϳ���@x��zEth���A�0xv��pE�1=%l.�d�cgs��rZ�ycW�ޒ2'��i��8�}KD�$Pi^N݋W��_X�m�K.���@Hp�\C�TI��r�d:Ϝ""��G9��â�,��ؔ3�bJ�{#�/}F5���Mˣ/zW5�'w���":^-�8
��d��@f���AN�0���Q�yJ-�����/Í͒���y�����X��	�T�Q���c��>�6�|,�J]���Ϝ:aw��n>D:S�Ыpr5Δ�]�ԁ1�klP�,ٻh*Tx-5�Z*��pB՛�r�5��j27��4���Z���'!�1�yV@�L�-yn�Ѭa� 곞���3&&s-@�W<�1R����xv�yC�Ӧ�����ϑ�%'Q9��L=zL":q���(&�u�e������W�D
>�h\l<'�ac��vS�G����]AHq���YBt!:Z�dݱ(,T�EG����b�6E�7�&=3"�����K�A�JTk��J���m��x �|���Ѝ_����!�hc�X�̿�{M�}�����k♶U!���s�s���pn���w +�2�� ��E ��L �*��T��7g��4����۹�����VVG�2��s�`����<�7��9�qc}ͦC�Hݺ�yX�o|j?�е6�V�ï�r@�ufh��\��|x�O$��+o�b�v�E��z�C��?�`�����G��Ɂ���� �{;�ݲ,YxM�G�YY!��pƺ�c��:(��B�����Ճ
�.���&^�L���M�����C.�n �Y�>fĎi���Og]���Q���o��q?����x=�j<�A��W7ڊ��	�8u�d����/�6(�t��r�]�<r�ȿֺb�fL��]]�R�E�8q��3���<P/Y
�"	b6��]:�\��93�H�8aV��b@I��܀���%��r�Ō�t0:�tL+�o/?v����4�i"�����(�d�{��'��(�'E�Ӌu�^����Y����<��O9H -��i+T����Q���D��Vة���T��l�:�j�D� 9�D���ͼ;L@�F)�M��#�	�₇��c���MYֵ;Sq�2c�h��=�m�:���#[�onW	X3eE�x���̂��FL�n������!�f�j�#򕄃�d�=S��N@޷/�?�W^�秢�1crҶ��x��_�����j�$H�7�uߠ�9>,d�Ƨs�Ș۟:Pg�j�>%iO�M7O^T�2�ca�r���W�b��f�Ib��}��D���\ex�.�j��婙�e�S�$�u������h�۔��ED��Gb�M:`��|�0���Q4�"���a�XQ�_K9H���y��(������au�Ș���%`����/��8kU�|�:b>���!�1�>?w����)v.dp��z F��}c��}n?�q�ڊ}�!��YE�K�k�È-!o�C�+">�r��n?�l��� |m���7���>Z�f��v���W��	�.L�(��@kJE�ez�XIג��!τ�g�S�nw�pJ(���@��޾�aO�x���'�I����wBaG��(�8t�s�C)\8,�-��A:;˭���%�coiU�8bP.{bw(���W�Lnu��֙F��nz��0�]z��v�fMkf�4͝�Z�_;\B����,� �C�T�@=�I���J����������f�c0T�2�����f�=�[}�]�y᜿7�Gy��g�ɘ����@��� ~8ANν�
�mDN��KC��:����Ҝɤ�͆��#���>��)���)��]^�b��� c�Iv��x�@�aj����򫓥5�Ѝ
%If���nh�R��;��W���R��` �Z����������w�a�Y�����}(���Y�yi}bӭU+���j;�,��Mᦰ�cE��=�[ǫ/Ay�P�I�O�Zo�.W��ԏK���:u�4{��y��z�OW
�m���\�Ĉ$#�nӡtf�V���;�m��b� �F��%��uow�S&^�q�>��<4��?�Xν�{6�@e��S���n�6xҫ�{�!�_V�{������^Y���	F���^:J�{!V*L���I�n��C�1���7j�����V��CJ��6>�
�|AnS�[��r��#X��y�ǳR�2�'�$12�ʜ5*3�� 2xUX0D�c�6���@r�/.�+����TbR0�sZ�j�agb��1��MRG�A�h�4��v���T~y�� f�k~���9mZ��W�
`Iu�Y��&�ٲ���L�I����<3X&{o���U�BV��Z;8�g�-(I;06��A���ܑ��fS= 9�
'Z�xUpFo�Ev��S5/�/��!�D�?:� K,(���4f�&<e�:�򑻴�XK�2���vR7uFA�X���"�(
��beyw������'������H���U� �H�.������9OM� 7�R�>��!?!巸���d˻Xډl�54���(	���ᯱZ��!m۔Rj���숄d��I����P�N�*���m�Z]^+��T�T.�3�c����g��������
�dbgA�ټ/�$�0�[�d"~Q�N9��NIp��?�5asZ>���@���W$2�t�Ľo�|V�h#KP:=&N���XA$z�>�a'
���Q9k�e���]1��l��F�s=�Z�(0m���ZW�����"5�:
b�.��%hcZ?@�^>iy�[E�z���UE1�	/�J��~ɢ�|�3&hzq.���ƖQ8S/`�:f����p�1I /��� �֘+v����W��Νv�8���G=f�X��G��嚠����fmɛJ;��淙RV�igv]hFG�+�L5@�����?=���K�l1�Br4�1w)[N���t�'m������}�{�M�U �ZM���L�zBw2���/H�����)e�#��ᔁɃ5Yub���]�3η����[� v+�(����~L/w�#+��,���pHl&����9gp������Z�+_;b��U�c���Wl�:���L�Նm�ա��M�з�I�RClϻ�� �s�8M���y�u��Wi�ag�.d�p�%'_5qE�b�s�(��U{�}H���U��sXT3hG�S',�A��<��3S%m��uMة��M�v*	P@Ÿ�S�}���{A�B3�����$����ϲ�s����Y�,�%�]��7S�3O-�T�
�:���J2};K�od)=����}J^�}����B�f&�rRa��H=�^�;��C��-ں!�K�G����4�?����7��_X���\45I��RX �!�?I�<���U�H����=��,	V���_?ީ�U��_�{c⁃͟�¡+=����&U�e�=z!��=������{N���:ǉ�L�%n	��\n��1-��m��Du�mv�>� �vYߩ����v9��q�� Cꆿ�k�r�g�s��F����!X�8F�N௵ ���8f{rb�TS��?M�	�=���{P~�vf!��t�S}�rzu$�����
�`Op���@a���GӢi_N�̢r ����^ad�����jp�׻!]�j�d�W��*l�=p5��2����i(��2�l%���i�[2ә�x���jb�Σ/� L���M��F��;6�h~�Qr�F�������b]?����`��P�f�:`ƣHN���'o�7_�`��3.��,�4������Q-)�ca�
���{v�wߛ!��q�j�xPp�ݩ��<����,W�7 B�Z&F9�Q��*�]�������У���/�S���u��}��,�\i�����[�
s����,���p�d�p�����`�[�E�{ݠ;+�{�͍�y B�6�������QӨ�A&���T�Hxr���p����:s��Ap��^|��;��B���:9��ø�v �=�����v����)%(iH�2	�E���7Ð�l�Y�͸�n�����筽;.+�G�rv�qt�ɓ�, �o1:F!p�%q��0��o� %�o����F�i�*�x�C�~��P��D_چU��6R�
�C/#I�˟��/l�c#S,��pz#�`[Jڕ�4t`$�R?V0���ZY�% �K�_tU`��j^t�(
(ve���^�:�:��cD�x�6I�~�*��N�E�y��'Bv�_�<힔�Y&���E,xB�>7�,��}%�R����Iz��!�tIX�iP��J���P��d<_Mx����<����R����A��N`�)��Kck�|Zn�P$�c�ЉXCp�������T���c��'K��ΰh ?���5��x�y��vZ��J�Z�̏ jɷt�%1q������O�kT���>(�l��m��98�L8��D_��_�9 SQ1E���\�չ\�20xJ:�!�d������L���Ѝ�g��]<�F���mA@���0��u�9�.�8��<X��iՁ���2\�li�IvC�8rŶA���S���]{|��z2(��%n��*F�h_�@�w�@�?4�郄5�s�2 ��@�y�T���}��5�[�[��:Lj�Sz�F.e��61���[h*�9�\��H�FM�Uj����t���b����n��b)1A9z�w��{� 7��y��EJ����t+��g�L�@�
Y�i��C�i�˜!/�{􌭜7����r�)���2�:��̉Y���F.TU3�� �4����~!UC�/e.� ��@GC	>:t]��H�pr[���N��Ήzo�+3�������,����_�����೺e�bA"*nfô��>�:ϛ��K�����3`C�3�@�̄���3#�������u&�#?}�ƍ���ܢ��G�d�,�
���L9@�Qu�)�G�.�E�>b�j�Y~�������z���c$/#�}뻦�kⰠ�v�h�zħ�UV�'���������9��+A�^ʅ���c�P�!\-��5�2��'aa��|5�?�Q[wiK8����G|	��@-�R���o��Td��%ͣB��;�o�(i#V�ۢ��*e��N(2ҿX���z7�.=xz�ϔv��̄]1k����.$���q����6��V�1Hb�z�+�(����ʁ~�ʴ)���!���(��w���h}�ϖ�GQ�q߾� 4��?��i��|U�i0W]�����f��~"0�v=��TF�چh�6>Sc�U���h�-7����<S��"�8d@���@8�ŷOrM�4Ʉ�����~r��p&i�&�����@���gV��M�?c��0�\s�ErV'��֒gңœ����3�8IU�tM:�n�!F���n�y5V!Z������d+����H�P�������a���±�5aYl�62�4�� �B/�9����ҝ�N�-���U_��s��c�o�N�]����f���\���HPk�]M��zk1�]�ZG��"�1I�����l�c`&E�>��V�-ifCV�G�N���U!���fLy �dn��7�����iFǵ ��ɳ�6S��$	6Ej���!S����a�l�Cx�D�g��X�t�,�j,�i/0�����Vz�����Al����vG�Y��d9�ܓ{d�1s&;���R\�L���ĺY�JhV{����"��?�w��ORf��Zd���QT���o+O�0ש����ٴ;�9�i����K. �#�mV>l1j�/��;���R�����:����X�ĉ-��,��md[M��be`N���}�%v�n(7�G;r�\�}�K`v-�������i秝�W�^��j��Z� +��wRA���1W2["Xl�i�LTD��\�W��I��8� ���P]'|�c6�U���ω#�Zs"ƲƆH���(�x"	��Э(_��|)�4�-���uv��H�sȞ�>B+&2gf�F�XQav�C=�qn�4��jk��ڒ^�.�+S�!~"�1��I[z>t�a^U���0�4I@����Ysq���7�L��Ǡ�k�LM�,�`y�{�$�+�O�<~.�%kZ%>
��?aY�i��xۛ�/.��C�(!'2gV��iQ�z�7	�S�@6�X�窷U��,��n�H�X�^�C\���Mb׿S�uup��0�S5�bAԑt�0xf%Uȅ�cP�CŚ�p��@B�[è�%��/�eW\��4m�loc�&�"3�O'!Y����;Q�Ϗ�k:N2~���
���=@�_6 �>n�]r0�:�fN���Z%Kl�sY��u��e���!'�!=�;�o�3��?aai�,Nwb6�B/GB����!��/�^A���tC�SOF�+�u0³X}��#�Rw�<��$�
iI0R]��%u�d��e� ���',��7�����|ٝ�&/�Xk\��|+�T���B�:��h�P���}���ut�C��~vYU�%��N��E�o������o73+,]�/�8梵�0��W�۩a!ӛ�ʵ��	�u�gPo~s�hAL�c?��Ͳr�>�A�@�0��n������/�Zrn])3�#d��+�q��߀��O���y�*�r���8Y�(�K�W����v��\Z��	nĘ�,�7T�[G�nڄN;��)r����Fg����yb���R�Ç��5�/�N�Ift��{�xj����_h�Aņ,
J�T=�Qb�Ġ���=�MM��w� �e�K|������m?)�F�g4Gյ�h[V�����-�9�y���YD�0?	K���d_��Κ��˲S�,w`$�@����R ����;�w]�`IT?"�D
�R�v@ �~�+i�8�JJ�� 	e?�Ǥ�J��E�%ơ��ۢ�Sk�M�� ����r.V����R���{�,F�\13ٷfw�0�d�K�hf4�y*Ĕj�JW+mW�+��B��(���?����>?@~�����-)]+����*��:�@�J*�m��s;����^T�$V���E�U�!O���� <M]�(�xo�v'�"q����V~��u��~*6���,�M-��LL&����[Q��Fy��[G:�� �/K�I8Vs��o���ɿ���1�-'�N1�8���ӵn��)�ɻ
�</W����bc�� 5_���t�O��?�Y�[vd��4mN�v���R��=k4(0&3E�e���k�^��qς��$%��Ȯ<����rC�8G��rm�^��� �F�]
l]�;���YG�h���楍�?�`ԖBYq�evjM gidhd
 QS}j�Y�ꚿ~�����V|؈P&���$�
ZBo��κ��n��SK��~��^�gP���/\�J�=��܌u���ޣ�X��a��	 hէ��^�������t�P�m���+7�k�>DsF��E9�n��5T�ݪZ�߫���&�3��:��W5�~C�C$&���x\R/BM�ʐ�)]5C���D���4�)�vE�q����V�����w�Ï��z�&��C�O:�:�8�Iǉ�" �'OS�v�S�����b����C#�VU " �S7TO����~��l�8� �UF���J��]��1ȘX*����i�[S�����e5>0�۴���Q:^--=X��h��(g�&3�R%M����Z��	U�H�L(��3(
�6���*�t r�\+6��0��d�9���K���SYd��ʮE��o���IU��!�g&����nⴹLd��NM&��BM>����y�sQ},�س��B�#���k�V�b��3���2������.�CiL��4$W�.n����Y�̒��!]�[��cب����֑ ���?����x�r��}Se['��7�X� �X�h+�ր�h���_���H�Hq�_�S���J-���P�L�-۾	�[��g������p��cG`��Qi�{}_}�����-�tk����W_�%%��� ���(5׮����n	e�;�b���2v��� ��4cn��.!fs:��֙Xy�)�˕ֵ�� 橠|�wYO�ў�fT��&�3Y�����a�}�H'���v�"&ʽ�ϕ��߻XN��l�<��O�W�$#�,;��g\U!��a�"7��ɀ��.��j����B�>��S�rXP+�Ac]���~z/@�Jp账%�P��LE����Ս��ʲ���|��R*��!��2�k�	��^�_�h��k�h�"��P��Jƙ�5�F�)C�l @�{�D��4�]��N��Ze��O��7 E�mV�د��2�̞42�YQ�;M����I�|��)sX��_}-v�������}�p�7������w&;�t�a��W��=D�B�aR����"��C!w�r�,�! �/�QH�Y%j�ս�ir���$�	�` !���	�{n�W9<s6�z�%�x�{{N�Y�w_�d7h(�ڕ:�L��A��r��ᅐ��C��藦��,ʟ�(��ղ/�MXh`���w V�CB�4�0��<($uf3E�+���{�ԇt��6z%Srj�!^��:�o��nq��{�][�
Nb���A|@��
��8C�^P��q�J�_1m{q��)DI�=�4��͈��A��?��Qw՜սJ�TՀ�@�%�y�e�ӵH��n���-��[m=w�ʚy��?�t1�G7S�g��O�2�Լ�,�J���O%�P&��-�]���bp�C�Y��q��e0��T��To�W!���2�z���I		R�D�IK��sJ^���+��0�2~"���'���A�L����Â� ����T.�h�+����
�ZX�e?�-\���:�0�S�1E�8zGӕ��މ��F�m_�V;�)�ϧ>a��?�[����qƔz9C��\��Dq�7@O��Z�k���龱����j�bq�O�"q�Z������=�He�K�K�:%^�%��z�FӶy����
!K*ҷEƉ1�N�������+���n�c��%� ���ms����z�>��'�E��+���x��^���4��sW�r�ډ�x�|��΄�C�4�?J��Z�0�����8Kۯ�N��
;�ܼ�9��(���I������P+w$s�!�v$.^���3����,��*z
�/h�쑧�{��$J��ծ�����#�_U#��e�`za�>�E�l�(��o�U&c&aF-��������+��rV�^J�A��7�9�D�&�x)W藌���ż.�9�T�哽؃���D�B}8y�7.�Yz隄��ՠ����-��r�RQ2K�Lf+JI�I��gM�̅Lb�Y��90���*�[��#�����l�SЭ�����PZ��_a�����נ/}/1kN���m�e��=�'L�-I���	���X#���q���暣�#�*!1፛;QgL-���t���\����Or��0��FsɘDg"����6�A^��[Nu��Iv�(l�U/Z�1�!d�S�N������m]�Y�&4�b9���Wp�^�G���I�C�$)�ۉ=�+���ehmDD�:�M4�Ծ�;���~������@��뾏Eu!�:>�)&M�Q���g�K���L���U���ΰ�w+�.��!�V�����	��n��~�"��.�!9��H"�H�Z�W�&��MZ^n�&�'�y��ų�bT�����d�T�$��e�����}���(g����5[y��!"�z����k�À��u?g_)��υ������,1�79�G���j�p���]r���-K=�͇�~�b�oİ*R���'��YU���(t�z���_�wb�j�`�����Y��E&���o�����&Mi|�quT�8�dC��<�;H�G��nk���0����Io\���z�ˀ'����L�I��$��>H��ޢ+�����{z�����]�R�c�SO� �X��]�Tk}�O<����-�Ƶ�(���:.�q�\Pf4�4�P�V#͍KTy/o�G��7��M��8þ��y���0�`�A�[j���;I)s.��5z*T��ɾ@-g���(�[��µ�a�V�����<�E������w�Uo�/|��`�5f���;F��\�s��l�t���%����A�%���}5{���� �jP�� �z��~&�����p�rVޕ���t����ڱ�?JS�����	z�V����.po�R�.���6Y�M�������"����\Y�z�2�̤��N�LC��F�v��KF��-RtP 4�������'�y�#U�m�x�ꋻ`����Q��C�I�\��D�xT~��sQCكW_ʰ-�sst�}��a�c�RG��[ ��K݊Z���U�8�Ǆ��$�LSl�I��'7�߰!aM��k��2�Bs��M����Xxl�	w/��Non��ؔI�2�w,��iPG��;���$M�X�	u�����l"vN�&�%����1l�f(c��jm�4��:�]Zd��g��]�~�=�O�8�`7.�w�Kd�i����zY�r�$̜��?��S��{��&ٳ+U�u���l�uP�BZ��qu�$�9|��*��){DИ��c"�.=�ifV��@"����%�V�J��*��<����^{_F�{dS��("ok����.h�3+����
���|�3@!�\dߙ����G�_������5«	�)R��l�/��S��PzS���W�1�����&��ﳧ5�w�u��غch���#9���6R��ؠ��d����-����Aq�w�|�U$���_*@�n�#��FqX�U;��9��2n�\�r�'�����]� _qU��l��/)�gw��1r�e�nՑ��t���s �,k�!ʝ]\ެ(sAc�gqR���?�@�iQN�"j�������P���7��j�B+01���r���KYx��0�����&�6S���Q���1�(��up iۿѵ�h�gE��U�%��6�%������˚��*�&ӣ;,.��/�#��Z�3�W�
�x`z٣5)g����w:���qDm��K[��j�+�jI� ��Z���A;"��W�5��E<�6�[E�.`�`*����<��S�ZvY�w�<���mA��i]Nxm��%@�~~�ρB��㓽- �ȠSx�X�i��hi�\Ik�)(���4ь|�i^
=N�;�O���=+�O�N�7 ��7��Kl|��v���>zi���}}��o�H#�ñ]��T�����?�3=`;Cd��mm����~>*L�%
a.�z���M��z���Hb��)b��r���$������J�V�r�SU��-
P
�|�'0~��d�����m�N+��^����;BQ*+60�LKڵlo�}]#�۳��/f��iϡY��\�~��W}b��)ޔ�0B��;��ubElx��ݺ��V�$���ɪ�P޿6`�Mc`�`�Ny�~�rgr�F�އ"��2��9�1���l������2���{t�i:��s�Oi`�~g���i��4��)��
�o��[%ڑ������Z���E��8Y����(�!�и�J�8�{k�{2]�����5�|77ǜ\cȈ��l�a�i��~+G�sm8s���r���L_�«1%��}	=|#&-��okN�3M1�.�hpM���U�D�z�2u���p\C�fW?Ӯy�Ҽ��'m�O���J氄S��퀏H(IKDvH�eO_۟#��n�t���p��׳��ܽ���H�CS��s����E��Ct��Pg���*q��U�+���O
�ϥ��.��(��w�Ӳ;Uc�S��q@��������ٜI҈c��>�Q�t5�leB��ʁ�Ut�9w7h�P�k�[�lu��I��Ϭn���n��������0G5D:yz��U�@���^�>{7��6.��js�F�D�}�R:ToU�C��,���(g�qK�n�q��u�\5ۘ@ ��dʷ�=����g%����d:ɏ!������;ȴ����Oh���C޽�ΛIߞ~��.������^ud\�ڛ�k��5'�46g]!B���	;��+07��ؽ���b-뺗�[.ww�@.�ߍ��G(s�'��T
�y�;�vz�tYY#��Gg�;ߚ#�5l~P�<D���[��x��ǟ�Щ¢^M���!OR�d `0���#n���g���`���5Eg�#F�~˧ 0�\�^fqHSn���~�]#%�Vb�B�g�5���9)G
�kE�]w(Wz�r��]��Gu���-\/�z=Z�+M��o�Imԅ�%�J,bTi���=��ؽ�����4���3C���.�HS���; �1����Y���ӆx�Xo�ǐ�vd*Bx�^#��-[g��n#���������Q��lE�i.��w�-�Y�X�Ǡã��`�5��K��ČD����o�v�C���fPL�rai�~V�z�8�\�H̃��7e��Y���Aˌ�H3CPvNw���ܦ��Qy(b����R,�C�79�=C��ί�\{�ʯO�)%9��F�/aG�2@O$o��BG�oB�>���'&�@�1��7���/�/")�$.�j���Ya����P�Nk����
���tr��)~����!t5���z�*+�Ry�f��[�̗�'��Ze���f.����eQ�@��Ӂ�zw��i�]��X��f��פ#q�Hu���W��U�::�K�Ӗ����T|�Ƴ�#�ӓ+!Y�9�S�����c����F�z~���ݳ�܎�sjO2�,~nQh�K̻��O�Ό�#��G �t#(j^�{��2�����)� �b�AUi���l�_�[캓Մ&�)'*��X�Z��ۭ�A�]���î���c�c<�_���0����P8��a����3�lG[O�t�Y<��0^[g�&��9u��h��3�Mr)���k�BZ}Go�(h����#η�_��;�V��ۈ��D
V��)�*��U��Bd�%"��K[��Pa��õ����l��!�7�+��u����I�j��q�]�d��I�po�32�C�W]9�wiׯ��98��?w
ۗ�Y��@��U�ˤ˝�q��sp�����U��ܺu6�]�p�����'qr|D�V�.��7��� �_�#v��1*�D)&��ᩛًlÞ��i͒T-�X.��dZ+�"��+�}�xu3IC2'��$tS�H�fk�7�c]������a���[�/`�$�0��󥊝e�Z�XELQW�D��6�x����+�>9Qd�Dg���}�&��~�9m�9����W�E
�������i��J"EV���Z�~'����^��8���_1�G���P+V5�T�x�� �:G�3���8��nd5#�eDm��=�\� M���D�S͖5����Txޚ@4gӊ�2�̢\~�Pj�0�ΐ�Gf��a���r����by
u/�����h}icV�d�>�uEo�IL(f�+^6�߈=�g2���_���꣠��%�e�rg���������z�zDچգ�˫�z�$u�'��DkGBçu���v*�~ـ�<��1��pQ�_XF��P�B�=����Xp{���ڱF��n�I%��[����
�p9�*���J���0������=�d\���%�n����Kk��H�!�����˛rew,3H$�2W\K�&�nK��f����i�%�cڍ�lG}��*�c�H+� 6Z;;3E�����l$�8y��v���,Ң�>��d����o4p��p��h�;`��7fM�tCԃ�j���ȑ؄���>G�(��Fc���� ��Hx�F����w)_��S�l���}+���XO��z��Be
+�v���s���[�Ms̷d(�1esҒH�%qM���wZ�v�ş�uOTkx�����dM�sn��T��K�&R�3p4֘uj�,� �ы�t����{h��q:;{6�pV�4h<h�sc�s⃟"���U��R��: CXF�7z�+^Cp�P/�$|�&AeB�o:�*j�w�=�YS�yb\�W	���7p:M�̂
�ۑ")/pDD(ͪO�4����Ӄ!y��8��0���GxE���]�5�$���C�1��Ŭw"6�y+�e����"�_��NA���44�M1^y<m0�<w�6N�F��b��5��=�F�=�#dc��Z�%	4���Q��X�kG����2>���2ߔ���qend�͇tCNm��]E2����¶�*�\_��:�C���P���
����{�g����p(0�/�F�Y����6�?�D(���ߪ񿛙@ ��0���g��k�N�z��jz�ࢹ�z�en����\kJ�n�sN��IsV���um\�G{�y�>�Srh�� e#�&[uf��vV�<?4)�3a��S>��}8�V��T�}s�l,�7�g�x��%u�������B8燮"ǻ[��]F*���o�o����^��][�
G��������]m_k&�������0��u�(TH�Ŵ䬾�@toc��(�)Q�H�ٸ�E��6�U$2h!�5-��Jk �zX�� ��~V��&Uf >�Wdhk�K��sh&�E
z3��tH�}�
��_Nq~JeNR�kߵN%���f����	(�yi�?J	��_��tp�i%9#X�o��I�Dϩmm,�:��.�&�2���]x�����oA���S�6����T�������\yB5\65>O��ۧ��^��Bl�e?�����M�4`�kT�T�s�������}��Ӆ�g�{9Vo����4��B��Qұ�D�#:��[#тv������z��Ȏ&�S�ڝ4Ey��AO�AƍZ��r�� �P�"��=�F����%��9��H�\�����e3�O����3.	�6ZA-�8n7�=�@B�YuX#�<l��7����[s8@�b�Ÿ$�IEA� ��x�4���+cZR���i�C���E�"�]Ύ���Q�ia���[����(��We�O\��sǶ���ȣ?�*
�9��fD�@Q7"���� lz�Z�����Ɔ��]B�m�i_��v.i}�Pg�b�Aھm�h���b&.�uђY�L�z�J���:�n�ߟ��Op�"�i^��Կ�"�x�CJ?�AF`�gm�%�{���:�\)0�Q>������L2��_�EĹA�JN���j{��N�H*u��*W�����	����x�a���0��'=t�cD���~�n��둴ю�v�T//
V�,	y)�I2��ս���O������B__�bh,rp�>�y�܊���E{��"QOTI�A��K����֡|Ѳ
3��DD��m��� (&\OQ�J�49��V�VG���@��=./�YtX��w�D�;��E"�6����m�����#�xE\�o���G�se���#P��F�)v�گ�V�) Օ�*���L�9���~��qsP���u�0;xGz�Y`8|��=�#/q��7����0��E���7ӫX�h�-pHWt�N�\��)�i<�@��S�$����.��.�D �7{j��ŝ�-H���+f������\6��2�qVE�Ď�K;�ͥ��� ���\M����z�y<X�L [��=�����C#�=����q�aS=#�y�d��e.}j��XLd+����=�����Gca^�m�������6pEA@n��%A]%Õ��r�=3�Iz'!��M��o�b��wĶ���2�= ���Ui�(��᰼������0�=���l&Έ8���vU2�E�]���[��ƬV��Ta@ns�
��zP�j�U{'fi6���2rq����˜�P�� ��T���t��'�_�8D:Z+K-By��ݩ.�5ښ�Y��p�L��#��ڍZk�m=ȅ����n����]����Q8�YT���+��$	-�V�V�4�)�e���r-�#r�n2�/`�1f�e "��5
4�͈�.SP��J��n&���:6�� �*�O�|N!0� ������+��<�>���M!��A%��(I.�Qp�X��A并����,!F����}�A�g�����L��Y�@:��b�3�X)�-�cKM��߱��R��T��(!���D#Q4�L��}.^kC���(�Vǔ<7P���zzp'>]�%��`H{�C� 8{π�.�?��8����yag�)�H��h,S�����J}d��΋�Fh4�s�H|�<؈�q)ю��]�K�D��,R U��� �a9��1F��^�qu�r[���t^���`�����z��0)�L�|	�ޞ��y�Yِ���}�������6uK�a���-,1��f㥥�\�V��]G��5 9s���&�;��F�`&�Ծ��\��+|<�cEӵ����}�G[�t��V+P���~�o����#MW_�9�F��<9n�A=V�G	�e�E\�@�WuW@$4��\��K�
f�N�\�6�X��z�Y#�%�e���v�Aw�=ǴC�a�&�<P�y�/̋0~�	�u��i)k��8��<���N'A��B�b�-����ɘ�T3Y��JB�mYY�sq�l��62�ck�Ȕ������_U�����ɉ����0\KU�,���ϯ������o��~!ș!�L;�9IC_�Rb%��y�Fo�+^6��K�:'Z��Y�`]�믈3�-�"3�G��-��V:�iX�Q(9u�P�8J�_���iCk�i�H=~
!>S��=�-'�dqʑ�#��ps:�1��D5Չ�K�QL������C�/#�Uo=;�F�u���+$�Z��Y���}���8:z��?��o���%��\�$��Z��	؋�W/��9P
1�r%A�H��i�)�a�ӣ�60�����L2)����RcAeD�������ð�NC�ب�Rg���?�����5q����vS��^����3����h�+H۔+��J��J8_��bg�u��Xf9N8����>�� ҿgVRHE��w�{�G�a�:��1��:PL
�F�\��k�˛J�&�D�M��@�PPagH��	eBl��:��k��`h����d��7����% �]n�ܝC�	��sh�<��ZA�
Q���+P_�����]:��W%�l:����������"im�F�2=-.&�vQ�[!�����*v�èM�v������J�^�^�P�q�2�fC���I�X���@����?��~
�q�Z1��3�θ���Y'�Y��Gm���������H�0�}~��j&�A�C�� ��q�QBʞ�8�pa*�K����V\�Y��`���z��װmMfPM��� ������W��q"�֏f�)|��6�`�UC%Q�yO�(���z��7���@���p��ji���������|��d�d��f�*Z���J_G��~42U���#�x��%�p�Z;IN���b�t3.���� N��n�6@�e5i�<���L����/�_��oU�����N4Z7n�	�q�|e���$fXߘ�bʪ��S���&�pn��@{�&~��V�㴍�z>=��禋�U��r��/�K?��x�G�mO���e�Z�=��q�WYoH�ni�z�����w,��,)��{N;|���.e����l&!m�� @`���IR���w��}�'�盠�=?ؾ�WJ�q��׿��t-L��p���`+(!퟾!����#lq��U�_S�y&I�p��>�B�B���u˶6��*�r&��
����2�vKl���N���`��%۔A��x�ծ�������\y�m�!�ҵ=��H�.L@g�� <F�b&�l� �&n����~�3�P�v�%��6ĥե�O%����St��-���>��l;��20-&�~:��K4ۑG�����h�h��H ���Irq$����W^ئP:"�3]VDPEH��\ߓAf�[�n94Y+�l�c��uٝ!*���+�iy�ŇxЪ��ns���T6�[��ud�����}�ܤ�P�0�y�Ǌ�{L>ޭ�����8}�.���̂|��q�n� �"��젂�,N���)<76¦ē��(^�1(zi����E�	K�P��f��8*MX7�mO��0��,��RY�y��Mi ���;#�\��C��-b�Hf��x�x���h���ȵƞ@�R��M{֞��.��q%F��m��on��a��RD��]�1��4�������GZq�@�EP��%594��4�g�n�=tݻ;��^q�レGX/k��O����9,��#x�˒�n�wו���3�Vcư�O��M<#�J���k`/0�.���`�u��i�����4�zB������n[^e0�bC�����$9ZU;Y�yPh�d�q��c���+�v���8�]be�N��l��Ɗ+�AH�!?�U tk��(�<L�}�r,�ȏBg���D� �!�d�F:���?�u�s�:��z�� �@���~'D?A�j�׶�	&l�j��ǟh���X� ��F�� `+ő�$��D0g?L������ cЦr��X�u�!u�工������ed9x`Ym/9�s\�E�(g�j*�gݞБn��\��D�ڙ���4c9�uI�4"���Do��c&�#?��YE�o�^��FU���!%��j]�+���֒Gg�BR�E���Ҩ|"�+s�O%<$�wPDD��H����y��8;���&�l��H��ׯ�4oH t[���A�*����	�=�^�<���농0Q�rH�	�(4y�^��m��eӲ�.��e����2H��hS.�PǤk�� �K[1��Ea�(C,�14��.����[1`�]��݁9�F11IE�}��b�����w�0Z�=OFNu�x�J*t�B<k{r���7������sG��o)�Ws@3����#n�Z@V5��A2��;csX�9YD�VU�tY�"2���4�l˻F���αB�)��rf���C�^����@,��k�oX�1~�g����:�+0�$�3��=�v��~~�vG ��*��A��)�*�����j���[,�`w��s��No�m+����˗����
L��ql~C(��'��u�N~��߳��6�TN����9��F�7h��m���?,�%�,�L�S��:��Cج��G�OJs&t�}Å娀v�m��A���轁���E������\#�}]u.����h?{�s+CZ�C"�#�rm���f���"��_�(�g�;.�����Z>���V^j�6C�m��P�)qF�f��|4��m/�I@�*�{��>Rt��N��hM��.g[�q��h�F�$n21�!����S�`TP�!���1���@q}�V'�Zt!���9Ȑ��1*�>�'��᩶��[tR@@�?�T�����ކ��V&�'~����� k���_p��ǝ���,c#*����6
&W�<ͥ�&���i�|yѽ}ec��G��-��pi�T�K��eJ����N�\&(>�K).9W��(������F	|M�d�)�ԳJ* ��
�&�r�� �q�tÄ�Y:���v�^�]ӗ��|j";J=()�`�x�l��d��UHl�����d�j]�t�0�m���a J7�#`Z!�f�q#rڢ�����	���n�pl��B��gP-{���_�aˢ��Ɓ�gHI�' ���1���.�H+c�"��%q *t��"\k%�|[�ϞH\@�]t{�I��A��]��N�;G+�=%9u�T�E�n��}z��3�i�S�D�D�}�3�<Ry�� <�蹄�׎N�x,=׺RD:�P��1p�宑����v9ᬠ�k�-��7�wr�Wg�����v�b�zD�9\?g�D,<�U��J<E��%r Ë ڼ�9/fE���v췪��!IB븤ӂ��{�a��W�h��M��M�M��7�TA��������ƾ݌Z���
�v24��4����[�%13���x�n1QJ�N+��b�Qy����M"ӯ��Y�߄p�g�"��0�>��?<� �E�U{\���!7���R����jDkl�\�m|�SOs�F�Ȳ���9��`+��:�����9���Ǻ��Oח����%3��k�1�e<3U�fj$�dp��j�bug�u��]��qya��O��H���Lmj�ԝ� �(�/
R��0���6Lz	|7���@W��j�?���
�)b�C���
g��g�+�z�
�0>֔w�R�rp���(n5."쳀-,��"j�N�J�tmZ��_��v_�\�#��w����C¼��n��%hI~����L�ϴ��M�!yR)A�_��T�`^<+0���P�t��K���`����Z�	S_k/�w��ʛs��dMW�:DB�#�s����07��y ��p�$Hm�����H��ڐ��>�o~��^4mm]�M�;�h[�����M��3�i�d���v��~�a��B_3��P�F�K��a��̢������'q�)��lן� �jLR>�GTޭ(n�H-��L&r�]���t�j��r���<�^�X�M�7�������%���~�s�>A8���t�7	�ܷE��N��#���%�+[���R����Xh�)��A�m}�vة4�?�(k���� � 8��c��:�be�g�ʖ2���]G�* �"���s�ѽtY�fUW��I���6���+�g�8��f}�&���k��[�d�0�I{:b��1��l�#�,��R���OKf����!r��S���Jxnq����S�?�s��sŜ�RũHa]�x ���f��.�V3�2��K+cI'%�ީ6�L��h����O��fJʽuSr'B���vN�U�����!W����qG-膢���T�L��C|����, h��O4W�A���&���nf�9��:&I׹Zx_�Vr�=昬��ٚ���bf�l[ZAyh�&�e1��Oj�숣���4����8������$ �E��d�:�>�F'�2	Z�F�����¹FE.��'�۠��0�+���2�mE��)��<��x�9�/Hi,����
���[��E�&��';�Z=��h��)���W���H>����FT=��2�0��pL���}/�3�]�o����I��=Q.;���]x�oW��<���!�`��IQ�v�T��$��W�{|�;=.�է�|X\$�kV�d����c|���J��#PnȒk�^�|ȘI��q6#]/�a�#���{R�2=Azz�\9�#/)���Ȟb�`p��+i�T����S՜*N�������|��M�}�f��	h޿��I_.�v�E!�g�g�:�t:F�Y[��]�Y�����2�E{{'�E�d���n�̴-�k����pX�[j�y[l���8إ	>OS����e}!
��w9&�e���;@(Β6�O �_8v�m��MqPeg+��ۀ*;Wq�^=����8�C6"���@KF�aM|3*�>eBK'��Q5`�j���2� �o��E�X�!\�p_���"cR����p�����a%E�i��'���<�������V�w�c�&g�|	�Dw��	Z�����}��7n��t3��m����#9���s�O�jB�N����f]$nE�!�E��z�,��F7�N*���.P���]�����cM�*���i��?|�X9u��hI�uj�m�$���&����;_��:[]L�Yh#��[|��b�,Xiem;�1D!g�us1rtۇ/\��dt30�}�J��� <���������&��������JA-��T���� ܪ�*V�PT�y�;��'��q�{�0�n���g�ݜ�d&��zL�D�Y��l�iɌj�Po�5�C�����C �u7�h�(�[�����!`'+��YV	�C��]��:��e]�!���G�J6�fJS�e-UGͮT�����,�㻩���W�q�?�W�1�K�0�YӖ���g�߉OE�`�9��_*Xo�T��B�r7��~à4L*]��_�H��mO5&O	�\9o��m��a��'P�hF-����u9d)Ȫ�x�b�	�l�ϹY��KiA���z)�A��,��H�b��� 0�ھ�6ɜo�悧�������t0Ԣ�B��{�^���j��W��os�Yr�P�$)�cS�ĿU���T�ե��/@�KdMi���S��$������\ P]�QMq�-6?�k^s�g�>�
����X�K�)���]4qC� �����s��0������p�:D̼�0檌��\T"�8��ț:G�Jy1dI�b�M)�;���r��J��o���j�!��� ��jV�B��C����Q�}�����=776<`��w!�Du?}�����cox�N\(����eA�(�U����}��t4��<�n<>�B�L�
���e��k9��@��Ђ�e1�'�l�l:��=�
}�t�#��9����X$���ぱ���^`��7r}��
�ܭB:�u*5��l�� =�)}qF�L(�����udWu���v�� xClܘ0�-P#<�E����˛����.�=`_]���E'kЎZ@=w*?��I�� �R�ՍMAI�\S���a���(g��u��_�oӳ�ql�:D�$=���4G����N����Hp�*�i��p�=��p�l���A~���oa�V�}L�R�}�Ap;��f;�x��D	���n�.#��B���]�A���\i�5S:��^�-���h��$��7r��7���F{�Hr�D����,�#:�O��i���t���M��̓�=>�5\z�\%z�^ʺsM�d�q��#�k�āA��%.���0sfDe*�äo��")Pػ�ڐ����$��d���c5F�.*|`�����N�-�3���ӂ��b���F6teT~�6�=H������Ćr�P�,�9�<="�( Ì�)��"�'����}2Zze{�z�� �/�O������-�x�ȥ��}5�
y� IU?�5�sq|>��0Ej]{���J +�'c���ݳ����:d��-4���^�/�w���e:���Î9k5 �L���E<D(9�C��H�7����U������a���yW�����Ms�2��x�>�I��Ėa��J�� 2�c�ñ��Æ��v/�\���1e����{�]2޹1&>Ʌu�3˽�B"�������fq(�΁7�$U�;K�H�iW��Yd���.'׎�����ܺm�9I�u�{��k�'�u_�}��A=}N`C����`΍#W��5�j�oDI���v����XV3m8w���9���h�1�"�2�I��'��@0�"4����d�6��_�xF3�.�C3�}�'�ٷ����E6��;��Q썤=�DI��y�@�cR��Ӟk?�ċ�< �}�q�lTl��m��`E}*���ѣpHz��pbI��'��Jۇ�K��n ��'�څ١��ܯ�ڣ�O��0�I,o00�v�Ok��i$�Y��n���i��A���pC���̗�o��{Z�|61z6�Pb�N_C�f&@X���]�紺Z�
7~]L�a߭�P3G=�P&���L��$AOӣ����f	���l:���g_iC�'4hwi��ɀUs1�ڼ�A��ؐX���ެ��*�r��]�����%�/�!B�R�]���l�:����c��͋$�tC��]y뢾K!�յx8���@��HP�����q��svt��7HS��d���_�t��RM]���o>���G�ъ���e�p��{o�yx&\`<�!Y��o�R|���a�r[ �Z�#B�:k%��fK��	�29����1��]<�}�,�nzKp
^�tV�z�
cd-*��0Gi����\c�hí����o
�#��xB��[���!�D�_&���}^T�_����f;�@'���
�!lA���;L6�#"�y�
"�^��DN}��x�kD2(( ��ꏰ�����0T3YM��lGV�;��ĞJt|}ǍĒo�� ��޴��a5d-���S	B5~[�5b}Um~
�ɟ� s(5���l �����k��,��M��?�%���D`s@��F̡���HQ}��c$��#�O�?����sl��I+%�7>_/)�ns�6����#S�{2_{C,-��]��9�o��q�z� �
<5&"��׽[���t��7�����.\p��?y��)���-�ԉ�ӄRV��q�ͷ�;��^*D���e���Gel��^;i|��|�(�9�߻���)z�<막ק	ͤvAmS�W[t�24�F��͓����}M��9�e$�*��D��GifMм^���~���}���x_� ىͯ��G���[�_l{���?H���L�A��q����ҮvUE��X��B>���ԟ� u)�paH��񉑪��v��p4^Ue����uX[��_��WΨ��]+�<ߓ/���B֠���=��J�Ǡ�c�)�k��0G��맼wj�&�١u3TQ�s�zV|�����.��5���	H@\"#����SHx��p#F.���$�
����&�M�y#�z`,.ݫ �����w��U���8�d\�d8;�3��H��� ���u?�8:��,�i�D�C$[@���w�2��_"�e۹
vQr&t�8-2Z�+��p�:M�U*�3�9O�]��i5e�X����'��4"����?k��Sjp@�6��.��jlհ�&ޖe��%b� i)U8G.�=J�&X���p��BӞ�v��	�Tد�u�2�<̩uI[��+զd��Y	���{�Z8��fz���� �/b�4.��ֈq<E�=:b'�R�!�a�wG���
�9���r�>�`�*��%: H��r�#��$�j�����ЬX/��yw֦�Dj���qq�O�A4���d
���ð�ʯǍ�8��)�����ߓl����������;�E�$����;���!��4�A���`�-����2� �,� =Įa#��CK�#*���{�戠d&^���m���TV���0X�(*T�$^�����bf���������A���=i�����=tk�æ��h�O_�I�U���)B�9k&��	���@�Aɟ��TO�����o��3v��7ݴ���%�|����Ϻ�������C,Cټ��6"��>ک��z0�=	�/7�G��͕*"ho��h �X��E��j��&�?S;w�H�p�6�����]�M�[�]&����w/쾼@y#�̇a��-~�L$p��3��_ӝ��YL��T�h4dI���J��e	b��$6��x�4v86K<S#����a~����8�Z���;�^Ԛ��i�yС�����!R�@���j���u�LU�) ~t��3m^�&ħ�Kာ�t)*�,HtO����j���.����K�u��ŧ��wNJ��u&w���]J*�J�0��)ѫ>^]y�*�?*@��l�oT��.2ٛ��`3^vQ�6�9yS)���P_�\�>gq8�l�9�8�RI7SO��A\W���9����%���M7�@8R�j���ӷ[^�Gw���S��{�^�	� �/[�j4�ګ\KI_��n8S#D�LB��G�v,2_W��T;�`:9M���_�]��`,ޒ���*&ү�z9?��}��q"`�fN���]w=%�D���P �R� n�N3�C�&v&8j��`�lG?�Ӈ��j+uig���e_b��7�\�0du2��C���A�]}��T�*����H���]n|(�3�L+y���_��=ĺ6HB�ꦤ�����q�_g�$R��xk����y�����hl��J�}#�bpa�M�$���$�c`9_�����f�4�(d�D,�	���(M.�s��h-:;�#�O�L`���L�j�֟��Wq@������)�F�3��q�yE�������i���]݂�c/�V�7Oʹ��T)g6S:��K~
�����V#�բ�dJ���s�9���-��K����Z#M��vm�R��c t���8��Ac;���Ć����H�aM��$9�)� ��EY�WR�p�Ų{s��$c�Q�Z7�����1�}�+���������}y�.˩�W��$?�+���5ߠ/0/�l�D	��w�UQ��^nv��JA��3�#��E�`K�������d��5��{C������V"oR�2��󅦆�WV��p���)!�-���U�6��~�)5[�ǔi���[�F������MAoDƾֶ�Ȱ��P���4uHDG�1�K�l�dh��#5or��m���N�����dY��dn�XkW˳���]"ӈ�p��z�e+>�j������h�Mث~v�����Hu��R� B���s=�C#� 9F��CG�X�� ��]}������uT�=�\���-UR����k�����&�� 58�B���A�%�~�&�zn�_ �����{�A�r�=Lx��i��Y ~�Զ�f�G����e=�F�/�[e��͹ρ�C
0>t�aIHl?x8)�(V�d��"�s{"�4�v�⪢��S#c.Z>���9�aJ�}���d^8��Bbm_E��2k"���ha��K���Y�K&�eL����
A��G@F' �QTd\:eW���|UeSN��'�~��2{�oc�l�p��O®>�B�$͘�n�9�\J�̋Vl$�{7N�Y�ݦ�z&����<6Sd�_F�)�❆)�}d��_?�T� %_f�����͆�ۿ<��]���}������a�����������RT������3�NC~>�"!�v�BG޾�7�V��EG�	�eW��xU�er��ǆ��ANC�F���\F��Hv�C_{*MP��H3Զ�5���Ll�K�A�����a��hQ�vK�2�q�I&5�H��
��/6��0���;�Ϩ��ė�.��0�ո�o����m d�4T7��%�OIs�ܖ����
YOd5;.U�=��݃K��k���1ښ�pޥ����_�F���S��R�]�)'��QU��Q�j����u�5�\δW0�,�qn?���d��J�x�5��!Z�uw.5&�p�hʒR'p��`�KX�x��Ot��< y���&֯ɗ[.õ����d�C��v�C݂q�$z�����&�GZ(�U�ᵝ����<F��D��fN>Nm�D���` l
0���t'��q(TѴ���[�;� *kP�@�v6(���׫��z5_3��^��U%��~��P|w�Y�
�$��G��xA����!�B�������5O���
ʻn���u�I��EN�ɒ��������.�Fܥ��ҫ�J�d���;��!mu�~&+$Mn�lE����`�V�!���dt�P�������l��"�DqJ�f�l	�-W�=�jR]�E�md �nc2w�si��^�hH�$~:5(�Nd��{a�6��(oݤ��eڕ8����i�U{j��*��vB�m��LqD����3�,�ϼ��7Wv.����&>'����Z�%ݗ��[b�q�e� ѹ6���!5�����	��:]�����o�?B/
�b��%�ퟝFw���BA��>�t��48��t�(~�Փ��2nC8��~�w�I�C�O�$1Dr��hMF[��xv��l��d���V����-rb��\�����R���I(�'4�p[ӷ3�� ɢ��cJ4R����*6��AZ1��¬�� ���z^�T: �RI��N߸�@�!����=c��R��Sh�����BVp�ȭdI�����^�p��}}���Rq�p�y%�玮�����!�,2d�^�;�5��&�J�t��9�
N�����f���rED��+���m��C-<�X�)FϦh!���n��k�K,�M��q�,�$�WCF��g\��;��I�@��F��S��pYb��Vnq���۱|��N)���.����L�p.47�[�u����;;3>����X��$|Uzb3l6�m����,�xB~T�8*l�lR X�a�hbɡGۼ�'A��� ��U5]u'���4ݳC:$~HvcG�
-'\=���R�(�x�M�	�<o��#�k�pq�n������3�=1��S&U7Y����s@�~�l��� �B�5f �J��8��#+J��@�!�y@���[d��;ğ:�ʏ�~�@�5S�/LW�r��f�D�j!,b�T�3�|:���"<%'-@����
x!Gjo ���~�|���%?� e ����I��?@
���>_��s��s"�F�2���/�.���B_��%}aGӁ��	1��O4�S���Q�zs����K�ȇ�������;�8+�3f�X��R寲Z�ܗ[a���U#��'��k�Κ$J���p�Џ�i�	���w���/�i3T� t��i��̒��קM>?��N"dg��\K���^�/�����8��bI�u�9�n��æ
��K����D�H�
�|�=p/��A�Q��
G;���safj�I��xO�]gi��ߕ����>�=%�JU� N!)��].O@4
�b�	k�U@v��>�e�5���0'4�R�@�T?+��ϫ�s:U{ ��U�zc��]�.kt�ƿ\?r�y@�/asD�a�����6��i�G�QD��q�W�@�C�v��b��7g�/ׁ�m����i�m�%?�c'�P�]ԡr�Z
������h�Lg]P6�����hB2d�<4�c�A�TY�r۠���M	���O{DD4{S���Uu�樍X�
��A�d�oO� �;���%6'�VX���y�"�yllP�jM���cw菳��-l ��$�U8���%|��V�媄�����Xx⼝�=�����l�6��r���o*Z�\��H1�l�>��")F��P�hg El{>ﺸ*7�A���C�5�si)&o1��c�ue䞽\���>*��{��8�V5ܑo�.[�,�450�C�QWyPP*����E�g��u������༼\K �ЄЍI�I ��a���3DޥO#���D�p~?k��0v�K$w���_�F���C����eGk����v!'�D�ۇ��>�ǫX��ZUD��QP�r$�jC����)պf*��M2ci.�D����lՓ� ��8#oT�RJ��˿��*�N�I�(���"\�;Hq��e82��|h��$�{:�#g�^
�Y%7q=���{%�s�"H���-u���E�aa�+����C8_�cPu'����v��YV��$�:����-���^l��Ll��eO8L)�x��c3�5(����q��D�(������Ϗ�+>� �䍼�q�@�a����\�4̑�-�3���T��tB�HG�t7�������~����㛶�@Lia�$kj^��0�����y1ܸ�
M��*_�Vk~����8�B���`�f��qKl�S������ƢS��/���/ ^�M%h����!��T������M@a��8��;!��pǀ���-���)�l�q'��"��4�c	*8&\��%+�}m�dLW��ةnvCdWjH`t���g.�8�UV�$yIXf����ws�Ƀ�D�N����=T,�����Y�:�L����1��m�Sg�$-~`�t�P���7]ґ�N�H�DB�a�+����8l�m%&GE�,PS|<�т@��J�+ow���L�:H{r�f�I�o},G�Em���~�Us����r}z!�"%2V �]�A10���=s%@���s��\�i~8.QFv�a:�S�n:&FZ\����uQ��$֫u(��iW7�E t܆sR�5�<uC����A����fSC���W5�:�S�t;H�gM�e6�8����D��X�b<Q{���1~7��{��j]��Y+fG��sK����ͩ��r���/O��Z}���i��ф��Rt�,5�e�Ӭ o@��i�Ƥ�
�u�vҡ�+�!������`��,�^�3`�;F�(�����{!�3u�	�C3k,��N�Z{B��<�L��z~`��}�| XE��(���iR��#��Ӎ��A���O�S�����.������9�4�gBWU�m�0͛[�!/�~��T@�(�|��K���m��r�sӐ|��i�����N� �V�C���9%�P�\Ng��-?��>�)����e��'2���N�s�1}q{����^����CE_��;�~�PN���"a��mv/q�T�=�� ָ����`d�4h����=�I�i��0ЉEW���\�(��3䠢awO���B��A={���K&���V(Th�7�>"���4dܝV�>TEM�Q`��e��0.5V�ޟ�X��o�\s[��OtRŶ����fJ �vPG���M_	&㟏 _�OH-J�О��| �Z�΁ '���?����8v��ߣ8d1WN���0�l����f⸸#�w ��4n��;o��ٮ�^%���8!�_ ��?Y��2uR�u.SU�*B��F��(��`��L#e�b���_���%8ѓx-�HA����!/c9����3n�L�!(�Xck.�U|����Q��?ɯ������ �x����'��ir��&��Cs1M)Ff����@˪�Ha��fJ�4��U�l��h2�#ʒ
2l2T�bb�P�>���/I~�U��0Jjѳ�6D;�϶�n�ꮞ�}M���a�SU�םX٭�͠V���b�|�K4+�F"#�B�]NϤY�ɋ��?-�6~��uRa���O�=�Zc�'t+���v��b�xQ��6���*eOS� ^�" �����Ȁ]�T�`�TX�W[���G����<}�qH�?�$j��{�n���	���Y�~Z8��Qs��@C
(ƛK�ц��/Y�BQ�gXYַ{3�H����[	��8��a�՝Gͤ{s�b��D��' U���P�tp�����N5��?`��1����.�T�s���[
b��w�;8Z�����c�������X�Y�&'��7����bq]�����dɈ��pH�\�2�Y�;3����G9.pD]��i�W�O
[M⥣\'Xov�wYS��O�1�% ��pi6�y{��0[�'Ґ� ��z���l����e�HKs�hx�'Ȓ�f�p�!aT�v���Md#��4 ��-*9:0͗2Cb��CQ�L��c�X�O�:)�����K�?0���g���f'�V��@�P�LN�*��=�H��?Δc������X��}4[1=�j{�-w"�"����8�=@a��#�Zs�,���z��Qx��8+-O�@�2�ڳ�Şud�u��)(���d�)u�a4�D��۔͇�|�2�{���,��L����:�D��`c7�N&Rw��_��o&���C�NW���0hT^o�&���t5A�W��r4��8GO;4��5�ջ��
DD�m�gSK��L�7�W�'w2�Җ-�g��]�JT�N�����-
��欈hUBd�G�L� ��h�0�zӥ����k�l�--���E�'��8,�A�)��$4C���zG�u�-L���G��D0������ )��hb�I�c�]~�0nt��t~e�ٳԴ���ED��H���_U�S�V�O{k ?�:3��n���ufWg[����J��3U�T ���v�������5�͊�����x�w%D��L$,�!3덾�GS2���P_fr>�o��~��'>��.e�=*Ɲ(�����"�sc��@�9�BA�lU� �)"9�C,�׀=�h��2n�o;��Z�V+�M�"L�?�gVM��� tSN��4wn�Q"]���J�7U��M_�X���Q��7A*�9 )A#���+R�jq�<�
����^٩'���`*N�{
�$��V�{U8�{�_+�Zc0��)�r��(����rkЬ���ʰ|7�M�:H�Q�g|���O�}��"��4Mle�`|�M��)hsc+4��0r.�����͊��XIh�%��V����m'��ѷ|x�t�6���o�P�<͵�!8�?`�/̞BV{+�
���n.������x����K.i@Ѵj6��Q`j�!�0va����I�npXrNϴO$<��_�L�~�&q1`�F����e�VIŋ��-S$-W\�D�~[I���l����ʪ6���_!�9�X��:�>�nb|>�K�K�(ƁN�{j 8$4����>d�2��zt
.2/�L�>H1�\1�Aks�k���
�����A1�I�6��!�}�q-�KL&�������Ŗ6�����^���m^y�#I;������0�H1�t��� �.*���p������n!�r0^��Z��b�p�;|Tb�xW{�������h�"�ð�\C+�P��3��l��-X��.0to���q����͍��VH�&.��Y�a��y��QܷsZ��U���i��bt�}^}�P���]��n)�UIE����!��^9y��U����:�H��J3�^Jف�}5�^�.�#�N"I	�1Q�W+c��f;��G���q�=)�)(�jϻ=LC��S�5����a��\��Qr_�Y�����NTV��Q�4h����w��������i���$�W'G8��}U�ӄ��4�/�K����.�y;zd�KS�Aʙ
�D�F"�����S���W����AN����ۛ{�!��������E]��v�]/Rw���C�*�JL����Ⳅ �>�a�O^M��𱰗y��w<B����N�=:���Mw`eQ�+��uzͦ���t�J]a��a�+L��,�-Vt�q����)�zN���2�li:�T<j�D���'Z+��v��X�.E`��"�A��J��|����:�Y�5R����%9	n��g�����%Q_�gE�VK�g\��<�8���\+j%!��=?�q"����;�Q�2R)�ɥڹ�cA;7w3&\B	�NE*�6[�J<� ��:V�X<G���^Yt�!���"�x�,譞[J]�j)N��+-�5��jt�.��h\nt�c9����z�#e���SPm"s�2B�6aJ~
R�<A�֢d�y'�8_v)p�ie�AJ#|b0��n~i���R7k 
L;b���;*���%Q�Q9�XO��p��&CS�5�B���p�k��$�%��W3�9�1��~�������i6�d�� W�r��;@�hbwn���x��q���MtX���u��6�'v=uQx}+�B�e��&�=˴�)�&���Č��L{*��|J%$�m������R�+���7'i�`����l3��X�\̝J�����`X�1� �"�*gޖ4L�V�_%nyÞ�:�&��зodx�pv�N��W.��/}�;_�&�	X��8\@`5�Zְ¾�1v�	�P���u�b�D�����I���3�]���/:!( �H�I��uQZs%�,�4�uz�xL?>!�H��~$K�����/k��I��蠰�W��z�s��K@URD�H�X����W��s9���C�.C� �Nn܄�t�ߵ�0��~�w��_�zv�.^��
;��y4�T���9Hs���{,�B��{^�_�ϯ�rz��C�t@�g�#D}=��*����
O��b6��5i:<WM��"�X�a�Vɩ�ƴV���� �͇�t�oA,<�s�oo*���<m!;��+r�$�hUc����A�?z�2t(�E���*�h(}�.�WE�{���������2�^�M���qE������B
���νT!��h�X	<u����7$�˪4[׬0�ty_�
������*,m�w��d�Q�[_~`�&�QUL]�p;���/@��. 0���k$+�}=���ǘ~��ٽ�[؝����q��BR�e�q,�=���^h��5�O�e�V�^߷�ޙ�	��H��b�����nݏd|�{P��S�!'��t�3Rf�5�n_&4�	(+�����^P��؂w�w1�<ə��̶"蜲���Pu��ЇU;i�c��w�I�&c͠�j��/���+C���Z��gqמ@D�F���T��[P��F�w���h�������P;q�칙p1�����r��_#�6���$�_�2�Cj����s@��l��~f�!�oB}�^IњĎ�+��d�R��52R��B��J`�]��V[0Uu��=c����C$��#��
.���6Ckr�v2�X�s�H^>Խ�4����e�q
����&��sq'f�������;-�%;�"×�
�ĩ���kqV�����9K]����M��D�y�~��\�`���K���)��DG�/�2%��y5�HpN7y	�uH8K��:o��B�5���<�A�@Z}�����p��&O����F-u����
�WP�=���Oy*����ۼ�Z��������j�'��μ��XF�p'��P�d"yDL��?�<[��^�ך��V�(���V���>y��@̰Aj9_3=X^�lW�ɺ;b>�<cUPt��&Yuk΋�fd�q*��ذ~����3x��H���"��k���?8=�x�RU�?���d;������>ay}�~��Iҁ@�
�&�F
׷Ðoa�?�M����8`�S��^ga��r_5��-'ٺ��kݫ����}$�p�
�2�K��l��B��2R(ygܦA`�vZN�;��\�1eN��U#2�9�~��
���ĶT�Z����:�_�5�Eܭ	K�D�X�
@�ϖ���x��#�0��5ϐ,��1mB@̿��ڜ���o�(�a�D[��̿�e�z=�P)�r����,��+�������x�A�c�� `�������-+�	tk <]�GF��*Am�<F?�'����'���6g �cO&�Rc���:&������>�9�iU��=��T�x�d��&?�:;I��"��P�/k���4H�����c^�k�jM��z+�9�v��D��z�=Kd���P4�;�t��������l(I�J'�L��/�>�4,7�*�U���LT��+�9&��|�P4�X���%Dϐt�v��U�C����w�,%�n�P[Y��������-�6Ǖ��U��o[x��2U;H��j�W`.U�@e7��"R�����dFW2v�F�,%Ҝ�i�@�_�ҏ��Z�f�~eS'%Lר�u>���M2��ۼ��>:�᧷v�M�c�@v�*��b0򥲮�s@ӆ�G�
��Z5:�I��{6c��)��xk��@���~��k�IB�|I�a~|�)L����;v���M{y��E�Ý30۠l 0)�*ւ'��x93a�˟:7F�@�j�� �+�@{�K3�s��#2�kb8��P�C9� ��/�"�����v ��^��k�[�
�� � ��5�)e�����?Nr�9��Bм�~:H�5dܕ}�i�
ł�WC�^�#�	�����Z�y"	l�$��ߋY.H���
��X��=�����F�p�I���R�h�؇0�oY5V������d����	Aq��\��p��V��&ֶ�X�u~׉��E�/��%X#J��~쿦�e��0RcE���U��'���mN+�șZ>��Nk�5]S}DA��Ɉ�%Xߛ�8�>���K��I��}����o�O�|{�ȯv���ˆ�L�/ ���Ҿ;���Υ�s����邂�}�j�c�2eNZ�U�����m*XL���p�B_�B�*��e�<��[�0�~�*���7 W�uA(����ꑮ����1ǣvɲ�Xr�@�XG���o�¹�^���SZ�9Ċe'Տ�o�����(�)�`��jo���5M;��[(P��>NVp���R?>A�Er�߽�N�R�`ld���0��w�s�Я���)v$�� ��YZ `ڋ.첨P�}+�d���\y4οr��ƀ���ԩk�L7��o�����˩A^=�@?�Nɝ��Tg~�u�K��\�&�O�M�,BK�(� F$%@��=�N�GȞU3���ggX�2��uAuQfAc.oY���@�!��'D����]�Zb�^0�0��# 0�ڱ��c�����b���6�e�� �;
v��	�~�G���@����?��Iԍz�w��ْ7�K���@�x�s��"��y�}s�����ע$}�>��.�m��B.K~�uXұ���e�����ʇ���d����H���)�40�;�����y ���}��Q�R*���&0ai�Q�w�Sv�4�;��kt 5q!�`��]`�%�I�[y�N7�ab����l�X��7�=I�wh�
�#�-�Dj��V��_��p����-s�iGd�a�XMP����S�f5ݍ�Fq����^d���/�����*���_��1����-!��΀$�% �[t��+@�#�-��Rg��YOlt"����cd�^�$z��j�/N(��v�؛�d��\2VǇSIٻ׷o�u)��7HL��/�2�T��Oj�!f��~PT��ƙ��S�8�������kMp3~�u�H��<�=��u�8P{�����/C����2��_�e\����u�hߘ�˨��i�Ezs��&�5���"��x�`n�5�o��`�±W�͖K=���d!�A�ip�X:���k-A�v�{��O�n?y��@x����Yѽ>;3�JtL3�M�8�k��@����E�n!8x\o��L85��ʏ}�d�SR��ݖ�D�&�X��R:<%d&��&�܁�Ʊ*�~���@K:[���}"n*���#I��^��<t�5��궡ܯd��ΐ����-n1�@��6��<S��Zt��`�V����y�~H7�-�eMK���/,����za���L������+G�
Uw�S�G��m���p�����;���uJ0	���f������pi2ub4 �Ah���}:����"FΣ��������l�E4�]���`?�+l������x7���aOb�1��-9�Lͫ*ܔk}@OT'܍�G�g�g�<W ȹy�����&YN���͉CD��ǐ~����h�����+1Җ��� ��C�o�z�C�r��j�Y�Њ�|6��wjؑ�.�9p�A2���U9��)�B�fTֿs��-�߂pP�.
�AM<�pB>KU�[Q�i9��3�ı=�(�%�]��J-�d�I@v336�?'�;_�<���