��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ�����9���������'x��~B�i��]��E0���)����׭K�IԠ�;B�
�g���;�bò����ӟ��%AM��=�����u��4w�JD,�r2e� a�ݖ@Vv��I�k�>�� ޿�M���,6i�t����]����Y�=��@�5��ęI2Ϻ�>p5��p0N���������
o����z<ڊ�0_6�Q@'�e������
���� ��4 �p�8��9�S�l����<Ǹ�U����d���e�q��ŷ)�#K#Ww$�n)�u��gǓ�����>�Kޑ���Q�� �C�l-hI���B���IK�"�p�*�䣙f�j�Uz�e
E�I�F�_���U������һ>R��E���6�Z	�b�SWSP���mV����vm�r��s?�i_)��]ĳ�"BK',wF�j��!`���^�:6#�Q�(�m�/��ZfO_�ك����AҚ{Vy�X'#un䒛_y�͆;�_���EH��QZ���By�	�z�gt��T
}%�=��?��҄�`<�ҥ`v�n��l`Z�L���F0�h��¤��!CJ?�YrQjE��͆�iW���-��*j?&eX*���q�Us'V ���}��f��Sb�Wf��g�Ā� �!Ʃ�E��ʵXJ�S[�(��q�#�M����I`����ua�t�g``�� N��t�E>���aٿLX�.�+�ݚ.����z���i]XRw����5�.�͂��{4_AN�jv�m{��^ϝyܛ�]��P��'8V��AM)��|�>rk	g�Z^���c\5���Z�?�9�ȬU����4	��;������8kfm�q(�֚/J�5�~��_@S�Pc2T%�b�6�_XY����@�aFX�fh�F����2y������2�@�|�r�~ ���!1��N��[� ���U_�@��ʝ��k�y�:���8=�N��j��{��4*pӂ��h�(�t6� #�r������i�A�hO�\:0�o2�f1;"�jў�L.����ϙ��\�5jLi��������.�%����@i�
��%NT�+1�1ٛgh�	5"�,�AaI;Ja-����˴b2~X�R��d/��$�Ĉ_�	h��K]�m�?A�{���;�f��^��b�Z���h��7�+]y����@�]F<-[�%>�����R�c����F���#Ų1L���O�����[�6In��L��03�{�tB��w�ɐ��\H�N�p))6L'��WG�_2٘n.�y�#H�}�N*W�ӳ _q-��w'&-b(��5������#�n��C���Eҿ����{���.�]����� �K*����
W[bDKk�0Ϯ,��g���C&Λ�T�8h��.ޑ��UN����:ץ���wo��Y�@��J+��-����4CJ�>��1��x/�35��圩7t�ӏ	��5S1zX?�@��]%�L& /{em�����œ�$��ih���Q�S�j3.ы?�5~�Ļ����v�D}0H��( J��)�g���x�rɊ�X����$;z����Lq�	8��X4!��
d;'j�b��c�y�vy-����W㗤��)VvYvv6��j��oD��)��#g��U���Y�$��nĞ{]��^�fI]}zj���~"����~�3�8���L6�1x��5����{���$�X6@�!�%`GV���+��76�f�:��}LCh;�����L���a�@��>�n��8����O8h0Vĝz��f5�\N2�;0��\-��(�*�WΑP22��c�$@��}�C$��w����i�ޒ2uh��Qa��$\��=������~���7�ӗ���Ч/W	���f[��C�3:�����d�hQ�WS�_N��/���ewd�!k��(��h���r�#�_����1 ��/;��͸�Ŵ��}�b\y{L3J��(N�>����P�����	���(��-�X�F�MuzN.J��$��'���<��H����<�48w�<��$d��w�S$3l+�k��ʏ��
�p���X���,�(}<�w��!���4\]ƒ8vz*��DB�=2�V��zt�}"!�[Z�d�|�"���(���pλ!c��Tt��['����uo.�f4�Κ�Ҏ�,�3>yw3�}&�NW#�mv��b��l���! !�lq��c���	g�~]4"���#�p?<F��l,wٶ�r��t�t��a��2(�M�/	�}��ٴ�19`��E|Q�{�6;��l�)S G�Əj������]8�x�`�[���Փy�i�pN�n�-0jx����I=y�D����"�i�n6�IE�洝��X�O��d"<g��\����Gx�&����oT1��t�M�ٟ�ߓ}�/r��I�Y��Ƿ�@XjUA:�Ǜ��w"�k%��g����*c��Hd�&�#����lN%�����iH�XAW�=Km5��"���3L�X��j���H�{����rb��B���_:�t�:��{ֆs���#�_�_O�C_�M6�ԁv�~*� o_����P�ш!���ǭǫx�K$
�~ȑ=B1�|��"��.���
#��2]�O�o=���͜[�OE���� �K�G�7�]��\x���^J��>��R��Cs�*-�j�:xk�b�/�$�2{q�ԛ����y���
��5'khz/�=-�i5?�wecXmJe&��pI`ߺfA�x��mo#e�zTf�+��]��?�Qo��Y��;o���\)�8Ҩ��cŽ��m�~�m��R��E�����.���<�7"\��Q�����bO���!/��I��^��"q�_�1�N����g&sdiTJ�oi���2�1W�v���:�y>�7�i-T	V(~=��=|�k�3�? /O#��^�Wӫ�`i��|�b�u���i�G�7e����Z�s�xN"�C�z�4%�2oX�.�^CO4����
7 �S�p����Ӂ���)�T��4�^iC�:m�[�}�e\|���޾<Щ�;��9c�tg�����y�]C<5K�-���̏P�BH�I�-�h~X[[��Sᴋ�ؗ��lؿ�.��e�OY��(�B�ha'�3�F&5�;47�`���_òL�'�n�M$z:��8�[�t-��h^�f�Cs~�B�3�yo5��0���?�:��G���9�z�5��vϴ�u��8AIŦ2�L9*�SZ%v���_�AE9L"!��(�眔y�/�QPf�wB?,%����D#��2��!�V(�]$.m�Ӟ�k�/�
~� �C�!*Y�EO~v�f�zb��ʹ(fmj�'�*WHÀ��-1v\sS:�]K����Q�-p��~��B>1	�"3�or}ZC df�y	����*�f^�����o睭����x;R@�
=�y{�)�V����^U�O>س^�g&�ܾ>$sK�Ir�U��w˄��#�x���3v�N�A�@<d5�B$kke��w����/�h�,'@����0��R�G��]�v ��hF��)JI�v�ߧ�R�c��d2����vJ���]桌�a���4�\�ۈ�I/b����'����k��;�o��:&�0��4�6�H�8����xG������ ;g&�u�4�t"�u�-�x�RJ%U�}���o�4E��k<j|��"9d������D�l�<t��i3��v$Y�t��p��4��y��ؕ��	q�w	�h�[��_�2�M؅_���玍�#��a�}��"�fڏ(d��r�ߢU/�n���9��z�H�r��T�M9�ũ��ʆ��c2�D��3��	���?7���yM��k��v�&g�0W����֬�p���i�bΪX�@	 ң�I��Ԛy6���Rkބ��PS�`0u݇e.cs$��!�*��53�P�on˖�W(e���^�wV��7�Z��Y~;�̪��N��~�11����-�tl#|8ۮ���\S!�k����[>aK
�JC3v���ٝ��%���h�D����u�2)}6�u��j��ac��^�������ۼ�l����	t��ɝ&7���� ��֏>�/�BA꾻q�,�D}e~�:Z��p�9�QK0��ǜN*�д�|b��,�t�Ƀ��Z�����c�|�9��" �r��̯���׊�	��/��h��ȊU����Ҋ��0�	Ӷ��>TZ8�g� �u��AYh���}�qØ������_�g�o�d�8"c qI �q������L��T��i��Б�"���S��9�_AWkƇ����PfrA�>��|���ְH�[��ۈ~���V>&���H�K9�&\��b�>-����+g���r�>ΐ�%�i�|�6��^ZO�@ѯI7�!��/�Z�`6�K�Ps�B��}�����ZA�q���9�L��\��l����QYj�	�(.wn���Ra�e2)�:�4\��v�� �N�P#���_	\���N�R����,�)�$P'�ÕOmd�p�	�g\)��5Q}4����F%'��*���\���1�9o.�@0�8�����}���\��a�"�0}�W
����P?����>����u�T5��Q�c(�j�g�\�,��Ige;/�)��}tZ�<��ay�E���8E	�d�Jͧy� HI=?V/��B}7D��U�p������������f��l�5+!"'�|
�J��0Ai¥�~�k��#�N���]r�.�fo�b�0���g7����vA�V�叝݃S� �3^��� 4;�b&LP'9>e?�j;S4u	��j��	�����+����,p�24?Y#��qё2�aMô�f���8�6bE\�ٹ��2*�����*��4M@]�s
��;�������[Xu�&��H���n�2�	(�l���1�E�:B>(IRs*����ȗÇ^`ZpT�k��g�C`/FoҾ��	t0v�%f�4�A�=�%�=�U�g��,�o����R+ȉ�K���u�2�E��y��r�ϧ���6t
N��d�-��t��58�/�,����
&���<zl�t���?�i�F��Z�˷E�ȶTwSL�L�� �!Vc�V�c"!�ʦ��M���'�����m�um�Cj7��#:�BXU�>[��q�%���d��{��3j�]���x���A��
�7��te}��a��DW�.�{�Q��j�f,��d���HE�$F'��d�O*��hrj��7k�?agu$��jӯ�K#髛���}�y;gdd(�ˁ��ކn��(�,�ZM*p��0l#w�;nl��.i�MoiODi��X�)B������2�	����l}J}
�TE/k萆ˠ>L������;��b&�# ŉ����ߜۙXB��tW>�ؚ�������V	���~B��ˠ������l o8��fA��T�,"*�
Y�ۡ9�	��Y'��Cx4�5��;�T	#��4�i*d�6���w��Z���~�[a��c#}O�<B���*�;%����,�Lٺ���𧊇�R!����.¾��y�pO�����E���|�?~{��k�`�ln��p�;���
��ڋ�X�ݯ"{��30�%�L�y�@+l����t���+voʊC�/�x�-R�n�ѽ/@�:e��.!m?٣؟[	K&T�h���H����ũN/�:R�Q�9��e���\��e�?m ��X<�Mb�A�ő����3d�4c���T#~T��" �>���By�z��O�n�����)���2����$���t空��j]�qY՝�5E�~���(�I8��Q����և���9zV��D�'�����Y�W��[mPGi�O��x����f�*�YC��zH�ܜP���v�R���ݶ�@�)��9|�ʯ?U���q�Q~�������S|2��8��qg٤��Yʡ��f����ck�X�
�Sv�Y�;5��^����6��0ɢ!e�n��1��I\�_�E;�vLP9�-�x���o�Em� �tq���9�b<�e�%���-���w��pTx�xW��<(:�g�ה����R2�i
�0���6�,5S\��f�	�T����Aht��Kk�+C�
���9��:/��5-/�W����i��ք˝�P�P�gQQ�r���g��:r��:ɌࡰNU�ft~���?z�o�qp]�&1w�a|�N�c�ؾd��4K`�����L�@&�`W�?�Gb�����(����&�y�D,�&0gT��V�Z��C�3[Hr{�^�����f�����~�∩m��6�r���1@�컖{�-X��@�e�Q�3y�[�U!3�P����?cv�KM���ǁ%��C�2���������F�c�$0�K��*o��Ps���uiN�����~ީ�ݝ���	�ʚ%Bh�w�b��t��B��j�HH4��Su.Z��!�|��+*<Eh_N�KwyH@9 ճ2
�)2�E�ˆT�L��f���[M�j�	h�[[@��Q�H��ExR!�`´�݇�|0����/#RK���%����
+5Μ<98p��K(�*H''!�Oyc�F�\�C�s�qZS
�Yl�t����M�=:��D�fx��?Ivgj�ZeF���)nT~T���h��Z�7ױ�H������'�5��De:�V�i���O1�2k��V4�G������[���D6�ɍ���cDI���D��H�r=��2�Ӏ)�E�Sŧu�����o"V�����1�]� !
�6�Y��j��Y�C�F{HG�����O:��ހ:��%'�q�3��[���ĩ~unR�6�Im���9�9�U��1[�� �H��]�c�ic-��{�-J�)�f$,�/����:Q),�f��H]Z���s�������r��[;}�Z����9��(yG�y4����&*HK8~��r4#ںh�l��Z
1��(����8�N�.��y55� �m��반_,w�N����][�g�_V"��`���Ą���aY4ع��U��z�p��8��I�癳��Q��a���wW�����?jg�A�Mф��
�I>��g/� �r1�M
y=)��*���).+�sv�p�lo�/ܽ��U`Qs>�e���F �5���O�+���*�P8n]�n��H��w��!A�M�}��ԋ���)�7��~���P̩=IPL�|��� ��wb������J�[ub-õ-�hT �����Q��*��1�
�=-�b��u""Y��Sρw�t��7�ҎC]�u�
�\�����)����7G��
�D��Ler�D�L�ȯ���2~LP�Ɇ�r��rm�gf�_6��L�ťy�"��2��tw+���E+/R�i��#=�LTzc�Rt�w�!Ģ!9'o��5*=�� �Ӳ�=��Ź�����B�8k^�x�g�����b�'���k�ӯ�tE͛<�����8&�v�t��5h��-��b������`X��'��[{x��,K��ܲ%O�F��#��,��9e��J��p�I�1˩����4uS@(��DAԶ��/�ʨ9�y�ǖ�%z���D\\_E���i.^��^�嫻Ä6F���V��N�
���0��Tpc}V�򨍢X�{���b��~)Rgb�[u����e�u�)`#�56&x��X�	c���S��4qZ�������ek%�q���]eZ�@�:l��
D��Dץ�l2?�iՃ�l�;�Y�ۮ����������U����wje=�}�R_9�� ]�-%}�;��ʊr�f�{#�ߪ꿃���	��K^�z�IE�U�np�m�R���y�x�jU����h����q��2=�p��١y�SS1x(C�<���)�H�TMO�vì������3ە�	��qYnf�c!;3�57��!%�J�p�8���Zѯe�jW�)�����G\�tU�����FuS���26��[��E�a)W�6���鎪��|q��j|��lk����lE�A�r�|��� ���z���CQ㣯�hj��x+,