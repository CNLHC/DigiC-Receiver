��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���մh*,�+��@���V�� :5_s���󇸑#�_$[��S\o�R;��J�u���E�	�B/?[H�z�n���2ƑRk�4<�R�i"�&xט��p��5'L��}�����w�� w���224Y�cD��QgLE0$"�((�s�E1;�Z�f*3w���QCG���,D��!��0Hdx�_�2'�x��V*LK������ѿN��$�C`& �BW�E�ا���������gyW9��\��8����Qw��Fֻ$
7�i�}G����6C;�sҡu���E���D ��&��+�����r�Z��0bP�9�p��J4'��xˀ��4t����Y�o��.+@�O�a�X�Ka�۫3Z_���J�#-��u���zHt�3R�ُ��~���F���i��]�X��]d��]�1���|�|����)W�K��֗}����ݏ�Y+�ڧR�"5R=�_��!���]0�b��R{W�Z��w\h+n1[���`�<R�@�\��Z�V�c�l]H�|p���3���Q�a��R��#g���-��<����m<��?}�\ƽ~�I��}.٪	S��]��7W���NB��U��v9�L�q�N訢Ws��Wv��fp'�Ϻ]y?hG�5k���4�b��+����[9��\d�Wu�⇯?12Bo/��w3�h��NZ����$F�W���τX֖�)�&�Mͣ=�?c}������Ν]v|��#�Ϝ�hP]��25�z�� ��d(z���@d���ک�0���_��L����C��Ob��ˌ�I��l�H�jɢ�����C�tN��-�ؔ�v{����yo�D�mۚ�%UlK�^����*��� s6�XĘH��a&]�Y�21Ef��y��w�0�cr6�vgMߣj�1�	�O7�i���0���m�pZQr�	̀�����K�����ӰQ�'�1��+:g��d�jh� ���m�Q!���[l��=�����)H��=���au����u��Ĝ^�\fվ�� ��e���t�b�me9<����6Q�x=H��y�1����v���Dη(�@p.x����Oiqo]�{ǰ��A��ꦒ�<"���
5�r؁�h!7��f�乸�;<D'��uƻ�"��q)ā�΅�N�o�ShlS�̽�B�D��|�qv�z]f�s/����r�8���Q2�'���v�E��q�4[͟N� ʚO%
�y���WwzJ��%d�K�\��ҳ�� �����y�����L5���@bd`߿`*�CP�ccE���6��Ce��/���P2�|�(G�-��g��w�D� 	.�h�R�v�i��*7���������ӳJ��6a��EY���>�_^*fs��¤��"mk���hu]�{O��Â��&.௳�ES�����2��4��An �Z��@@KC�W���� "˺{tu�-¹�N�1ە�~�h�Ø��s7 �j$��v�7w�	�|&3�}~�KV�J�jÒ9{'�3����Ft�؄
�ts}s	N$��B�i53k����	t8���7���3`�=��U�NM�7t!xh ^ �ļ�g택�1s���X�pH�P�'��6���w��P@g��H�7x��'&� ��^o
"1��̪pA�ܹ�X�xyp=�_�]�wXYCe��k��-�1�2� m4rfa3p@D�\Z��}mM���^�)Pn�i|��	��5��p�X�ݶ��A����=Js�؎��{���������π�ts�oD\M���ʃ����g�{1�IӅk�I�����=����n����IY�[�|Qӥə�({n��9���/�c��~i'��j�ݬƾ'�k(�M�t��tM"���Ԧ�u?j	�6�	Z�q��v~��ѫ ���S�{�K�*M�(�эڲ����Qm����G�v&t!����KD�<n$U�U��	������J�Ť�36� �{)�M�	ߝ���Q��1|~����2���O����s!O�@�7���8����O�&W�[U���L��.���^By�2*4q~�c�BI4/�"9�t���QD�*��vlڤ���6Ŋ~h7�C>����R(��W�ȫ��X���g��E.{�Z�9*������E��Xtm&ݐDHy&��_�n+����	ѓ�B���M�d��	�����W�g�����m�@ȏPn����d*3&
���4� F4��D�8G-E`usC똝H%�1��&�us�i댑�YP=��v�[=*��-�p6�[���	����z���ѿ��� V���[�4^��>f&�v	�D�X�VoN��i�@ ����}Zb.�]�r��[L2d����Z.>�h���^f��V	G�x{?��{{�H��6�:��P�J�fZ h�H4�l�"q��]�B{'LK��-(�}���r`8|�ti\Ȃ������X}x�����[i,00�;����Sj0��\�=�{-=�R��i�8��Lj02
?�������O���-@?D��0�[�i����h�-N�ןO���a6'}�?U�C�w��p�.���Z�`��uj�[t�]*�/&��f��T��s�j0�u9�N8X 靱d_ ����z�����ba�}	��Kv��K���Yz:��z�֖�Z�c�h��G0�&������$��j��n{�{���l`�Io�î�zE3�ˈ�Aox���KE�f�mX+��*�3�caRɽC�Ȱ�H�ظ�ˌ�Q�5IЫ�D�� �<����8TwXx[鹷�<���7V�O�E3	���{���k�~�?:�\�SO��x7.+Oڒ�r�Y�=��h��)at֐j�L[ӽ;D�*��H�gL���
6�Q�w`7͈��p�0�뜮k3�O��m=8����Q��o���1� ��V�d��#�0e*��ak�k���d�M��Nx>����x�6�����0H�~ޟ.Z�tJ����]���M�s
I �i3�QӕoI�7�U��C�����Š�$�υ�:^j4�$�3HDg���	��=��ѕ�?���C��G�X��ԌR>�=���n�Eh^�Z7Q�� ���������(��~­V ;KPa����@����P��M2�������Պ�G ���:p*�d���@Jm:���О5���ժ��F�*��+�L=W��c�Vu�ka��s�F��Dڡw�~ �=D��DDr�'�x�����,8B�6mқ�H(�S��޸å�����h6Y6�@[�L���ZlR�]�Z�Eܦ��s$aM�DT%}�=[Ѩm�㕫�U����M�;���XV�Va��jR��5ԺV{�����K14��{];i��S ) ��5����r|/@cn���O���&���OS(�ݐ#E��x��͔:�[)h��&f� ��@�� r��o����[��^D<-��lk���6`���2+�Ӿ')�n�t݋`u�CS����GT��_��Ǩ�A'޲�,��\�_m���=j���=ڙ�(:� ,<���`ۣAB�o~*{��أ��~'k�)	�B���I�&(����{�1�i�u2����2,C]��<zK�5���O@��W�X��jE��Zz�.�-�������/UU���d+�o��OzjR��0�t����X(F�Ƅ\�+�2��\l��i�/�5V�T���\Y�PC�h����sgto�z������c�(��VN�����h��I�&��O[�=hy�nZlQw�'y �Q(���
��îЏh(0�qT��_w)��Q�q,��h]m�NE�,�:\�ȟ��r��ܡ��i��4H)�<[���G�5�dk�+��\�K�k��瞇Y�]{Vy��*u#?��MmG��|�&�@�S+j@%ט��\�G���2�j�N��pU*P�/(�hR�r�&��U���8A^����p����ڈ.Y�]�PB�i9��������ߺ�M1�B �0�o�v\�l���*��(�� �3�����:0�k�N ��\F#m�e �
�i`m �>���ͭ��<��}F�GN��Z4i�Ո�ٛN�|0�$�I˲oKFZ��,�%Q�6!1�����:�O�ӀU�C�w-�Tw���3x���(��'A�YW�A�y��F`ɡv�Lj��@�m}�3�,Z�����i��7VD���uVD