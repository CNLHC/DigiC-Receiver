��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���_c='�ؙ9��G���0e��>�cGQTi]h
tL��m:�������d��+˵��$E��UV�������a`ԇ�4�����!8��ұ�����3Ѯ�����-(�ˤ�P��_����B��f��T��r���!�Ux",�q�����{��$���)w)��oc>��X��mcb{N�9�y�D�X=��TPGpc=��S	L�7�a����v�y��kj;ceԴ�G%�y(P�?�#Q���c����86��'A�bUcˈ0^B�eH�2ѳ��q�����{�7�ֆ�-b�~Fb���EM�ǔ*�s�#�����y4{)�/��o�9����_�Z7����@_�e�o469��ĥT�GDZ�-FF��I.I��xF��NWt�#����B�kq�P��4QN�\�v*D�+�Ʌ�2Tq������J�c��u�nmz�(����\��yB�Gd�����)�N�����!���H�BG�FaF��Lg�o���#���H�W���CSG#�&�q4��~G��Pi@�^�G8xw�TI���5剷~�����-��J�2-K�v{�e�`�
����9oS�ײ�N�]+:�`~y�q �?7�[:J�N�=s ��u�X%�2q;P1�(�D/;K\ܻrr�ț�6̠^ft3��<S�L|�]q�@ԣ#��T�`OJ�lM0�Á��Qd%�����踃��ho����dR�Q�,*E�i7��e���F1>�EܹCTnVﾳ��51o��"�7�>������ku��+���������U���ٚ���v�<�D�� ��2�YXY�:�D=_�Km!�����XL]Z����^Eppk�8h/���2��ⵖ1(�N��:�|e�1-�j�YTƖp�.U���4�llnEJ�_>٨����w�6Q|�Jȡ�*$=��>�Y�����ģ�1�5��ӿ j�V�}��d,�5;+���\Z�_�a1���@��(d��&�_|B���*v�9b�����G�K�0�8��V��|�X�=���uɶ�"9�(�hJ`����/��h�e4�=~����@�6/�d�q�2?�D��z�064tC���!s���lvf�箴m��3�[�5n%6 �:,P��cm��$���4㨫�c��u��b�z�>��4<&�= @��ʽH-�3+_�ֶ,�^� �?�zV%�e>�㱺2�6 NKc�PU�EI��a�!w:i���JK�c��B9�Q�^�{~x1 ��nP������c�R�^O,��3�Cy�'>Y_�oz����V��
N��8�p�׮�Ы��%+ ���8��TݦO�f�r�FB������` �`:qE��v�|�/�CYM#�������W�^������Z~�nT3"	���_�X�
B�^'��������S�4p�1���;�o��-�Bo��R��� _��j2�c��0�'�5Z��z����75���f�U���|'��}W�3/����K� q���KE���bK �F��n�[Tx�e��2����r�%��X�eK�,��q����r�$E���
]��K����ae�g������s@���Þրᨏ�t ]H.0��V�-��}m���l
�齈��j��HS�,6N�����ܸZ^s��>�Bջ8�3�rA�DH�Π�k]������_xh5kh�� �K̏
0����
BTl���]Z��w�n��*R��I�]+wW<<�QD?��Ռ�ݐ'^k�fu�bn�._�ʔCg){��a��6P�*�y��:��"Ãu��n�������$9qO2'@2M<��4�5����8�edch�4��N�A"P 6��C�/b�r'd��R����`s�]C����'��9��J�2�HC����ͱA�W��!ϛT8�mI�/�g��v�[/��&ۿq������$/�+�Pb���i�M�*���\��P|�-Y=�W���w0O�֕��U��d�^�G�D-�2���>H��W�{�8�H��v��)�0p��� 
��V���ƒ�wH���Cj>�
��������y�~���K+�<�9'�tXٯ����tn��P�� �+�>=ǁW�C˼;�\�փ��,�6���l�)g�uf��@P~��<_�s@\X��hn/�x�*��Ԙ���K�8ܹY@P(5/�Ll��2���%�Ƕ+�o�/:ʍ��>��'^	��y��R2�k#ӊ�REg����Ɍ���~����Eא$M��Ź��͊��֥�!(r'��8{=l���`j(�qN$>2�
�m+/7%��n���-���Q p���c��*��p�lR��>���_����_�D�D���;��.re�۟�k�Y=bI�z����HE���]P��f��E�I�=���2�����k����v�w~�;AWqآkv����v���"QX�j�Ϥ���b�����%���q4X����CW�P������wd";��>\�%k�<dH�-�y�;�R��X����	�P\EY7F��\Ĕh��Є{�:��WtoV&����(#� k8Cip��E%����G�O��D1�2�w�l�0�-�P^�&ߥ�n�@ q�q;���Y�񒓀!)��Wh�}ݹ�$�?�|D�%<��f��q?�����;�u�0]���1����6\�诣�tA�%.�X �KD�ˍ����'����,���z+����-�e3�4\���Na1�(���'��֖�ϵ�-�sCp}E�(�܏�4�{w��'(٨�ƻ���z:eX�l� ag�GT�On���f�jSMqO�mo��]�;�L�8L��c-��
_l!$3��ybF�.��U�tў0�8+N�� 0G	Q�?��:��� �D������X'��ܔ;GP����u1�]��������Z��;t�a:�*��V1�a��A�p��{�n'���
�KmO�.O��ԡ�![K���.���9��q�]5�}#��O5z���Q�"��,��bfm����xC�'<7v#�����	4u��}N7W^N�#h��	����П�,E���x�B=߱��2�H�_����)�����\� P8���ρkK<�ڂ�1��Pe�!�W�<����\0� E�>�[��=�z��G���u�8��D�*��vl"_����O����Y��x����_Qtl����l`�l�q"���%AF6�pO�*�`H�"֢��xI��u�oz�{�my9����v��2~$���I�PO�Bh.d���߀J�M;� #S[M�1�9�}�~��C}B6�<ݣ�����뜚t�E�mm�+�Vmh���E+��1�|��VK!�X�8x-�̓>.B@�\��
Fi򉜺KW�عl��a���m���7�A�v�����R�jƊ�㚔��nR��ȱ@�NTq��'u=j��y���*���=i����_k9w&āG�sc�G���!�Xx{��	=��+QA~����i�a���,��A�F'̧'��V��P�f`{���b��|b2�@����u�'uӍ1���@����U:^�<!Պ�n���	���UN-�'�X�3o?F[[T����H�T��7�(çx��Ӥ�lq�~I������ il�P�9P�%������ǐ鱠�%���ݴo�Tj���7��d�ў�Iǽ���N�/�-�#֤��e��5@]b�H+�*��a`!e3�@#1�0�:���[.���X��s��+~���Ƅ�7����s�Y�9`D:�$�~��S�N�V��'�]J�jGɁrD�|��hN@@ȘT$�1�
}�Y��V��4y�����ex�Cf��Dq��-�b�Zʚ�z���ܹ`�U
V���p���2�n��8���`�P�e���+h�/�r��\�K�ns����Ȃ��l��A�p�J�J��<1AY+x����"�l@ b�kSZ����}M�e)� =��HD���t�q����k�a"���A���yC�� I\"��mJ�׊-�g��|AY�I�}���F��-0�CB�4-������ߣ�U=�2��1x�l/O�L
8cU�o|��F_�����fu�,?��PG�����h������p~���An���+֋FX�%خ��>�Ç}�۶�G��򞳯oet7?]���3@�>V�^fz�؆��=.�,J�����/n)l.��f�:�*��x�{�L9����}��i��/t����_�@e�rɽ�
�G[��wc��E�V0:�-�"�i�+�Q���k��t�@����Ͽ����C����I`jX���8��: SY#-�l8X��rW<LIL�m�'���v��\%�Y�NW��j���*B�	4�9��֝����\���W��)��|kt<�Os&�����7�-5�5���N�e��f����u�MF'����ۆ�f�7B��q�����j��U�"]��Ar��n�$z��9�����y������m~ �[�:M3~#ŧ�j��5#��Q 0��2�J1��*M�JЁ2a�Y��A1#z��y�ص[b�0��F�x�T�Hԫ<�yjR��%!V���`�i�c�;`)�s����=,�2B��^��<8d9���}RXu�������ٲ� ?,��^��/(��5A��ܮE���pnYݕ_�	O?QOW$���J7�h��M)�n�y��%�\�3u��/M�R �@"��w����J:6E�������]b5x�)��qc2���5�I+�Me�f�@*�tW�2��}&]��<Q��b�&���5���
��2������n����	��E���:�gVQo� �f[�	=i0�W��'2�N{톹�*����Y�¼�*xZ���.]CҨ��3���~���=��E�V￯�õ,W�,�t�hN���6�;�*d����^z�ӒB����I��a�fk�An�I�x5�z`�*i\|���1��5��P߿��7�����(�?rU�R�5\��/���c%���,el�U�,����s�毹�Ҷ9�
�6w6���xF�n���Х�Ϟ���ٻ�v3U�ɉ,�R�N*��uB#��L�֓�� �?}k�}�8��"��w�R6����h�GlQ��J��̯PEeQ�<�m�#�,��h�`1�-,ӬM����%PSZ�.xwO����\��g��;5Rs6�ؓ
M
�u]5[��ւZ8t��B�� b@�ɓ����]n�7a���iV~@w6�V��?
w]��_Mڹ�33$Y��æA7��x�7сc�j���q�.�(�/���%.�2X_�z%��̷W���	I�Z��}�Z�߯Q�Ue�XazMi���9���'q1!���$|�o�5�w�7�"��<�W�h�{���*���5.kzW�Z �/e�3s�ZY��Ǎ19դ^Nϐ,!H4B�0��Z���u	_����G��s�����!9_JT��[�d��?�l�_o�]�\%T��	Ib����vh��޹֣�|��`w&]��|����̳�+��b��I��Z ���@[�,h�m������.��X�y��ޱFж@��q��Q���r(�&�RM�ˡ��E�X<��^��Z6�I1�(�jw�=N���47�X�`äX:+a"�I�>������W�Q��=[1��k�^�	�۬���I�{����ɟAlv��V��۠�;��I��r���1Q�+
�c��[������\8�/��R�n��יEC,{��0�����R^�mޛ�U�	�E��a"�^��R�>�&�W��I
{�P�MjrT��-�HN,��+W��.�gz3\7�0>W���n|�荨�b�&���e6�"���u�o��3
�<��A�4P��K�"�M�h�ä�ן4�\6��6���s�tLE��N�1q�G*F�㈕�W]E!�G���8ŕ؍��yU�١��}��;����L���3��*p��Mg�(A�~��(��=��[�}&�,�i[40��'&�k���q��YSOVtfԝ�xa�%�z���]s�n2���t��6�~���+����H��c�[h	��iq��Ԃ����@����o��.�8��͚^88�EN#І�]�2��g�\YP8�:�6�i�'w�GB#��#������ �Q�u?᩿'A��\]� C*�p�ҡ��Ύ$��ЈVt���P5n�$-�ml6z�ӹ�]H�W��XTd]�g�t�G�c��b)����^_;�T3����`��@i��LJ��Q�Pf�l�r6�`##���wjl�l��\T ���oz3C9�n���}��&$�lO�'w�fo�..�e!��eG��g��C�kz7N;��LA��>��3'4p"�����_L�uO�5���IK���"v�|�p�d�
�jx\��xڡ��('=��A~m�v��_���#YK���W�}�&\d+"zݛ�q��j��D����f�̋#�+�ٿ�}!�f����8��3��$%�k���_O��5�G���9jg�p�Tv�1W;/�{u�}�6,� ۘ�!.w�'��D���]=�wۖ?ɑM�����^Bum�i?)�ߟyKÒ��Lg��4��ob5Uk ����q���H��&�F��*`�>D9�uD}3�ׁ��Z=W��8ָ��g�����O]i�H�=�3T�O�'%�O�U�M��ak׫�"mޡ�緐?]��.��5>K�+8��pS�Vk�*P��_n���!�t���%Å�3(Q��ģ�����+��B�z��� $M��؊v�2E{
ɽ4�����?��OS�@L�r�w�|�4��a�~����=~��%'gzT�#곓��+ ;�s����!�^�+@u�u,����4j�S�e�!��fv4T}VC8j��eD�;��L���c�n{�|[w\�]]�P�ۗx��8�n�e���nι��~�G���}<��T�L��FƝ�M�'��/ˀ�dɃ�5��ټh��z�1h�fK0���W-F�.i�C�R�G32�?�6��+�D!pݿ3l)����^�5]�M&�lq�!s�x\����A��� �m^��uׅ�k<e���R�ɩ�LE��������yz�a`]G��˨�uR�����7�OZ��M��e��A�aLe�����Q�B�>�$��@�����^a����ٻ�n�؀헌�\���X���H '��L�b���e������~`#�uym�H�k���,�Pj�x��N��m!j)�4�	ׄ� �_P�DE���x��Cӧ=�e*s���L'�g��.�`�P�K	��m�D��T�il���BN_pA H-�f9w��[/��� ,	JUQ����;F�Rv�ك|����n�%��8(�!�;��	��FjvX�sH��[+~�mK�n�Q�2t��°������f�$���d��0@+��L��$2	����XG��8T��bC��=}]ԧ"��XS�����se،_�p�9�����g��R�c�r*�ٵ��]���1|4ڧ�N}�i�o�?uN�¢x��E�i/�j�{:�|NzR(G��`ע�`����t�w��r��X(Ï2w��L�k� O�"y��y�ᗹ�U��X��57�8�$m�F_�4�HA�%�~��\9�1*`�5�HB�8_�
�Ο��	8*o�M,j�<�mdZ�]��)�!H��u� Rz/4��v�I�sN^��c���6��ޱɃ�-f�#��ಕ<<��w�LaB �D���י��n�T$�# ��X��e��q`S6�V/���b�&����W��ɼo�p��p�ѵ�u��JnP����oy�)� S�$f�|-g;ȯq���J��?m-��T���&1J-���ʶ̓�{�%g�X��CaY���_��֓�<|����G��	gETa��V�e@�6M&@7C�nۣ`��)0ñ:rw��b������_
Ii���xO��'|��5�S�p��u��-<-s��?ɯ!L=����Y�������.�f��Ǐ��ti0�8��E[9>l� ~��[}�H4����������n%��F7g_�=��k@�48�̙��'�am������e\�0�U�g�#�D��Q�Q���o�6��I�ʶ��C��?{�[-�D�H�>��2j�C��е�i%8��u[D,�VA�jB�H��¿�m�򏞂��1n+m�"Qv�?,��}���o���?��� ybF��P�Toz�o��s�嘼�6�h�G��S~�-
��N��:��)�&��:�T{U�;۸;� ���x��8��*�&�� ߺ� z�а~��H³3Dۑ�'���eܶ�?(.����(vė��4)�,�c��=���y���퀁1��æ̐?��懺�m� ����B=x��޾ˇ�5���Jubv�#����)1Ȍ�c'wL"��~�KEz�w~EK���Wx�/�Z�&$�W�;1���G�ϜuH�ۤ/6jO�:m;�gR_���x�!`W�Ch��)� �9פ��>c��̏b�S͜�[%�n����@�U�C����)j�X�X��*+�3f������$�����6������R�i��)�1&����9�u���8�I���NI%=y�,�)3w,�g?W��S��ۿ�$#�D��>c�7!4<���ۻ��O�i~ы�> R�]�( ,�QnF��* ���mk���7<�p��Hғh�,ye�,t���c�t��k, �7}�|���d!}f�,�lBx�ĺ��wA4�T�ε�dSnK���Q�;y�w��_�-J�)ʍ��LvGG�8��������#l��e	�����B���ᇽü���̷{z�x�m��f�V���!�N�%���F����&EQy���c!��N���ۋɅ�g\��=D`]K2_�h�$B�$�3�H�����B��h���HeEU�T�n!���8j1^���}��Q��{�����_��;á�[9�L�,Kb��(g�e��\b�pu��R|]���v�YG��u a�f4h�QӤ�T,�r�õ#�A�?�vL���[T�Ew�^����8Ѳ��FR�9�]�~��T\��}w!��#���$�,�k��1��v�v�0���e�$�#�0��.�u�,����K�I�$���u����; L�P͙e���aɵ>C*�`_/�v����E?�*�<�379l^��T��}~��*e4n��p��nǒ��b�+��cю��X�7(���(S�op�N1��l�w� ;�`�1ʓ'@�uK��dI�}?q��p�D��W͡Y�g��D�.�<����
��<r,p�M��[��[f�^+����=�^�����/PD�0`��w��j��χh�T����0@p\�0u����G��^��H�����bk$}&A	�~/�\�B�
��H��-��/���M��Dw�/�U~*&H �q�7��ť������nbS@ɣ?YHP�o@4l����T��v��[G�H
��]l�\�9N�L݆b�@;���O�^}��a�FWC����2���cmP��,��9�E-ėA�#�L$hw0�tɣ1{$i�U|C��ϱ~����{����G`�?W�ss��za���˺WT,��u(�̯&���o͢/�.���.�D�8�
؞hN!s嗈��>҆�<0�>�=�M�����z�'�E�4�	��Vk�t�X^���`m�D9$K�7�Ub�p����`�&����������h�O9��F��M#''sD�`,�%�~U���e�_��kT�Ŀ ��<�{
��u�Ƥ,��D?�p��3�J�7�h�?K^�xsҠԜV���Xn���&c��D�9C:o>�c�Q8���8���0첃��*��Iyo� �u�s@�������&#�1�&W}�HDZ04Ņ\�;0k�PU5H�t������e/8^*Xs!O��(Y���y��"�
��LQ��1��W��t�!ME��:����F�K@G�q�Ї�̟S�DkA�>���X�����)j��̤��*i}2OM⦝�(�+�\�:�:y]���ԡ�M�*B���,������J?*m���^�¥�i>�,,�TV/�e�<��˗BU]��"p+.��.p%�H����|�z�oT:A4�k͉��c��|��r=�u�!e��0�`5�/p�v��G�8d��)>.�
��j��m����L��T&�סW��wR��HXD�����M������:��=tּ@L4���N�xA��j����W��¡�OE��m�Ӝ.7�^u
J��Ԣ`e��-]�G��ᇫo0��d:�e��W$Y��iͽT�_c#�h�5���8�X� ��G���?m�Y��19<��E}��c�d��Һ#����%�P�H��J�4n�M�I����I� C�
�
>vQ���Mыh�H� <�}�}�=ݥ�V؀��'�nh�1�w�S͖ϛ�P����4�^Z�S(�Lm�㡢�>����"� �=��u7o��GV��q���_��9�0n�f�`'��$|ˬ��.��f��,�L�۾��$�w�X��)����6]h���	��F�t�7�'���&���g{{]���
�7T��v}˰t~E��Ic�v�B�O-)��:�b��A������ZH�4ε���������"@������&�D橭.��|���!� W��t]�3zoGn�]t�'�Yuo����h��2�!"pt�H<8�Ef �@i��I��f;�x������m��` �*��R��]FxH��|�����<��o���1�zf�Z�0��\9�g�}��FM	�)D�f#G�U�g�&j�t0�Y�	�s�)�`�^%�T�6?�Xc��=�ٗ����Nnݸ1<��Aqv���]����
�3����n#�n�#ضG��Khw������[5W<�_���U����AO�Z����j��lY��� ���s�