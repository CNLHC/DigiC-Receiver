��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��ǒ��=���pOwA�`.�:<���+<_3�� ����ӂ'����n�S�~9�)�'`�"���4�����[�3�絽n:w�ߟ9�N��-	�Qo��r�෎Ɏ�̤���%���q�#�+(BՋ�C�������ƕ玗1�����(T�c��Bc��3$�%O�������s�1�,����<��g�۳p�G��QDn��۳|�����D�����D����o�>���(�٥�{ݨ�.Ѿ�שC�(k��0@�pP��b=>� )�z�ئ�s�<������k��y�vT{��G��Q-�f���~;�Z=?��}%w�d�|���ϮJ�����C���U����e/郚��E��K����d�����2(���n�)T�pٮQ�X%��-�Y,��)�\\����V0�x��e�?p��9�m(6^�$)�5�R�[�ͺ���� mifY�%�ՔL>>�$�x�z�4N�͚y�K͑Ś��P7�@�,�cXI53$�ˉ���q5b��{g"�G#]M+�>����S��0$i���l7A�<��R"��DV[W �
�}�H�57J��2�}�biݒ&��;���<s��j�H�v��>9�j�KΉ��ʠi���V"l���3_P%d��~Y�{�T��N���&�>��mr���U�Ҋ`6ꮊT�-���6�r��ȿ���cT5'�Y7��4n��Ǧ&V
�6�`��'2��g� ���!اT�U0hv�����5����yCd�
=�}�1�[!]K��H�-��SՕR�#@=0��tVM�K�� |��'f��R���H��=�$]�A	[p���V����2�2�%>�^I�Z�R���듃[:@{���g�����e��?K�ڈ����ҵt�����>B`i�A\,4���Y���Ճ�@��^�t,���@�Srp���=bR.�Pb��)}��A�>f%f �8}{V���{t�ꏽ��U̴T1p�2��PkM�m�>D8:,�!�y8{I�&���ܛ�	d��q:��)�$�\��%[C��1J\�~����
�*�=�3Y*��K�m��oϊ[�2�BN+�ٿ������o����?u��V�x���h	����A~9UyB�54�A����A@�G{�(�[�g�K��Q,z��8�(a9�J��&�V&�a��n�ݻ~^��CS��x���zī$�tS͒Ԩ
sxVO� S�ه(�"�������I`MV�%ʘ����B�kC�+��6��A�]O�
vsz"j�S'��S���#u_�U�X�9�Γ����
�2pe��?���|߄+i.p�Uȸ%��~0���TҴ	�"�W~����h�u�la9g$xK�ftgD���.:CG-��*/�~����!NC"�B^T"]T�}�ԝ"����c;~��_�h[#�1���Ƀ�T8�Pf@���˫�Ly=���;|%����!JB���@u�����~lCٟ	&k�|D;��Ӧt����e��d���G����}~i%Cv�
����	M���ːOV���an��|;�����wu����x.3���ܿ*���f�T���}��7s��Y��賾`���Wwi���GG��q��l�QA�M��Z��d'�%W�]T���w�g#=q�8����+R���Rަ���b:ë���챓�I(ֵV���$3Y�!�W�B��i�o��Gk^�x�+jo5�(��<��ٓDH�SE��!S�B�@��__��~	���P�B�ս���{)v��}ͱNP;I��.��'e'j�䒈ۿDm/�/����(�4��/�2�ђ�O5H�(�[�8���#�F�E�+w&��)�a���S���9��$86�+b�S�>*�$���R�Ғ�#��iT�M�Ai,BǇ5���§*�ѥ|�� �	��d=/T�{G�e�2���N�E�Wd��\���<G� �[�ǎ+�׎�ޡ2���c\�wq�뽳�,��r�s�^!����UP�lQ(L9He?v�o �8FKפ��h+�5i �pi���<b��)W�%���}��*����KJ����3�G����o��7�;�y8�3'h0E���I�N��\�fJE,Λ!rwb�~�\�P���-����X�e+���D/���J�(/FK���V����n٩���63���8�ָ��w��<h�#K��j�nD��ҁ�Yö�j��59�&^�G��
�x�p�Eݟ��L�ۙ�ԳA��.j�(�{��!��ֻK���7"N��wˠ7֡����*�����?����C�$��H"N�_w�$�֯:�{<n��hê���R�g���tb����N{<5m\T�uj�M�
�ml���K���W�'� �W<�/���o��,�ڠj`����E�N 1ۨj�EL�$��7T�=�o���fQB/�N�r���Ɯu?V�zЊ��Q�����<�_w��*��i�NWz��p7jXI�r�a0OL����A#�U>k�S��N�Bfӎ��Ϳ�b�ŭs���`f����)\�_��%�Ǘ��M�6���\��dԀ*ά�*K� -���9��<;���V�������^��;�"�X�.d4����j�`�퓽x0�ֱ��z�kXX%��Q���%[�!������r� �91߉̝;9�H�}X�d�5�H�U�>�s�-��/K1�h�e�`O��e�h�Wy'�e����u,}ƅ�Q�?����	«����}	A$���cZ��ސ��jW�<_l����K�
�/�\c�FQ~�t���X��|S
�ᚙ�
2�ee��PZ�F��
�����-�7����MkҰn�Ī�m��S\���R˼�z�_䑦��q�!a��y1����=�cQ��Wi呠�p�u�=3������UC�����;b�Q��	��Ct�#D&>_!j*��֏h l#ݱ[���U}��F�/����&����F Ib�*.����UD�X��J#��\�P��!� y����A\�Q��5ձ@����ARť�I͔�>�F)�&�H�T���T��"��G
�4��w��~ۑ�f�m��Z�gg��.hU���k�OviR��)u/8����Mz]a�Aq����<��-��Q�:p;�P����p
J>���S`vI�h��/���
�wM+m��ZBV5�aS]�u�,���f���D���ݞ�9��N2��\�k���{�/�{j��9�Jp�`L^�K��^|��g�{
�Y��6��O(���(��d����"�c�c�)mz�=}���nOb7��6� ��z���Rxm���Dv���O�c��#z��P�I?IXk3����mWdc�Ȣ�R�2mZ
�e��s'#�ek�j��+D��Yq֔��F��ӿ�V�'.�{%�%"�n�Z��]b7��ù�yZxu,��[F��
gs!o��Q�u,�]?Cc`�[�~{_	�e����<�[9I�����܅G[W˝c(9�����ƥ6��ۆ��D �X@d,my���0�HE�@>V֌@Bt���2�����k�\��o��J:h���qX>EHgٔ�j���h�)����&�*k�Zm�_��ÙЗ������z�m� /�3�j�&��u���F������`GUH=#W�@6H�� r�l���p	>��zjoc�~�C�a>�j�~k�Rm�+O��^a��'�p��o`�Îpk�]�$h�R� ����^����R�;�s
,ߴ���q9ﮰ�A��q���s4�V�=������9�I��s�ՠ�T��c{	7��G��j�y�d��:��YtE[�F���s@ލSn��-{��j�ax�eu'��C��Z�Y��!��1�mQ����5F�S�	t.������a��K:�f�X��t�@`~v��S��������O�`��&yLI����z���"W���#bi5`TJԢ����4� ��z�u��!10�C�^H4DC�ߛ���2}׻ލI��Z��[e_�C UB3�ϹN�r��[�'���SCI�O��רAK6d��UP���w��ꢢ�{���RK��5a������?�ܧ���W�Zv>����EA#|*^Y	�ۍ�)٨U��<7\�?�Di�m�W�*wJ�F~A��U�M��1*NG�B	p7� �JK�	��Ł4��
T0���\�8��]I�X�i�c�{t"��j��O���o�4E;P2�]��Z�?���*��a�S��cl������'8�"��!����UU!x�G�#"��b�7v��x�t xE��������΢�@�]2�"�嗋�i2�����%��*
~�CKDB����1��y���1��_p^�F���!�	wId��S'�����M��7D?���g΀П2e1�{�����5��&�V� �;�%ĸ�L~Q3��kkxm��b�Jg��ϼ��6��r6ie�L��5B�6QbW�Ԁ���ȓh*Nl4̉ ��g�WV����tg͸��UNIO JgEO��3��m:�wњs?/�����P8�����e�d\<eT��#-�L���	��C��.t_�C�If!�ȭ����8|�Baتg����΂��kcG`
�[5���[��)��I��t���FbÃm�s�D���	]cwSR��gF���=8\��U�� G�Y߉Lqq�Z���7W�?�aO�޷�^3�<2z�i$���Ȼ���Ӈ)���%Q�֊�
�y 
�g"�ˬKF� Vcw�Vd���N�r�}uOv�<�䦌d�;�FU�;^������6S�͗N�/Ȇ�N@�����{�Ϊ&�-�	�<�� VN���,�d�8,(�[7��E�y��a!��n mw�DA3��������D�DE'���j�<;��/���Kb3Ѹ����H��\\�6�7f��)���te��2we�HL�z�s�nh���ʧ�!�k{�F
�
�@�_�Bb �-����ƈ��:�6/O��2C輪�6ޝ�Bwoh�2!#�4��)pm��t�����t��<X�\���=X �O�a�Y���6�'��Yq��?��%�i�L�Q�qh���]�t®3����8��3��Y[�����P@3!(�d�c>+G�q�&;<����f�a� !󨦫���dIQ�&��Շ�76�6�����gճ��&s?фfSdp�ۜ���C�9)`Ȋ$���ГUZU���C`�L��:��%�9H����_��澹<��u"�bZ�Kw�	�l�$h�[OdB�0��9<~�B��'�zm��O��Q�)P����C����W��xb�R\��
��J�J|ǔ�a!+�B��s���/�~f;���d���s�r��xMP���V�я+�'j4O��W�`��Q�;Ɂ��ڔ�h����e߽W�C�Q��ܽ�s\yiA�Y���O�sq���e�����hhsT�W����b}���J籞@�1d�c��*`�W}�~`�I��٬�m��t���!�*����J����y65��ӋK�.@�֯�H[�ԑ�ל#�;��6B��?_kF
�J�o졸<��P��{����݌"ri�Img%�D�W�h
�pS\'�@���TL��]S�:�P�S����1�t �����&$�τy�O&�T)�i=����(ʕ ���VG�JeZ�룋K˧
Y%�P��7wӎ�t(���	�)�V�} 6�cL��(�q��b��o 1!�a-xI��f�s)���Z���zy#Ф���"��°ȋufw���P���]��J�B]�n� &,&�<n�د��>�-�E<�:aã��?c`�-�������'
\������
l��e����[k�A�'" P��>*c5�uoGt���c��ǧmH��Z>���â�[!~������5bȼ�X���.�&�b�/K�3̖ X�w�l�雋�/��(�ԕjt�ADO�cN�+��k>�&�0�Dx<����{^}g\=%�H⺈��κD��q~�R��?�� �M�R�o �VP����-n���ZxI7���˟KPt�y.�g�����=5��@���~7_�T 'N"ψf*r�W
�ߴDeF �ؐ�v �4����VJ�u�:pE]�})�oĉ�`��1����ӷ3(�k����a ^�j\7��-&�C�=x��AI��3���.q�&4��G�U_��m�+���~��Bs��~�<f��}���F�,������j����[�g��#����?���6��Q�_�TW�Z�sl�30�������J��!'�E��k�c+.���&�f<�i@�@����c������[�@�q	���������q2�y���ѿQ(�Mp�������qE�nں�����F�V���V��l�g�O�h�lǡ�H�2�-Dw�0���x/�'�q�~"��Ø�'��?0���"�\���@p0��� �p��X���;����ķ��ʽ�E��:LM�nS��|��IΜ7�B��M��Xk�|\�L�r�z����y�b=N�Rپ�Iy��%���? ��(.Q��Ԧ@�孰�@�g��o��[I=���_�j��z���y�@��^�&���D݌ZW�	b��- H�}2g2S�w�K��8+̖����)+�]�Y��|��0%C���#:�X�\�H@owЏrߍ����1�]�E~�A� XD�ge�;���ly�_�ʹ*�4�s?�^V9Ee�[XR*�9M�ée�@Rw�5�w�y_����~�ff�*�)�zL��6@�_(��o'f\:	׮.�  �u ��Z����^�ρ�b=~Vw�;��߯,�%m�)�K��J��:�� FxH�?ͭ�>Q[��%�PBh���\��E��PݙP%j���Ҷ��PJ��C�s����M{�a��v�ѡH<�U�����Q�MG�7�����w�*mB�+�
ϡ���1�P<[U1��b��:��3d�惿��3
AR���p�
���8�}:��D��P�;r+8uenIk�;yEk=n��c���?:><ǎM��ϲ�W�"�S!���E�����hѺ�m��^
�@�;f��=#�� 8 �	od�k}k�m4��ѕ'�������MIe5�kyqnB��Gﳑ�ů�#�-���n[Е
�'F�ɜ�P�G�����;?�:2�O�I�%�~t�>�@�%��"&͢\,��#d�_[^���B����Z����,@띪&ˍ�c��v���	�(Ng��N�SPX�]Ne��yFs�PS�H�q�ӕ�N�
 ce������<W43��U
�
x3gF<��U��-�-��� 7d�U�0<�߾���l]Sڟ�d3�̝��SG��Q��D�����g���j�Y�z>�ء8,�v0e�w$���y�4H�e�xH�O9ݜ2��O�\u)����O���`�zS�j������t@��T����������W[��,�cQ�W���?��6�a&�sJ�X;��  k�$�%��OE�p"רk�}Mnԣ��� �W]0�����̫���ˑn�7�>&����P��B���1-_�Z��(q頻�a W����k�8�8%�VO	{a;�}kt=�i��0M��]�9��bs��*c(������o��0�-;�E��_#�i-�(��M��Xc�&D���\�3������B����	�Be�!�s���K�����HX:=J=2��8�ѡs�QV�>jY3#4���V�l�a���u�K�\-���Ă�]�R�Ɇ.�|t:O�Pɑ��߫2V�<����}�T��=�")5(��~�ᘾ��T�D�%b(�S>�S�v�L��o8Mv���n��X�bt^f±�5O������W�4IڔF}с��n�d� 7�>k:�a���G:��E��x�'$ᎄ��1�oKˌz��[�����棓r*ՉkN�}�	1��#��&�Pe1�c�����x�=�7�l!�k,�@	��c��Yy[+).�:-#陨XP@��J2;t�u��K����7 O�b�!L���X�U��,���Q��HC���	p�Ǖ)a`�C5Ec���'� &�<���i�k�X�Gr��7N��")u-zg��k�������!#��JCbr�K�o�k�U�=+���n�X̢r��:�Gpp�� �9X�z-�CGa����;z�/4Ӧ�r�Da�I�+y��f�r�m�Ix��!wN6��Q5�i.������t��zb�h<�X����O�4�M隲�IH�Mَ�*�%<�T��0{�<��]���Ђ�̀��r� *���j�yP���DV爫�D��/tőF��M|�����/���kh_))�|�c��Cw?d�|����(�2��~�Y���c��DR�o�
x�y��Q�uv�:C��.5��H�@mw8� �+�OY\���J嬨l�����*�N��K ��.ƕ�v/*�~��������O'����z�����A�7�0�Ck�|�n��yA��ek�>W_��܀�嶌��Btͺ�b_�ω�.�@_�4�U�����GiQ�}�0��L5=�s���5����·2URe�6�'�/��ۘ]ti	��0��|��鯮�*�6��V_@���@O�B��!�vB��`[�us_��"f"b�,�����r�x*	�7�2Am����U���!�%����5�59�#2q����^�<�U8
�(0�D��(��fp�WQN��#7��S)�܃�P�;6��-ɠ�Z��D�I��X<���4b��SY��o�bK��3a^G�]$�����Ѩ����S�5g��S-Z��zw@"Zx�|D#���Q�.(�g���l�M��P�]���0	�.q����c�#Ř,�� �{�M��o�Ob)~#K|Vw����,g�4%�o�r���kF1]iL �����c�̰����@!�q��_Qm�
Q���ҡ�U"�UX�66ʱn�`k�/�Pfj��BB�W:,����_�C���� ����gND���֞R&�^����5~�o�̰{K؟�j�/��՗���s��:���6�$���J���<S�u�8�Lh��s˗��Գ!�sgn�d�JT͌�bx}����b �>2?A\�)�Z>��ם�5R��B��*�1.u
鏞'�)��3~��>^����M@Q��q�|����- ��p�4����
�U�X�*�@P�Ȩ�w�H{r9=�rD��P��^�R�쎺6Վ7S"��|6�D\�OdqA!C:4Tp�cNEp�|��\
b�U�Jn�?�Ld+[�ޟ�k��Q�䏄�H1�:jR��!��؀1^S8clxR�[�>�`�H��;Ҝ�Qk��e����zh�Mk��C�����y�R����3A���vHIc74�&���zL(.#sD��f��$�|`�����7���r��d�I����>٫����Z��C�%�+z���I:��dk�5e]+5�TN9��$а5�"��e����H�9\�.Y��9�h=P��jn�t��s��d��#`��W���������B��Lq
r�B~��l�-���s���Dء�5�T�A�G�K���^Y��,�3,��Z'?�l�HÅ�v*e��U�\�>�3��b`��u���UV��
��(�2�`�L���̺�?d7v�[�Ve���"�'���2����C�Wg7�Hʧb���w�Qu-_�>ә��.�#~ ��R�.J���N�b�^$x�ɜ�}�͈�I��3��u��b��v]�^���ɰ1������z���,�/�;�뫕��86��`Ҭ�c����ˠ%�BCq�I�A>�(�t��y��8�\�`���b��z;.i�ո�5�!�3a�+��(Gti�wX�ʔD��R�#Ǡ�n�{
js���/�jR����7�C��(�Y�1�s�$H��1�Ȱi�<��o��:���]ڲC5�YFOL��U劅7B.�4�C�Z����I�ђ�$;C{����mP����L!cr�<5�j��J+����i�"F���Kto�v����xA��8w�f  �Xh#�^���ǡ�b�{A�+.5�U������ }��}���2�Ood�\!
�z��!_3hx'���$��>Lo���Q{5 ��:t�̯k䓾�h���Ep���8R��8�2Q��'�2��Ǧ@f��䳪��d�xɬ��<W|�F�>�40ؿ
�0n�$�\�i<$�[yR��7~�X��,�Q,4K��W�/_�5�`����-L�[�Iׯ����(������O^����菥�#u�e6����LO��Z�P՝�m�a࿏���͛S@J��l�|��=�!3inV����b&��?��ۖ�ϞT��*�싗�H~.)إ�M{f��k���<��--��75[���~,-����%-C'�⛎҂��b,�R�O���2��#�i薏�f/MX)�g�\g'���p�Kީ��l.�9���o��뮹��uP�|�]8\۞pz����e4C�Q���=7~U����s���4:�y�}i2�*��E��`5�~�� �6ܟ�x�(8���]o�87�w�=H� K2U�X��'���O3|$-l�sۨ�(���J�����k���(�ϹB�;]cl�<���ܨa�ܰy�!;���)���YRR����N"�o�$�6�"��D[6�ڃ���8,-�8�3v2n-�x�j)����1�@ˀ����������$��L��.[�ӓS�c^ �4+اn+b��DWɚ��ys�6y���в/6G�ҜA�J`�� �>SNX�ԉ#���S���Hu��:�"���	>�.�UIX�ܭB��Hr�DC��M���cC��1������I�~o������,�~��_o�3��$��;��/.̒�������������c� ��;��ߪezz�]Q����F�ࡲ��)�6��D����8�,��}��@��}Њ6��Q�;���E�ZI�{f�Y2o�C��TV&O�D��Bw�u�_#�Ag��<ߡz�`��#䤝#�dP��[��)bP��|z�x�vؐP�����@wv+�mMV��v/�����<�x	J�3
ܼC-�dA�"���}�����[\�qQ��\��S���[�y�8����`�䟾�$[q�q >��A��]����0��۴eX����
�bo�,��f;ho TvmV3�[��e�Q�2C�W`�qfɨ�`=��6Z�r�I]9�e1G�]��y�)����᭕��#i�j��t��<Q�P���?��az��Y��FC[^���X�'�7���j�W������2w8��ůN	>G���S0�:��`G��K	��Ͻ�o�0��#?�&ZHZt�-���:���u�YY�}fw����U���n�>��W5����>��$�
d/f�5�<���i��]�YX�Bl�;���0E�~9��M���2-}��?|d�p�����"h�F�0��?�P�.aMiv���,Y�8�u�ߴ�{�Ʊ��D�G�2����?(�F\���I:c%%���'�.����p̒;�X�#c��D���N��ē����2_}8<��xtF��IrC��s��[/Р����E��;��s>c���U�+��J���X �´��U!QVE�n�0����?'��Xg�/����0��̭����1^��@�<�?N}�Q�)�ϵ�8fΒV��6��P@�f'���|�q����!N�� љȳ�����ڪD_���q�ZU�	�N��Z��XB 8�Č�X�\g�B���Z��	?�g:+���a�ۍHU{�p.�O.5�͔�+yn�X���_A��]��r4��"��*��>�P;+h� 8_�=d���Sj.>UgU~	�_O��`|UlHr�ØLy񣶷�0��"�6,;�L3��	|��/�ܬ7������๿�?���e]P�Q�ӿ�j<�,7�:�F��֬�n���f`_�+Ώ�19�5���jӣ��"�����Q���ARU�!R���pƨۍa�����̃z�wCw�L�'�4���`���U�����X��?�,g���j�G`��0� ���s�����`��g˪��Ӕd�^�7sXp��DB�i�;�������"1P��$9�6�?��nJ�m���c2�*u_�m��}t�)�Ւ �]�~�����6��y�ۑ"^����q����^t�SS3d��~�u(NN�`6�!�o�ί�����fmģ3=���ڟ�ח��&��`n�}�Y�l0!�`��Q��=��TG*�7fU0��ԃ�yh\HFLN��(	En�N���^�=������3�l-b�P��U�J�ݕ�U��X�Yc̓8�� 	�PQ%�p�G��n������$�(�'�Vl����T�Qy�Y��	��B��َ�c��>����qv����]�C*�L��%���׼BB�t2O�ů�f�R�끵�{�<�m+�T��[�����C����r�.o�Ʌ��:?š�Yg���1
�ޞs>����2�_��ПFE+}�zMǷ���b�,h<�pp��_U��ؠ8)�nr�.�}c	�F#Y\3%W֜�;������Ivg��h��'���\���M᠙[�R�?D��:]�렽Xj
����A��7����N�ʶ����ǟ)S�$.���P�wJ@\x��0��,Ӳ�Ά&��Vg���g��vu_��r��d� �.p>v��3%H3�//���W�M�c���
����{�(�Y'���1��=Ӻ�j�d��|I� �/N_���/~�?�M/Z��m{J���\͕�=Ө�T�=/���aL�(xy}��W���U�1y�`\��qց�Q��"���K�-��]W�S9�<���BO���O��ma�f����-'�AU����T��T�t��n�
��p���f��Y�b�>�P]��t_l����f��BBM����#Q	?^j������c-7�'�mQ���u�Ŗ,S�z5ùG�|'�� ���x$$�n�_	w�y�A����03��E���
�^u~&1rL��L?s1z�,&�ws�D�+�SbIrk.����e�6����C��\U�e3i���u�]h�@w��o3����.q��e|�f�ӛA1�p������-�Zz���}mHaC��1��tW3b�ȝ�����o�H;�9�<t��3q�2͌Ƕ�_�qX�.qn�탦�� �|�~R>��33us{�ܲb��(m�r_��:�z��u��}�}�{Wm���H~�\�⪴�N~9+_�C�hv~D~��FBԶ~���wN�0lx������3�5kM�J�x>,zڎ����>���r�P21��� �E�OLI�q��t;�
�fl�b�<��:j/�����?X%���P Z)���<�	=�Q <���՞�fu5�ZƖ��K勻5�F�in��8q�� p���r����S77�HF���2�f��;uNv8��X3W@?�9��g���|�d���:�fA��@�,�eV����)�tt�Z*���Z��Hͱa�-guf\AsEjt�gŒR�'L9�gh϶*fM��=�(O����Z�I�H��A���E�k�F:kOB)W@U?� ����}�^֐�O��*���L�Z~�=�צ��Y2wG��rWO����6�6�!i'`��⡨�V����N� ?y��AXbn):-������`���l-ou""iY+�ad�ǁ��1Tp��8�}%����.Վ)r���᠈��)g.Mp�����p�I>�\w�Q!��/h�����av�/�%���j{ϣEm�w�]I��ꆧ�9U�4{���z-��{:Z��湚V���j[(�T~�"�KR���z�������M��Ƚ�Q�y3�M�w�[h���l$�4��g/:
jg��ԘGEɥ���Ѳ�J��](gL%�`O�*_I)��D��3�|j�~�a����dPQƮZ�����C0�F�62��~�����z�5t 0#�Ȋ��>��i@Y1��z���DCB���K	r	&�c��GF��=J� ���)�[�YG's�^h�ղ�ÿ�k�.|H@ܛ���A;z`	�����Pz���,�#��@��v��!e�V=۫翫$�8_�����R����e��Q�#p��bCgyt�d;`��<����Z�>}I �r��c�)6�c'�h�ߩ��@���a�:*���6� �E��G�|�i�Kڼ,��JDu#�:ZIK��졛�j�5	��iĎN�s�OE�ߘ%���9c��޳z>l��4�!�<�T��&�t�U�k�Bed�[���Ԯ�k���߾4�æB6�����N$,���S���H����CIu����
�+�2���=�V]~ �	'|ml�T���a�^tk,\؅�mm<��G�	���_���j�|���r����~��a�m0||�GK��Y�
��$y:SWA�J�`�פ<446������
���7�wjM��Zn�ɫ�?1to�uλm�����N�k�3��~��	�����E�]7���~������Ѽ��Ϲ�,�lߚ���6�8�i���V_�'�􀫇Q�˫$ܥ���QB���NG��!��>N5{M�&8���.MCd���yj?��7�f��%~%O�e�l��r�jG.㟽�O6zS-���k��^�x�s%L�-��bB��L�� ��&��b"�! ��������&z��6p̯�׹�W�<�UH��\V��]9�j]k�������Z�<��"�LrM6�8���>By���Ѥ~Рxy�6����޳�������D�W�zv�o�5����4S�7�_�%Z95�Y�Fc�<Hl�o2��wR����R��8lY�}?,L����6*ز$b<��G��']D:K�����J�z�G](�
�(ۻo���S<C�\k��bm�����F���^\��)�E�U'��ꩻ7�	j�������]yy�+g������~NKe1��|'I�߾<�$�-z��s��l�wy5���c�5P}$�t:N�0�"�?�m��q$�K97�ed*�Ժ���[a��i�w�XB��,����HB���v�nXQG�� l��^h�1�az%��S��k��<����$X�G�����㬜H�_?����%�ۅ�i<��7�YsA���D��kŠ���,�\�"	@���{IB�x_D�9]���ba��\A�\��|��l�����@�[zM���9�&Pf��z�X5M0��^�v���,�>'�,��S$R: �P{u�lѫ��b�L^!������Kq��C|� �BjZ�v6[X�#yy���f�1�M%�"F\Y����!��S���K3Y5�SpS��$k���C�F��"2�Z:�K�1::j������_;U����;my�����m��z�,�\G@7���W��a|��z���Ǣ��m���~�+�	�zq��SJ"s��{�g����SB�ˮ?s���)����r�I�NyY|�
���F�wP^�B�q��et`�ص}�&�!S��I��G����W�eǍM@�96X�iRQ�kN�Y34��rʊ� �j3�!+��;H������#]#Xs*zI>������_'m�+�o�ר�巢u��ڄ�^ɹ��D�O�I�8]���� �$V&���a��s���<�s�,�D��;����%p1�q��{v.(��k�C�$���v�%���pm�WB��V	�J�-�z�*My|�	����@���H�.��a7�DO��톔�������c���dq�wH�q!��EJ�(�9�J�e���j���u�{m,6�!�YI�Va^g��
r�d�s�/#7�$��rƲ�OO�4���g�5_����/��3U3����Z����XnSH~�]6q�u(����&L[��;�0؛[�f�j�#l��~P��p�B�4o301pMr��42ӭt-7ܻ��P9���9
�1��?�␄d	��h�sb� I�p��{�"�c�h�Bt���+�M�lu��6�mq.jl|�j�5�h���`ZL��iO�9��?lKon,���[�AI�z�N��"֗?p�DC�	����W���b#���#� $ :5���S����T pTA��� p�}����-7`B������"b��9FH�-������"Ao���X2p�O���_|�bSZ�u��i	��Jp��Ļ�S	����������Z*�7z���]���=!��S��F\�kQb �߬��k��O�%[�Xq�z�DR�t�2\���1?1�J@�t�A�*����cD0������]�F.�|�"y���cb���1���i8���?V��NGv�������ʧ����J7��=�3V3���υI��mᨰ�� ��!^�%Yz2q�9o�R0��pj�2����/ӊ�܆��l�>�8�m���9N	礥�96�Wq��ρ�胦�u����AG��gh�0#��-�{�-���_��'q����3��	�9�4j�$!�Q��h�sB���ak��?שV�/1�,~���,����VMn�\4!�M���_{й��%����9�����B����|�S<вBW���Yy�`Ul�;�U,����p"��גW"�fT�+"pׅ�;� �j�������]n����!�$�c1j�i�31�������uI(�,�n��-�R[qz޵8�����������x%�o�!��0��asc����L�S�Ȯw��*�rζ
���E����	fE��K~���/YM9����-�� ��{k F1���I�5-��0@)8�^O�O��Y��>�FR.i2����r�J�G�*ˎѐ	$�,ԑo;��5׶����]�$1*O(���U�A QaK9��ԩL#�qp_�x�E���ZW�¢�y*� �B%�)Kwy�����tq���՛�]�1��*K�o��c\ IrɼH���느�/���h�<2�/���vrҏ���G6U/A ;�'� �B>q�m�fӄP	��)�w�^��$��@�Hec=��������r��'n�/�x����D�e��EB0�v�8��↲28��gq_��d�WMs�
��y)����t�ec����Za��P�Š�Xjm��_�{JY[_]'m��b%�b�H܏�C�:�M�D^�\/��Y1,D2���[�_���)����"�-rz/�&Mt���cg�4�Z��e]�cfD�:��=L�����dtv���,)�vޑ�]d8�+��	P�_��SӇj�����F���=��9[.����4�q�<��e�@գ	����XI��(�T�bU���M�ԯ��t�1��'Nk�k�sli��s��N{7�����)e[�x��{U�]���D�q��8P���δ�o�[j�o{��0`���s4�g�p_�M	����V���:W�m��,C�O)*8�?�F�h���� +�\SpM�U$�iݯn�����@ihiJ��&h�vfX�G���"n�D8��2�G�-sL����V��ܭ3t���q��Dso1ɸl?�ϧ�`������j�9�n��ۘY,���D�p0'�M:W�̂6�0�*&��V��w�9w|�ʪR��(�����Q�U���;�����˅�>a��$�L�ZT�E��m�!��9�q�_5]8NT��n���p)=l�E��ٽݯj
L��X��n�5� 3o8�y,:�}��\��]�8�"���넼 �.C57.U؇�[U%İk��Z�����C��_��KG$�5-�/��*kS�����t$V��bN���pπ��YX@A3SVA�n�-�I�~)o2CN'�FE�m�x��"(b�*�;�%�s"T�+H�L�R�@�ϥ�`O�*�.�y(E��,�1lE���o0�\h�I.��/CT��l�P�A��X7n���\MB/rw$�(�*�9`9z���}�+h��[�`H*��,�j?!����݆�Ǳ��ۏ=���g ֎�,���$@�?��c����V*�a�q� g�b&H����?��;���S�*u'��bG�Ey��5J��ktב�T�����^��#��n]�����$�����s%[�FAţiC��G�+��!:�\z�g^f5�e:�+�͵�����:A�Oޏ{����V�o92; å(��1���#��s� P|���7^�����A��o�4��'�P���쉑�fо�l!#�ߧ}����T^r�q�^��5wDdn�@��1�u	��C3�љ�n)0G�S���p�6Z3��פ�	_��� �ڞd&�f3QP[���q,w��7i٫��Ɵ�;3�5ΒQ�Q�X�(��Yq�0wİp�?T]Ӕ8��C�[��P֣� z��'6�H�״���xil�L���:o�lMk1?�??�������W�7�"���rc�zK�`/�7ÅZ�6��"qr��|���<����P,��M3�Y�s���֬��ø����:-C+x7|�'bB��qJU�(�u$1!=5��G��E�o��IW��v���a�Eф�+D�؀G)����~����ԡ�����c�;��������ct;�>(W����5g"ǩ��M�ku�"���1S:)����/�g=�J�IA��{�t���~7�0�ޓ&���[A.Oo�S�kw���A�@κL	}&��Nj��a=�`S�x��kX���@��b��S�X{Ԁfz�`UQs����S�����X`�j�'0%3oj��W�]a�]�s���Jf&/�G�Ӈл�v���`��F0v"<�g��da�F�uY߈���!���J����Hv6��xnƽq%�ڂ0�J���t~Rw�ׯ�7��^���%:z�g`q������k�a��'_��Z��=	����
��
�Ⱦiꃇ<٥���)��\{�z~D! :Ӏɲ�t���; ��&$��!�
2���Iz���7�{�����35\�������E)�W�l[;���ثY<��rc�z�诬;��d<'�0�؛7����F�j�2�CE��f.s���R�����d�P�OB�[��m~u��h�hm�[ ���L�Q(X2���Za��=?ؠ�Cʏ|n�g\�ד	נ���-�W�P%D���m>E���.0
��ش�[�k�i��Xl���-+8�@�f��N0/�r�n�������`Z�����y�}^��Vč��{"�/���= �h��p.�lP�&B�A���~���|�bH�󠽲�L�<n?���#��8�r_�rp9wS9��N$
,T?X��e7�ʐ
�e�x��6�^Ŧ�U�{AL�������G�2ˉ۫8���AvQ�~��C5`����Ջ�9�1����#��G���ͅP0��'ťKH�=�p�[�춇��������u4���������g��!R,Q�����3L�04�Q=�t�t�;�3j%a�N���m_E�O�枫�I3���]���X�7.�K�Q^?@ެ-��g`���g�G`g��N�l��?�@��=U��B(��?��a���sǃ<#b�q+LLG#��h�F�0��!��_�R��A�
�i�B�Vr.�na�� P&� *�P�>�W����A@RF:<��@�FV^��
h�S����<��9�RF'ҋ��9굴B���׬|"~�Q��U0��XN�5��p��.D�^Z��� �;'�A�$�6�s��h�Ɉ\�R��'
�
j�:�%{��R
����.��u}���2$	����
��x�6��ߛ��O�.q�@ǐĞ+$����?�������7;FD���bm��}��B5��HP�r抈ї���:��M���)_�/�@�2�(�爒%
���C!�Q>老M������2O�!����.d���$gX�����4�K�Hhjz s�D�Z�LUgA���L	��v^�̊��BڤIԬm��H���p�Q��W������tXH�� ?
{��q���-Jj�g��2POǻ��'^��Ӡ��Pa�ez�R5t"I��$��5���v�:Oc:>�%���I�M����-��D/d���5*<!b�o�ͺ��*s)˞{��Eʾ���F�x������5�%�0�pMwv1�4�(��K&10�;�b�#�x�	R��6i�X�:~�(:v�Y�@�hI�[9DY�I�L;�B�,o�tc���D�*�A�\J��[�0g���j_@+dERut���:G�)�ON��Z|�wJmF�B+ؾ8���r�{z��S������bB�1�ΑIƵ�p�2Ƒ��i\������-�"�e�J&��1��57l�nO#�V�Z0=�Vΐ���i%����2�ܣ��:�)�_�w�1keZ�0x�Q ��X�$=UQ(�q'�z�!��E�yAZ��"��%��������I+�a�Mt�j�U������|�����n,��s�3���`Y��J>g�s�s�OJ�����/Jl7��	�E��O'��B�r�G�-7!UT�w��k�&�WVW�Y���|ٖ��McCmG�&$L�L}�"�T�Ix�7r�9��˞W;p���1Lę��|�	M��垩�V�V��	��M�X�c����P�.�q20\�y������� �K�����' ���[�����i~|x��*�ײ2Nf����������mp^��<�.�n��'�����Y�i�CŒe�Gp�4���f����m%*�sM�ter*\��yN?��5G�_��.ş�8="���G����GVJBE��٧vzG"��^�^�5l�'�a��}-���O���Z*���Y@��hO@��ڜPn�k�=��q��skr�jB]Vm��I�i��=����fp��I��)3!�{����S��I�V�,N��K˨J�(vl��A��%��H��x�[���:i��=�Js��ST�0��?1�	Z��3s;��^�,{ک�#�G~��]�ax��x�X!�֠=$r���43�t|˟ƭ�8�340/�=�wꘑ�8f�Tn��h�w������gy�Ę�<�m��[Tހ�O���Ó	��yO�Z�&��Ƶ�D��魽�=X�V��F�&����d{���u�3s���I6	��G���Z.����$��� `�p���1i�1l�D�L�,.9����n�	�ӱ�3�9��GtA�3:�њ��[���Ӻ!UX�4�j�����b�i�t�����7��~l�9n�7����Qw�pwKk��72T�=]��|KnV�;?�yV�W�[�g�h�.6˦�qK�=LR�&�>Ew�ۙwa%o;�_��C�ǉ҃̭	
�K$���u�6 �20Ǔ��ytF�{ �R�ɉ��l&I������u-�d�D[��i����=�������]�7���/p4�}���[(�5�Y:��rO  73�j�1�|K�I�|(�T������o��H�Y��<�����9Qa+�*F��;ͻ�<G])7����JNh?H5{{�����Qg�;_Ƕ��"��4�3����/��Ii�ڜ
��Y=�,l�Y���t� ��܆��/7у���)�9<�#�g�������Đ9���ǵo��C���_���.�8x(P^���w�@��0����c6q��ϿHg)[�4x�w�,�8/7��?�����#-!���T�|��;�[Ì�)���Ȇ,�Z�	㣓�x>v>����isR�+,��NG��}�HD�	
����v׭�2���j�~�t���];�_�>j�8FG�*hP��򷖲�,�g�P
޹��y������+�&g`"�6;�[��:�,ް��(Ktd��4:/���-r^�I���Bq_7�=�jF�_����;q?پͅ�E�A�-K%x��V'�5v��.�w5��;����oA��02B翈�]�����1$��[cQ��Y@��ifW0��3��q��ݍ~��[C��Ư�>�S��A7�z���+C�=�Ig���s�W7��{L���c�y�;�dG����Ti�՟�+c�e��gkz�����O,�o��)���8�crw��=��.��Z��&VY6��_��F�7]"��
҂.�	cq�W7P`��Rx�O��P����.�Tc:�D5��F�(�賥��}�"F��cԴ�2!�g�8MNO��Q]Fw��:@m�>n�"W�W42�h�^꒎e��6.��b�ۮ%O��An�{֫CD}T2�A �����P �	j$~!�A�6J�����\q�v�j1ŃD�:��/y�����n-!�#���x�4��K�*���&,�"�#�%"o�lq��a)��q/�!���`kWn"��D���Va�s�8��M��O��h;M�^� Yn�hJ�!�QU^��iↅ�2�Iq��AՙHg:5X�_#�l'�u��v|��}�EV��{oY��/���IMK@�hZ��Êt�� +��n޺����h�l�f��UE���lSqv�,y]��� |��' d�b��kFEx��e�	�#���]t��}����u�F{Hi?J�V@:ec\5xs�j��#�����3N%շ&��S0�V} ��KP�%�V�7s�6��]Hd������䗇I1ރǽ�����5��N����&�&��.T����{gn%$��yh]���f�*Msyc�Ec�,�Z�D�V*̢��Djz>:L�F �:�5�c�;q�P�