��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ�����cY�r��|�Έ�bE�(�Ӭ'S����,W��_!�2����~;�T�G䂢(%��¿op��`D�|"�d��L ��GFܫ����h��e`H��.H��ד�➁�,��b���>��
Έ/�#M7�9'x��<�������?��,�V_謏��κ淤ZH�[��Z�z�+���=(��r7^j�ϕY4�UŖ�Ƒ�I��U>��$�v���VM����������+�S5�#�p>�K��-J6\m3ej������*j�	�RS'�ȱc�M������&�,�L�ߙ���^nU�-2�+?i�	�H�V�F�h��ס�h����(�]��,ܡ��O�7��)�F�(���Z�)�kTU��C'��+1�v�eD!���aj�r_�����B�Gb��`fW��J%ZKb��:A���_<�g���rE��(�s׬���d۵�5n�H�A��.�'ć�����ڸ��7=�o1���>������*���gh��'�w���BE�{���#��]9-�)g,�G�2���ǩ�4�#���/YL4�ʲg���>kr�V����3�z��9YHcn61�;:��Z�u}q8B^��!zզ�Y���� B~.��k�Ա�:��I�{i��s3����?��L����32��8-�i��D���NTdi�_3�"�������fg��Z�H`��&k�U���u����g|)Lg��p��n�3r�������uY`:�i�C��t@W�݁t\h�?��K-�̥����8����cL�����tt��Tb U��a��'�r#�Gċۡ�$�^�]�t߾@�z+i"dm�lv�R�&S�y�&C�f贩�Dg�� w8�a��� ����@�+�e���ۄ��;W]���]�U�򟩀`S�\����i���c6���!2��4������G������]5��y��;x !j14���y��Lރ&�T�Z#7Ğ��wVL������9�S����g�A���f:S)ͯX(C��w�j�r�}J?���]S���xѮw��+Dx>�F�>����rFW��+D:��˩���b����f�[M�"�����
3��S��q4~��1��0ހ'/���G�6�c�������g{N�-!��]6�{��/�dŮ��k�Ms.�����jAL��vH�5�B����Bl�"���G�:�Ui;���Ԑ�0m����ؕ�멼�p���G�JI����j��>	w<���.�D��q��.��	��j���'���o�>4s���'����vB�w'�����o��g���"�r*�P� �9����EJ���-�E�w 
��ǰ)���G�3�#`�d��>�I��^�;��f<̏4��6�<�a.G`bpG�3!R�*/R�K��y$�hMK�#_Oކ&�r���M+��S��n����_����������vӾ���c����F�L�S���X�w�6T4>��顋�C�� |�����:���s�oF��SW�E�i��k;|�@bV~S{~t�y���Μ10B)�G��n��(��R���N���2�yӸ�Ő��*ug:���:ހ*�H��w���R*Sw�Nr10��y����6�ҧ���T�g�n*�K2��Q�D)`B�5hU��Q�4y���t��9��72��#�?d�I��vB��~c�t;�,ڊ�(Ȑ�꿚8K��x6k���U9E��u<�$ͽ�����%4�u�2�<W�4ީי��#��h��@�?�RX��B�ѫ��D�VC��:���n�L�N�F���k��Y�<@f�B�M��1���rӧku��ܟ�z��J^�o
D�X;]�'��7��Z��+��Ws���ev�)��aa/���G�F"B�ݒ����'+,{�\�,��洏W�0��t�/���-��YhgN�o�?}�����8���23M��N�[��t��q��[�����v�UI����9lL�F8(2��r�����ΗN_ �*�M�H)�[8� %\dCa�0�֬~JRо&��L��=Ed�_/1���K���J;q!�(ں�؆V�~'3R��ڡm37ø��)�.��aQc��z �Aڿ�U;�&���x��8��i�Vk�������/l�G0%�T�D/ee9+&�
�BFu<󩝳W��h�b���m-z�A<�t�윟-�p�X@q Ƶ��=�Je%��1�h��ͤ�U&g.I(}<����4m����M�ؗ����+�k�2�X�k����	,W�D��x~�D@	B�յ���)$�Ť�Tñ[M?^����8�e0��t�r_�A�/�bZ�JҶ~���cN"��1����֯?
+�#ʄ�7a�56�����Z���w%b�y7�� ���������4.�
#�q�pd�=�j�Y��[ʮ6L��U�km�\��%�m�苽<���B]=�k�A�hN�mC
T=ޥ��r�ŕְ�I?�m!���c����!#؏f)�^����D8�ɵ�8M[b����ȴ�%�s�0 �L�o��á�+�#3۱p�%����M�Q�,���Qi)�Z�K���,��a�.�ݛ�tle���h&�;P���4�8���0Я N���L�P�����%>�~�כ����q���g���Ul�ʃB��g"7�E��?H�^Y㔕��<���o`���]��N��]�\K���&�W�kіk��L�M2;�em�:.��c���=lX��"���QfS.s�gX�i�*�"�	��l'�h���}���#���q�]u�ul�Q�����ae��_��D�-�1��'L�I E���-� n�w�ңp-960�ߏ\m������lKGO'���!D�˛�@�����@U$�3�W�'�o&���^�x��7p���~�c:���l�_r�p�A�k>ON�k���wZ"���O�$(���7|���_`�>S�h1�H`��Y��Bӛ�P��M�mek����n���?����Ke�;*�O�)M	tIEo��S��@����;)����di��&��~ӵ��O0}�x[F�_�Of�PfQ[��~��pu���X[
Y�R� uO!���+��h;s�������fb��(&��_?p�gҴJ�P�������C���%D,*��rM��'TΙ���W�C��(ģ�=H弟��	#S�Hȼ �"f@�oE�y͘�ïN ���vt�g��D-��-1<{�p۴��L��J�L��'!-շ��z7�Gk��lb$jxvlB�ڏq�W!ua��7Ri���Q.� ���l ��_/�➊�j\�hD-���[�����t��N&���e��P�r�Oǜ �x=@/��L�����_l�y~�sE,6�H��>`�N5��z�b�^��_�ԡ���MRބ0xM����Q7��_fi����`M�5�F��m���+��תB���[�D��s�	-X�G�r�ذ<u�B-0G.�w����}
�喽������p�X*V�]1�6�d&y�n8u�h��w�j^���+1~ެ�+�{�� bn�@�#��RB����c v�}�IB�;9�8�eĥ�?}�K{�P����1��-�-̘����Q�U.�,M�
R�..���u�^=�`7���V�������M��^�������[��H���/&|��N��R��%��ʓ���laB7���N#���ə�5/��v����R�����7VT�������0�*;%@�...�m�w�o6�ؓ]��Z��/��������)+��B�)Z���OȨE�#L���0.���Y�2"��K�6�6��e��N3�����ϟ��*֨F!�+�r�\ǆM!�W-��-`����y9FL�c�.]�W�'_0G� 9��8][;ݪ�Q�?�[��m�Y�\ �}���m�%0���z��Kv�sEU�Y�enu�����oo�e��|��UᘤU��[��
!�f�jɲ� ϦTs4G[t'+�U�幪�����G���t���HSu���)%��R�݄�6��ro^!���
�2��ك=�d�/=�ێ*�)���k�م�,�������O��w���	�3��"X�hY�2�?�º*Q��q��9��j�Ɵ*xG����7b�E�<ڟ��+jJ�+�X�H��FO8%�0�r��P���I�^��$���oh����b1�
z�v�����-��g��S�p?j�o�������m�2v{Hgv#F�sLU�V���	J_�<u�����8h�pˎH9����9?�Ԉ�p�;h���+)[	�-Yڛ޷�ȱ�He*�%"�i� l�̳g̗宩1����i� �ɝ)X�&K���n�z]��}�~�rd���:Oy��T�,��ԾYɂY��OAy)֭����?�JC��
V�R�� ��0XI$7{fw"1��|`w���>l��qk�-��a��7��V�J�O-`����C�Ĵ`�&�	z�!���?��v����Q�7G���B�nA�H�_�)�v���v ���]��t�2��)�e���+j�� ���A�T��N>|"��z?��G�L��kX���-���1M�.��g��Yr3y�����(u��B:{�&2j�^�S�B����c�@��
+c������w���A�����a]�cq`QW^�l���0�R#�'{(��2�E�W��kE�	`p^��z@���7���H��@C�B�>�,�xT��MBd�?��D���.
���-3�����B��� 
-d��Fsl���Ɠ���'�N�M���V��t9�o�Ȉf?�x�����
y��kL�����Cm��^h#2L�� �(齩i�Ǎ��l�3�pL5�L ؖx�3PKK]�ڐ�A�"KuHE}�����㶳MT���Ξo�v|'E�w��nC6���.�^���Z�lВVѹ�M���%p���uSXP���4�&�]����aEN���O�y� ���m̺K$!��?��z��y�p��@`	��f6V���e�p��#�߁c�)s��
:d��ш�$	9��d��.�]�����Zgb�~ 3�e�9H�/�{6��f�>��DK}LyQy�1�������Q9�/���N�ȧ���<��\(���a�@Y㭉V�"���9בY��N�"�ӗ�@��6u�xv����pB�a �>�6�`��I�� ��<�)�GHqJx.?3!r���.�Ӥ����r�k~Rn�-s=LD ��_g6����q�)t�Y�-���M���|���szW95F�XPN��Esg�[�1T�pd}�E&��v�v+Ǉl6܈�}����!Ul
���[���%��Ѓ������1޴�1�ϤN�Ι?�vN�.�?d��[�B!��m3h��!����N�!����_�"�ź��^��K.F�.��O��
�K�$%}c�#s1�M	`�ϒƳ��]����4�9�m#E;����%͔ˈ)L���l�����9(����%��5�,	a�Z:SŘ}�ת=�OyGO1��rZ&2�-���	C�Y%E��(��>���BM��1�\��Ɇ)��leɂ�nuj6jl4:�tWN�p���Z�4�QQ��%%B4�L�*]9�g�|��_��Ź�/4&�.���K�t��n�D��z��K��f�}����:��(�['�%��A��9�&���[G���N]Զ`��� '�l���#T���J�A�Bk����:�'f'"e�Q���S;���K7f�.���ڠ�������8
Wg�Q�`)*(j)L�����$�jc6λX^�`�95���~e~�?�/���t�Rg[����s�Dը>�H�:�+@�5�~;b0��[mI:�=��2�	0P�eћ�p���7B��a������`�P���^�K޷����Z����0�o(�+ ��5k�5��ߴ�ķ��%�����Mb-A�L.�/ƺ�D�^����Gynޕב����`�Z�I���L��l�ByXOg����������ɵ���A�D�wu��6�i=o
��ڊҹoW��ߣW�.�p�"G����^��g�5�:�s�G���4��oԲ�F� ��/(p�#t��-�K�W���U�xҟђ�g- ��Ӎ��:Ry��H��yuH��0j#"�N�#\Mwx56Y",�+]HA����~��'��]����?�ߪ�w�H����V����Cc卨����E5���[�`���������0,~���ť�Vp���l���<f��Ly|�NZ�$���_>��?�d�Ė�mU�*��f15k��3,i�7�J3e/���Ra����i�T�X9I�<��Cvtv��{�U�r�"�zo�@vr���\@Zo�M��K�w��f+�d?v�O"�pK]}�B�[1�5�dt<q��?���WP��˭B�*�!�ٝ<�t�'�7���yp���f��}?��N�Z��Ϳ����6�_8�����x/B%�����WS� ���P`?x;(lq4I�6�b�m��GA���l��fܔ&DH�J��gͩ������O-�_�23�|q���p�KsҎ?��`{)���~�&�d�S�j���{2cJ�o��W�Y��Eg L`0'�ٵ��%�V1�2�����]����NZ���-C���#�T�':|�?Bu�pi�>_���V,͙dA�96�4&�*z��P����b&Za�)�5h�2��� �kl �c�o�}�F;V�ֻ��u���.(�9U�j��y�/��r%i<���1���m����5A@��:����P�%;$,X�x����y�C�!�捫!pk�nPn$���PŅ�mE�5�5�phgYb�����R'�� ��f@'�|��G�	p�t9��P�0�y��B�VKO/˖j�̳��BG�00;6n	ȷL��Vi�x ��_��K��$�}�����W�j����1}�w���>k*�w*Um�T
��,��ݴ�� v7�(Fj��7I%CVTS�.zu�H�x��ˇ���x٧'AZ��P���R�Qb$7��n`e�o
��V>$���*�I}�o&UhS�G��cx���8�^�lH�b~���Of���2�7�+YM��(�L7��킹-����z�DZ,B�9=Ѕ�7�jMB����P����UT{_]x�Rt�L1!�����LT\�����N��,S��dW��a�B���
I�����i]t>��h�i����[�[J�ň٪ٸčm`�l�R���i�G�XJ�7��G�ɱg�I[��ڲUe�����$ ��EЗ���M��?���M��x_	͠�7��pӬ����nnh�����S�9������!�Tα˯�>�5r��T�2�M�_z��%W�Rۈ��v�?p��랟�1$h�Xl�e��V��ԟ���!���h�pu1Vp��_�R�)���RB��k.�%w�n��2j#�]��ym��>�#��ܣڼ��\���@	�|b(��r�hhp#O�u�)VTU������F?%'�H-m�˴���d�5�m����=e�k�:ݲ�#v�n�j=�<4ylt
���� �r[��e� �j@�J(1u��RB)�U���]Sv��3�1|���1+����h�rb8b�ڭBlŨ���*�o�uOL#$�i�i@�����ǁ��u>���t�^�8Z�3�MKr��).�4�ߦ��d�1c%w����m��y`_�����@/�ž�~�¿�x����H��jvHe']�=�吜�!�3��{�K^u��y�9������?T=���θ�7R�U�L:�u�;�yɐ嫰�lNx@SBL_���$�~XO��uawr�,iQ���" gu����z���㌘��7�w_�6l�G�\�A�{H�j��T�u����>B� ���Ԇ��f�����\��6.�/��yy��a�T�fY�(���&�.����60�F������l�_��l���3�m��-A�a[D�^�/�9H,���vj��9��d�k̪qkY��'Gue�?{8<����
j��oJ����(kgø�і�,5M�G��a�rGAVLk�9���X-�n��7�}�#h�k�B��]n�v�䗇��ݬ�`� �`��g.��ݜ����|b%V`p��"r�B�����6�~*��.��nn���ΡSh8V~����=D��;A�G�ҪNbX:�0By��g'�ǧ"�ʇy��	���
�h���-RES"G9�9%�IC>�<M<a��6ߦ�q܆�c�?�p��ThA���#!���k�{FMe��k��F���?>��W$��;����c����G#��-��G�`��?����b��k&��m��ݲ�N#�����<\�6�v�9�5K��������ĺMRO_sF�w�$���w���V�?Jȃ����}Ø���G
?n�@��I!������Q�sעNG� ��&p�v��@����R���+����g9�#Z\'���5�	<'P�)A���@��r.�/srj^��D�y��8BM��wQN�&�2Y�z�P�᪬_H�#��P���b7˟�og����ضˁXF��"l���{?ds�B���*F�W�J�%��}c��-��y���"����ʰ���t|�K`�/�˭��,�5�A��X6\�.4��ON�L���CK03]ƂIU��ˌ�oG��s�c���xV��<���R�=tVR�l ї�� ���4,��k�4�`��_̚v�ׅ�؅Ģq���cI��\L+;����K7>&� 7"�n�IV��?0|gǱv_9]�s��i2N�JE���g�֊)ޑ��f�萐s�DN>b�@ϑ�V��z�q�}���)���̵|����!d5��TW�`X0�H�NT�`�͚^���L�X�m���b��T�/zL�.�̶=��n�p�m��F�o��ںR���/fG�r,�Y�(� ���r_n�]��d��Lw�7b�$f��и �?�k!:d�:�JObub��������d�?/yN������^��H�is͚@q��m�ˇچ{�N�#�6��_�E��=.5|9/��J%8P�_�FO�0�����~���n��p�d߾V��b�ܬ�f��ҥ$%�{e��s��r_P����r��Άm����Y�xt��΋g�H2�+�v{�#=��~q$#
>�T5&�~�Mu���[u>a}H A/�M�<	�$(bT����k��+���S�BrZ��Y� ����/=���ׅL�w��SCl���0���q���J��//�6 �@���koz|02~�r��� /P{�(v�}���BӴ�N��=Do>��F�p�<������3��-�[��E�v���rx�F/�D
���,��Ѡ��K���,���u;��Js���<�+�n[x�v����ihx���$��{ضN��z�9�b���s�m[��:
�ݪ�����x��������o%}�62�x)T�@�	C$Y�
��4�@��8����� �mbia1r��_֤�Z���D`E�Ii(�#6�V��������Mx�19����|DM �R���"9�4+ tsݹà!�<_�������h���f����hH�P�#�P&|K�I�@O���L�]��q��.;�δQP1�O���ܼ0+W?z�y���Ygsg�����? � �G ����]�PV]�y@��
�G(���sX߮^��1�ж�r!�����I�lM��p�^��R�����=waK�P�"����8�W�>[� ��!�1�sP�5���6h�ڜq2gw���C�:O�i�ئ8áoP�7(�� aZ��r}'>G�0_�hB�Ա���s�ة"w(Z���Ȼ	GP)mk*!6|�?�J0��"�x<5�D޸�](ŧj�{�{��rp��K��j�D��K�2�v�ԅ��ESgU2���n�p�dz�UK�"ޔ�~c�gUw�]<�X�Xkǻ�&C�K�pС��f��X��3��ڨ�X�b`�K�֛ H�"jT���ދw��Nz{��̈	S��ՙznq�J��v~}�㲖�eXC|�n/��S1�em:S��0*��\���4�S`k䱇���3R��v��Δ�e���>�,�8��	g��@/� L�^�a"��Rkdt2�?��O*�Z��PvӠ�^��T)�_�-:��/��$/��L�"�hA	�`Zqڣ�ԫp<���8�\�`?L�a7f}�i?:i{T��b 49�Tn�#���I�c��g�����y��Wx�A�J/"���/��\Y�o꽁�K�6�X��9���S�pM�b�k��]��Wn�OR��E�`���.�/�����R����b*��,�<���웨WM�5G(��2�|��b��M��e�|�̳��8��g`E�p2�����˪�\���Xv�Xu3��w��,�S�5F�,��_j�o�V��yҦ�Y�����B�������v���x��F�%tb.@�0����?�J�U�D�O;�5��fǏR]�m�`��@+<=�W��.�H|�I�)xۈ��i�1�h��/���e���}�;!ݱ
*&��t&�څZo��¹+C�?I}ޚc ���E����k�A����ËeJs�4��l��'��˛i�:���Մ��F��Y���a#�$p��^����8��磈��sɍJ�����dy�<���������l`ix��Ӿsp��T��Z|�:!������dM���G!�x0�Q;�H_S�k:GJ��L��=�GdZA���en
e�B:e�� ��H{2��í�{5J��Qvd��4�m���-��7��۝>iu/M(Q������҇�#W�����󯣃(������\c!o���Y��������EY��Ē��i���`�Zko�c5��!�Ef7����uFv^V���v�@����f�6���e|*q+B��j�,cl�@d_���(u7\ꍆC��֛@ ����n�����B��AOJ�i w}$;�)�$�.��V@��|�!Y\�Oʠ��G�k��N65�qb��>�����5 ���␊��~C�O"�/�ہ���n��]��$DyH��y���$@&��-�A�׬��L5'�s���Հ݋BS����K��~��s��v����tQc�/���J�(h����p�S��?��1�k��m��e�וO�af��#y��K�t!����*&�t�����hq�<�t0�U�F�b�,�Z�QA�rŷ��7�)�A0���}�|��j%	� A����P�'�5&���G ���$d��+jT����U{y?vH���q܎,6>Ǡ�q"[�.*���M�NϜx�"�� �>NPpM��w���Q�gQ<gD��$qQ�t)T-�5��U��+�~i0c.����w"�my��3�\�Ay�ݗƣ��{�A�*�����ܪ ��#h�2�޿��H�`ݞ1s��vh#dQ�L�`�A:}�)W���ZrB��ʍ0Z��o�>)����IV*��GWd9�y�g�0��Y�m�������`��C�	w�?���IK�o�,6O2K<�A��J�)�H[�����*;�r|��̱��3�y���B���y<y������rkcű�Ө��cU��t�0D�G�������u��!D"B3dC:
M�G��,G������"z��u��/�z4j�&L��u��F^��/9���7����8�7XC�o��2���T�N�w�z�K'L�c,��x�qǉ^E��t����'0*�	�+�B��?��s*oc9{y��S_����~T���o��\��Ĭ�ʵ�<30�n��ßoa�����S�E�;���ݻ[*��7���\�%��ev��|���/z�L����� ��1��'��{ȥ;2	�}ڀt����,� ��:���h�:��v�ש���q�,�YJA��?���-�Դ�˴eyFAU&��^�wpI�'����W%��wը�3��j��+p�Ecbi�.���^�n��3��P2urf�vA�I�^T�3TiK��~5<�y���
i�o�PΔץ�ޞ/��k���}LQݤ���#�V�Qџ�.���M�bIvC'Ue�N@i�B����>K(=P��8V��\J�;FYkk�����*,�▼%}��w�н�����v�����@V`@(�B:�&+�%x�hE�Ed�g?��0	��BT���F�5ZFǔJ3�W߻N���y�!OQ0V���@u=h�.ĺ8f�8�X��O�_�����C\`�IXBVY�(�|0���]��]#\��;�j�Hv325�msC��;{$����|����t�h��B�p�R��Y'B淭j�:�aq�I�x��U��� {�!�4W����v��25�v��f#�^=��4�����1 �����Ǩ���X�S������C)Ĉ���a/Ӈ��IB˛���H��&��#�<K���_�����Dnn��b'c>����^0�РWf7U�Vu}� &mS$�g�ЪS�΁p��"	�|Yh趭D����%����E3��or��HQl"���M����SE9�b2��|�u���`�x
î���_�rE_��܆.���IY��gu�os� 9(ql�m�>i�%=�A� d��f�2<���
�v�i;f� �a�Wc��T.V�u�Y�ZS��>殺�^.���������2W������&8����Ld|���*�s�>օ��+5/���t��^���H�Ez��/��w�1�}��j���&�k������H+D�G�h~I��5�:}O{>�c�:eJ����-fF�2Vo��{�l��#�P�/`,|�7է'jy��q�����t�i��rʿ@��֐��w�V�?r�Ȯ�.���٦a��n������+G��^��bu��
9��|?WN���ֽB�����o�@�ay��8���� ;
>��d�H,bt�r��Cv��&���++9�����U��X�?�ؔ�r�}����nh�+�^y8�x���0��K >��^���f��,��z܈\�L̯i�& ���[�����Mӿ�]T�p�;` ����Sz_�,���1�cS�ͥ����2���	p�7bJ�mC��}�al0ޠ�5��n�e;���=��^?ጴ�`�E�x8o���B�<�����D�>0cʟd#�el!�Cz��Z����c��I�]�L��2]��_e9u0bX��D�&�Ѕ��%6�"��H�h�,r�M\z���o�|M�=w��?ṖO�AS�;Y����H��ź�"��Km&}��֑�F�.P�׉�����W�c�������5��K�5��@-
/��f�y���?u��m���M�ϕ������O+�v����])^qτ8$�m��[�G�;Þ8঑Ɉ�"TR�+f��B�����v��6���V����y��q�t����'������g�����$����).��JR혚�(�^}*�X����#����9��?���2+��6�7���juΙs�f�?i7�%[)�gfWX�W�l���
�;/w�#�Wv|�sS��y/���ؼ���J"��[!�:+o	�r�N��BVƋ̲r����Y�P#�}�)�nc͉��+{����3t�8ip�<?3�L�������T��0y�0��<�F�]-���Q��d� 6֑}�!�_��w=��Uu�`�Q1���%�-)����E:YL�3O��I��"���l2��BZ�1�]4Y0��C��@����$�E �I�^�e�I��!�WOJMd�uɐa�����K���9/�"���u&{��X֎��&�Kb�����}[ �m:�ҡ�}��T�Ò̮��k���30Op2f��o�/7�v����6��BWdD���t�����bI�k�6[����;?�2
jvp�
t��ۀA�`* <�WE���E�0�1�T� ��!�Qu��o+�a�b��S�c?"3�<L��(�;=�Ey�9���J�� G�����х���$`
�-�J ��dVb��4�!Y�@�7�}��Z��:b >>��Sl��H�P�����?��oC�)�/II2H�
�|��ul�E�'[��e2\����rĥά+�!��wg����@r�*�`�H&`�G�h�$`W�8���@�Y"M|mUu�v�2�_{g���,�nx�-�Vs��Ty�h����!�gӭ����盄�ko:A�Β����3>��q����I�e���V1@��k���WT]�2�]��Ϟ�]�>w��ǁ�ɟ	���K��B�����0�?����!�e^k,;����Tz�s@ǿz�
?���:����"��zѶɤ�9�<�����ɺ} �6�:��K��/E�@xu���o��k��^�ߝ!e�@�(�=����xbC]D
�$��h�X�.{��P���@���������Q�� i��?�rm�ܐ@D�6 �Rm�j��)H�N�I���
vz��4^�oD��o�*nT��D�L�C��I�㑒%��{���R�Y(���vcV@�}M�� �h�YL5;��/��k����葜vPp-�Q����]�Y�c�ah&��?@�SJ~*��9��a(��x�u���K��!mv�c�|���,��#w�e^mFo�*���B�����J"�~ntJ�$������X�a;�2��7�ֳ�����?`ǩ=�{*Gi��	�70��M���k��m�}¦V$��[��|��W��s�q���� �r.���b�b�΄Y@|iBWX���5�q�p�*�v��`�e��EWS?AB���|�r\�z��=�;C��|�������<�� �w��'R�'����p��O�N� c�S�*\�TcB�z�7f!��U�6<��	�R��Ew�ߺ�/pzb�ͱAh�����T؛l�& ���g$oZ�4AW�U<�\�����<J���"/`PE�U�Wy�9��I��mʣ�|�- �<��=���Ѫf�k%:���&�����Ϲۑ�;L�P�����V2(�#���l��	��mI���/���������'���5#�gŒh�Gm�*�nc-0����N5`���	�T0�+<��U[;��g�8�>}�Q���x�|���,�� <n��V�>�]3Uj|w	���޺���5���[�8vA@�f��Fs�M��u�u��r� �����n���t��$���c����US��%��}���I�SĎ2_�n2�yQYiv�oB����U�z5������Ҁ�n�3w.���>:,P0�P�}�$���԰��kn��/m��n�*���տ$!��6u�
�Y�Wp���n�_c��K�-T�:,�6���)���*����k�8X�`�pqq����Q��/_`����s  ��|^�,�X`1/b�kf�}�C���ԉ�ەP�i�sg�"��>w�N�U<��<ؽ{�S�-�h/d���R���'Q|�ɪgB\�z��_b
�b�t��QA%���K�{�B��8�#���_�!���Í���{;hf��f4]�vF'\5
���G�<,cĉ�F��(�%YoQ���������~4L�6�i�z}���&)8+�[���MWk��z��5IV���A��K�~�i^'����� 1I��q�a�仉���&ġ������߬v��)2$m��=e���y�Si�}#T(���8�xZ[�����^���+a;�6C��Pۧ��\�j
��[���4Z!���R�[���i�	xA.�\/W���2�
�L����Ie�~�pc�ZW��c3r��K��5�%�:�t�tw�@�I�쨿1q��}�`Q�#e�<@������禌��,J=��M �1��c���&���	��f	u9\��5i�D�e�Y"�����b&zR�_O�*s;�ER�S�p�qu��Tu։,����ܟ(�6�6������p*�A>�T�};U���@�V���W!;��m+^�!��d�Km� �]�X���)��ɟM⭞|�}�=�{����2�^����C-��d� ���V�'9��Y�{�{4$��r�i:rq�)�CV������?=��ח����`��~�h-��z�;SVxxh������t�In2t�L���δ-+&��|,��L�G��.���V	n��(�o�ƨ@���u<X��PX_�|'�o�X�޶�l�nP�5A�/�r�2���c�u�.l�}�W����Xƥy!x�fO`s��҂|���P�/��A)oC�T�+�֘���fEIXD?hq蔐���z�p���|��{CV�3�iQ�آ�,��w��w-Hk����<e�3(���{P�~��;���閕#��W������"�)��K�J�_��TZng5���%A4�W�8�P�·�vO���w�Zh%�=����s�|E����6O�c�@��l�����tR�[��g��)���u�����3��m��lO��z���~�U�=�~P��,���8C34S�����hX]�*���Tq�Z���i�p�Я��JԘ�u��/���W��V+�ˣ�K1���ΝŴ�CJ>�I!�����Rǿ��nCMP�_����*��3,�7#���f���Mk���K�֙�����P	��Z��<��M�y�SM��B�gNYg�+���'g�DD��ăm82}1Q������7�`�R�~����Y��r���"�]��F�S,����g�mMMXn�7DA�n�j��P0 h�CQ�"����8Y*�p��n<�ޢrDC��;2C,� 4�2:и����q��C��!�������ԋ����e��Z`$p��aJ_�����sdfOF�ιavh�
�����D�0�~�|���S�Y�X@��I��+���S�W��_�"��&̲���+�iz�{K�}�f����ws铅��K���pD��y|��ǢvU�Z���6�r��d"�H|�7��1���3��-$a�"$��"�7j��MWg��w ������:У؀�Щ�%0���ʢ�[������AJo��Sa�14�(���a�9e������ى�'�����һ��Ttri�����~��3 �<�Q�h)r}~US*��o�ɪ�s�;��=q�u#��{��$z,�C׍��o��U
F��X��v.`�m@V ��^��a;<QX:�Ǡz-�`f�|�fP�I̠N��S��Q� ��8��Ї+�վ�w��,K�^x��S�b��ݏ|x(wm8=Xؙ�J�ߏ��K�[�_Jly��b���p�I'Q@�|����$��ӈr4|�o�\�}�l�۠@��aA�.���]��x�H�N��YG���H�����5tSz�-�fP�4��P
4��o�#i�8�G����<�B�^�Vg�W�y�ȝ[+�z}��A��w��veMg�1��"��lZ��%/a��)�����Gw�)G#���<z��%
��я�b�+�:����*�b#�3�70��1��M^X�|��cZ���a����	=�R\/�F!R�7�����p����y��&
�n�S�OiC��s;52d$�����Va�.�[�S�v�3�qPz�7� �^O��(�P��Q����߁\h����[�0����l΄��-C��o˚���!=�'�|�K��Փ:]P?��ue}O�3;��۷��JX�����Q�f#8�T���+b(���hk><�8̿���,T�2UQ��J�QLf�'y���0y���&�[�:��UMy�����y󝗨�&>�XuJ6F����{?����7�"�q��9�{*l�Ƨå^��`y�����������5�>9ώk�|%�I�䓴u	�}���̌���݇������}��R�����Y�v�_z�(-��Sʋ�	,��oW߁(�f-�����x:L
ǩ�U��N���aj��G��@�O����d�iďD�}=L)�;�K��π�1��/�a$�s�����r���b�N�L<|����bx���I=��\;F�\D yUo����9���o�k�?-?]�|�+�Jƀ\�k�N�"���\�m�s�
h�ߜ@��vZ���g��Ε�NG��^��O�g��t��f�0�<~��?��{��ƅ$�\���ui���jA�Γc���b!Q�V "�di'����*����./z�N�4u�&HC���bɐ�*��D��WuyuJ�����kofŝ��SM�{n�jy^�>}��=b4ז�/�z=��x�%��\�ٯ���Ƕ\{�<���@3*��9cRYD�_���s��z��Nd'��8PS���hjپ҆(�4��t�n7e]���5s<�,�U�D�g:|�)��ܰժ.U=�9�4ټ�%v�I]���@�������q�7����I*/�1~���s��O�����>��e7t(HA��*���g�m�����}|��垾��6���e+KtСQhү�L�	���7G��g���>����F�m�&L������Y����ȕ���c+I�i���ylhn/��P���g�/��,��
��zzϳA�d�%�?�j�R��x����"��ݜ�:�k�kk%�2\�a�h�f�&����R�:4��nba��eo2a\̩����ʊՏe����ؿ��G�2!��Q�Cԃ�Kwr�.��`��laj���dF����=��2�6��|WA<��[����5Śk��C���dO��c��~HmF}]y �D5����DVlf��|B�.�0��i��sS�&�1��/@%@�8��1��O��J̤��<��iK̿A��}�*�aqŶ�r�������"]�M�Y^�a��t�	g�ܴߵ�:�2�-ɶSx�K�az�[��QD�pM�6rHT����I� C��}[�2K�b]]��ٛ£�l.��8���ʂ�c��<Ua�Q
�c�����:C�/��)/	^fO�����8������1��)�l�G�#L��[Z���M�*P��@�����(%c��j�kM��E�yq��1v!�1��>�tД#	����.J��������E-o��@MڧE���O��H�8�O�̓���#~ɺ�'ʦFD}�����2�����}�v%��^�Ԉ�r������p�.3��\� ש��j�R\E�
F@�����UX�=G �O��#�B��m[t�d ]�V�H������Ѵ���գ��&�a������C!$�fW�RB#\���K�V=��~��'w!$�Jx�M��cH?�kP�O�`_$�ۭ���>@�kdO��(�Y�Q��\����R��=@W*vN&z���i)^>�x�xCs��!)k�*�a�(nC��cǢk���Zbt�n>J�s3}܍�j���U�`�|����o��*����&�����]]Z��^����-����\P�`pw:�.H������l�f��#zTt���kk�0.�P�A����3��Oې������
�t�<�]���N�s�af�R���@l�R*Tz��-�m������b/B�$�Q��~�*���WV���e�f�� �D�
Q쨏	(�f�唴�Ԫ�R%DpVy0!��61vN����4XM=ҏ4�X���pц���LH��ӲBɲ��rĪv�aI>�d�!Sr)�w�� KOA}
���Om�Æ�E%�.U�ۂO�nAV6;$�y%���������6����Ix�ie�AG/9PH����[�O�>��VM��9�2���_�-�#V�t�7m�ؔ�|�u�tR3e㧟5w�[�`E�+z7>kE|2�![$;����������R㒈�N�F5�Նw����:�^�~��*�*�V7�d�bM�>	a|(���y��s��N:֪�;d�����@]p%iL^P�q�K�H�j�\V~RYHIbt�F=Ut3��L���z��5�bڲ3�:���/In��W&?'�@�����j�����Z�[m�y0!i�RD��#
 �����ҋ�	cA�7-'���ZSI��J�Cy���H|0�Y�"�����kҊ"����rX�<����ʌ����}�mv�d�Z�޾�kh&A�q����b��� ��u�>&���7�;���
�&dF��[�\��_�HSpc�]�#|gBqv�Ux��� ۜR�7��/�6,���I � �1))>#��*���jG�7{�j��c����gOqg�٫�Kt��w��6m�TÉ�44W[u���t�|��f$\)f���dw_KVH�a�Y�?��W�0g��Ǎ�	V� 	?��:����_�"��X�YP�f�8�b�����h�Î�Y�W�"���Wh^!f��[1L�e�2-޻h���S��}C��UO�K����<ݖ��Lϙ�&���EJ̤W�9��u���8��s�R_�!?� 3���{��I��Q/�/��bu�?��r��E�TC�{?���(�v��]�7��!�)�(�'ƥ.�����@T����xe�b�����[�g4�`|pz6�|��3_#��'��}<�W-����^�e1*B�u�ȫՏ�궗m��x�s}rٕ��=��ASt��8X�xY3&'J���Ch�|3���[��oUyF���+��� u�1�ˬr�E;/�N0�y�&����+��⒢�ȃa����ѕ�d�wy�yc��y2�5�V���*�!��oͭk�8W�Q߱�d*�` �7�-8��Sڹ�h١:�	;��o6�Z��肅b���:Lp��-��Ґu��]| k/�Ǹ�2������MBћ���/�4�NT�����[���v:�ߓ��?��v���h�c�A^��m�̈́uX_G�T%
��h�*���#hx^D�]�����PH/�����/�������Z����.���Y���q�y�H}�&p�>jT��K��W��>����f����5(�����alW��ȃk���uf};�	kϗ�O� h��A��*�F��Xms���de G�ز���4�Ul��aͨa ��Eb��Jl��-���f�wE��+lh}�+��&�񭅵��OG��b�9N�*���{+j?���� ��Kg}E�C��s~� e��D�_���J��/t�~��&�N0Q�!>M�j-F������Z±��Iv���ǔ��J�1����a��G�[{giT7�DWѐ>��2|����{�����D
lP���q���k ���Yǫ .+�t{�o9nM&��[#k"�ǣ��a�k�`,�8ٲk�]��?+�ƨ#��uB@��K~�I�����)e�`� � ��md}��ʎ�1��IǷ;bV�hm$+n�\�-�s���Q9���;�<^%��l��_��&�V�J|�h`\e��d�Q��hI���/ҫ Z��'z��Ù��h�6����; �2\2��HDB�[+%����a�g��J,�>��o�b����Q��V�X�2^�F,�����s˴=r��M�iy�+OU��*��D�>*�����5��/7ٳ��}��<>�\~�Ve�����x2c��@ �1�n�=�*��}B:w�{~���O�����O2�Oi���+��ň��$�1��ty��|�>�c���0a������=����w�@dK�����(61��wݫ����M�����}G�u��&���]�*d\�Tn7�7�G��4�p�ɡR�P�Lz2c�8 ���_I$�a�MZ�J.���x���EtÅ�Ftɶ(�ǂ�X�!�Q���A���%N�D^��'��YmZ���Ț�Ų�&�E��������a��f���f�hb4���J�.����ګ��TwUl�!7Z�n+���`�*��T$�X��k�?4�$�/��s�U�U/x�8z�:�-&X\�d����ۙo�>C@p^�$|n!�?�yP���5�7q��R�s�s�hC��'~R{�i��ǡ���/�/��!����GAU�l�ء� �d���e�LҮH����	ݱ�*^Zx��8�9�g�#�y��R
᥄;���u�:jcA�X}��J��g�Lމ�#.�Yk�W�Vl�R�fE�L��_�a[$@��"z��n�r�#%@�SY��5�j&i 7�x�PGzr�j����L(�=����r���w�V��+����pL�zF"�DV�u��98������'�-���7��S^a� �_����(��2��hƃC�!�I�㭩c0O���g��,Q%v�2�W�j���0��mPW������l��wG�A�<��dit5+m�D�6�h�'�;ƃܛ�b�	w�E{d���!���p�S�e�2�ctYb���1s���8g �3��	Ff��+BI���&$���"@��]�bpǏ���k_�� =T[���a��,7_�n�pn
;��T.�nط��8i���&��U	]禔��o`��ZI�$\Y��;!uE�����:g����ɷq�G�E���U9
�S&�������7����V�	c���`�H*������F^����}R9�*��e�*�<b>w�N+U��n>L���C��Vr�󹜨V3�`��9�����J*!H$���ڋ����P�%�u�m��7'�m*�d�a�e_s� �]�E�p���)���jC2�v ן[&R�?�F�^M#�jE�����o�TP�JJ��А�~b_��Ecz��v��-�x��8<I��9S�x� �rd�D��(G~�j�ԝH�4�ƺŀ����&�P�\��@R8�u�JVBXf,V�c/M��O�W�^�E���v�wM	��)����|�6�1� YK�,�ట�[���,f7�Y���^[��/גij��5�:��yAgi���жTL�DGu*�����c�t�!�=4�" ̸3������[`����H���"�NF�.:�e�'.w)5��0��F���'c�O�C�Q	~�+�BXt�o��\щryO��o��.�^�?�`2(��_����Ӱ�e�m͑��O�Tz�������	�2\7\>�~3��Ƨ�������m���褰�5K7�:�8�~�J�F�M���9�W�ܖ��Ţ�'�mi��G�+~�?�G)��K2��fzD�cNvl9.K�	�H��QuѮ���$��O)�p,�k�7��o$@ﮫ�Z��n ۗ�0 YV_�R�R4�Ql�e��
���z��O�$e}b�f��������O��gC2�t�f؝�B-P���7�Sg�jb�^8>�S��SQ��b��}j�|���!\��W,�%c��'Z:������NV:�V;����ㆃ�{lz���(� c6F5�>�ldG4�[�ڞ�
zj�j�P�2H0�d"���>��(�C��H�q�]7�r݉4VRR�(����}�PG��7�vk�7�j�ݟ�j����LM� �Mx;��<�h��� ��D��`:��q�G}v^3]V��{?cӴ�Һ/��&��]�G͢�
��C�E��2�ox���"p�bof�� �a��($�u�g#��h�b���G*���;����_
��߯���7�x�y}�������)�x��M�"n�j��g)� Q5�˙)�c��\��)N�?�X�1��z���t�����vKN\g�2��������Oo�a�Q���[���3�B�ˁ)�����G�9��iN�6Rmgݷ�Ů�GΫ6���"i��
�R�n�I&쫀�sd�����ޠ�h:��[Mw�_����2iK,3�U};ql�q\����y�lski�Pp�Mqc K��*�M{/)x��.�p�2�%�Fﾟ��b{��Xcc&���(o6�����-��h�#Q�?
�����R�����q­����E}�X����j�,�2�~��t��AY(�C)2�3[o�+��Ĩz��n߹����N(0�<?�:$�U�Ȓ,"8�� 
%6�o�$b�j�7�������zl�\̻sɲ������a�cJ��c��h��.�+���C�]YK���wz�_�>��lP�RBQ��ī�mѴ�4=nl_�jU�I�۞����^K�m�����0q,�},[��@s�iޓeCqnt^ �ʂC�1����m1^���a������܁��|�$P[�׎��DSG�^2��mP�}�ԟ4�\j|ݲ���胘ʃ $�G�-%e���2��C�t�I�1�}�?���>�7k!�ב���L|���V*����* YP�4q�L�U�e�V�����Q!�8�};"�,��ބbCIL�lmJ,s5I�W&rc���5�B��ȦC��¼Ԋ=�H�:�~�$_����+1���r�w��P�0��f1��0eۮ��S��k�z��S�'Ys�*��F��&���
���8/n������h�SI��[Z���ī�l�/�B�}�u��!�^��!�2��`��ʘ0"�\Zy�}g�9߻}�="��v~.�l���/��`���\?����j�[:Ak��Iyd�ۨ�����e��b$�"���mB���)ך��"�L�����Xh�L���X��`&f���^���8{H�6ߐ����6�7t�n�=�X�AI�ѐ�F�Ɇ�V�=Q�{11�d�#�M׽�_��ĕ��~���'��F����x^�)�h_��nyC��d�LZ��)�[0;�qv��c���#�龜�K�'��b�σs��s��?�r2��F��3&�㞺g�7���H[����J����k���I�\?�٠ǐ��+	A�u��^Ҕ��IO>��Vt�{˺��>n�L�S�E��;A��~���A�h�7���xY�C>=���بE��E�n�wD��!֨>η}Ӝԯ�w4A���*\q~�]�&��q�Rً'����fX�C};&�ND�� �Uẙ�&T6܌㊌��u���ΐBO�,�f�s��$����ŏ_��o���94�q���(� ��۷�떼\t��uu�����w�h3����X_dQ�� n��W�p[���rĴh�'��#Op1�Y;m)B�9~ ��X�����S���U����?Ive��&5��ٳN�1�J�{�Br�'&x��!r7u@�������v �/����J��w�Ii�D��i~=�s�6��c-J8k�ؐפ�D��������f倇���:%�"����&�b�M}]�����S��ɖ��tw �h�Q���]eq�Iڸ�}[La���i9�ɗa�������dЯ��.DYb# �1�ǿ�{/j��8oI�:�	9N����\��f�	c�&��I%at-T8�~A}\o5tHRl�4� ��;!	�:m��ߵ�������C�O����]#ڗ5hm����,�B���LQ�L��%�����׭j-�zݳW�� �r��f?V��j�&�X���zz8���f��3��g����'S��)���g��o�+�u��fq�C���#*c������S�ߠۘ��e���`����'�e��Se��V���H��&Z~ר�.>\���Mh{�o��~���Eű(*��m^ś"�BQ(1���}�z��hd�TQ����W�O�*�{EP	V^@byƟ-��XL���H���۸ ��������P�?YQ?x!!���{��È_k,$Ջ5Pr�h��(z��b&C�x��4��p�ܮ )j4&n$�A�q�b�)�$�4��:Q�>��Ox�B��Kg�z���Ie��NM��	*����T-J�q��4�oi��-@4�q�M2wEj�AJo�z�w�gj=��gc_%��,�Êhd�C�?=J&�آO���j�vЮ�d�9E�������y$���ϫ��������I<2,��+��m4y�&ۢ��f�9��c��j{a�>�-!�/5/˸Mj�r��u;����U�&m���.=b�k�P�Ͼ�-(�|:�
�����J3C�Y��~֌/�{��OG��.�����C�,�ξ������'�����_W��������+Ct&5Fɟ�xl�Z�%�*��c=�0>�z�����}�9������a�0�̀q���>���hy�a$a�1��/�Ða��:�4�1>@]�x`}Z��=�.A\.���@P:��j�&��
�{�<�΢e>-
��Y��J�f0�6�\N2L�7�JФ}�&��PZ	� n2��
�Jw$TAB5/�!UY:�W��7��BH�f�ZʬXjkv���U�߾�N-�7�<]���}Y�G|}���x�x<��(�ږ2��Fo'�/�I�WJ)�C�k�4><��OE51����$��Xu <�M�c�����ɠ\]�O�<�#���\�󯊳��qH�z�R9+�mľ6��� o�7R�% _����ԧ>�L ���1^W��2���os,����Y�}���&Ռ�㷒�k�^Z��E��<$]5-Ҧ��V���ٕ��S�����ෞGT������0�%��i���R~�S��� �Ϊ�bڙ�#a{���&�d��\n�=H ���%b���G����T�_?�rk���	R���d���w�����}�����A+{ൄ��'_�r��ͷ�
�@���+D�oB0������za���J}��S�U��ڲ������:��R�d�>�(ٌ��.�2��EF͠�ڐ>U �|�}Yu{��1�TY�]�	w�r�i��k�S��?�Y�V����M�ᰤ�qӓ����w#U�f��^:�W�_s�z@�b�@��E���t��(����F�����c����WD�� ͊��Zˤ���O{��Ů��[.ؚ�|t����Y��  dt�?�w&;UѼ�e�������!$O.��G1��2�Ѷ�5(lh�0	�7��Q T	��,U�f4g�W�ڢ���)�r�1�;�|����J���3�}�����&�.�����$ZQ^`�T����U�k���z�0�e��\�|�Ye�:����
RC�w��;��1�d7�=��Y�QW��RG�4��#��6F��W)���1s�N�Qn�ҜS��,\�����&�C�5k��:1�	��7���>[&7��e�,sc�Bb���ී�L���=����o&�|�b=�9Gfbw�욘�d���� O�4���uj������`*�'�;paߗ�D�ԍn����{�|��=�26T�J���B����Ge�1���%צx="�>��'��@NT܄�LY�P">s9�O���ȟϕ_u��R����^���2��%t�;�b��Hc¯�:�UC�'�Ci^P�!,�}ƹ}������Ė��8�D����Y��׎m��,�(�d��ЀzJz�M/�����F�5�`�6z��K�xnVʙ��Ģ��l��e�pZ ��N�j�$�v�/�9��O6渒A�1��|*��R⧼p������CG�o���jg�r��Q��!����J�M9pO>�����fbꓸ��C?2˙�})��*�����A
M�U��X#x1�`K֘�f�A�+�H�j;����,�����_��]�T{*�V)�+[f���c�΢�_Q���-���F.x�T=�^�u�o�5sX���M�	��`����a��t���;���Z����m�l�v*��D��^�3���;ۓ��l��G���,������LvT�X5J�<ޥaM�D��&��`���j{����JF���{���lL��ո��e��7��χ�"��ۈ.�z�c8���3�D�L���Z���� :x]CI[�T݁P�+��2@�q�hiQP�Fj���m#1��;o(�ގ���g���Ӿ�O>C��%xjI��@W�j��*�J��	9l��oB�<��H���+�;&;�)�M~���oyeq=���������A�8�C> ����J�X��J�7X	�+pK��{>'׻��f���,��Qo�G��@?�p�z�Y�N]h�S�����2O��V���S��*L0����e[}J��K��,>B�|7n���t;M}�#�qph�V�,�b�����E�����N�$�d�r]�ʄ��F���d�>�&v�p��W
P ��R��]�$��k���{��4�tc�5�/��h�Fd��1��cs�~l>$�����|a+���^�������A��B$���5|���Q�7��i!���xZ�@�vyKB7޺ ��Br]`BYvѾ=��-42�Ԉe骙r*�� @�LP�#��~1i�r�%�.��5�ft��T�@��D�a���콛
U����Q���P
���'�	QG�YUS�]24p�G�����!��DAݮ�;�1O9�I�*uD}���})[�ص�o��G����_V�"�%^��'K_�
�������n�OVxv���������4�]X����(Jz'3Y؜!�-�YV��Thȧz��i�=��,f����� �X�DO�,�tʀ�Ϳ�K��$<Hm�e��X�b���@1���K�\2�lR�D�,>������#L]Y(�����#�}���h�c���Ɇ���`���qm��
t��0�\� �Ԁ_!:5+�h1���s5���ZbD�5�h�C�d�J|��A�-�ɷ�-뜦	^��Z�bc�]iF%o���𳕘��Iy[Br_1C~��2��eT�+e�d��qm��� 6L];8)�ܤyb=�;��\"@C>�����ʆܲg�8)��?�]uU��ʝA%&�(�^�3��^�#�=�R��RO�1Y�s\ MVz���MN*?�f�9y�v�ښΰ&[���G��S�9gH`�s�ͱ6�I'�˕�Y�Me�����3��{��y C��S0��\G�V�E��{����N$Ä�.,�����H�7��/��/"�c�'�ͨ��e����z���ac����N��������qA)u5�Q���@��8�P��m_Ϋ`�ރ��L�k�Ǌ��}X��Z���=(�I����Q>��H���i�_�#[��Mϵa,�Ӂ���P���%��C���S�n��%o.�6��Ҽ�-y���}��ڭ>��왴]�8V'��轉�H���A�؁`
姢e'߫�D��t右kK�IP���Կ!eܵWIv��5�Yx|d����rs���K��`�הd���K�F�r�/�_ӕӶ�'��X$yp 8���_��l`?c�	�딼�䛶���[�D5�y_=��2�tq���`P9�RV���^ ��[g|�
j�*_W�Y���)��m��Y�s~��d�7� ��+��=qL�É5h~�}[��d��LJn:�נ�u�$�R�G'� f[�_K�tnK4��M ܲ�V}q�YJK�K�an����f����}�ZM��	��yS�h>f>�A�	kH������vE��!i��ͷ&L��	6��ب��>2��l�'2�5b��Pѯ!���숮k?������1{u���3.7[��c1NI�ݐ?O	��Ԯqɜ�����ۙ���c��"!��[T�"��o��qݎ��HS.�V�\�O�A"�H6���9��n3�K9 �UO�ǬΫgA٘�>��'�@7>B&u��3��D4�}��1��ˊg��Z����7QBsG%[t�}���NhB���,�!�r�σ�Q�T�os�\�ع���H�y��q������WhSWN`P�j�J�-��e�[��*�i�ӾX�`�.��}�O4k�FCMEI�/0ê~�f�gOv�s�=��Y��a)oЎN��a��Nw؎�Ӂ��$�Q3�䞶�&ʌ��;��#���T�RQ�� qT�0�3���N<^w ��ShH���0�m!ҩ^c|iX�]�{��c��x�D��]�b`�O@��|u"��y{s(J�d���e,Q�d��f2n�Q��=1p�s�^D�L9��uPF�#�\��o��G���E�N~)H°B��%�������ch(��v�%�d�"�ߴ�P� PWr��)��,P��b�s�k�0��l�W�l(�,@4��8{�,TIu_�&�8��d�#bv�L�V|P�`�Y���҇\���s&�,zA[8��JK��y�uHF�.6�Th����h�`����'�"߼�fL�cҺ�qa��z��*)�%:��"���3����v�����@�P��7d���3�S��$�>��%�'��n&�Rq�@��ۭ��ԯ
�ܳ�2'���' �����`8K5@mI�U�������;�q �X��&*t��t7�]���Q��dC��'w�4��gfz�f	���j[~�������^jqr���?��ޮ�M6i*:��ީO�eOhyH/+ġ�'q���'�dB��/?,H��feeI�.�rb8[�&���\�=ۃ�~~������z�@���φh�Y?��v��A��NYM�C	<T<���)�!�0�$'C)_�	L>k=v�ϧ���4��W"�W�v�`��#4��C6�ܿ
�'�As]���4�6�׺x^�<��t������d���S<�)�hK)��)�n�5����P�X>�愭!��Y$yfu�:7�NClTeF��Bc��ީ�HRM?\��n�,��l�vo��>���KR��k�V�Q��Ro�ʶ�Z�̗C��/���R�ހ����c�w�����v�/�b�Hc".5����p,�j�՟ڏ{�ߞp����
�{�J�9�~pϢbt�gw~�����
Cp�LI����{*��J�]�����ZIK�g�Pe_L��ā�3�_�_����Eؒ)�z�H0#�ljH���*�6� �ٍ1.-���v�Yy����2�|G��_�5�%�u}�1��q�X��ra�4$A��e}�j'	�y%�*�h���'�H��|*/�?��V���KxM��xOq�8�	�`(I�e�$��t�32���O>#c[_�ؓ[8�b�� 4�	�@�J�A�4��"�Z��9w&�I���i2 ��E G�g��x�Pҙ %�.5�a&���b"S�i���S��L`�;r�� {��(����]>������⤒Ir�p����w��>�������x�U`��[����r:r��uq+�M�C"����;� 	6��-�a�%P�z�r��y�c�p% IM��+����� .Y�h���3�|��D���G�
��_�4ac5�T�*�Ҍ����<G�Y\ B�{ �CZ�awഇ��|c<��Y��0Ի=��ٸ"�Ԁ]C�x��B�2gPC���X��#3�Ԥ_D�&R�Q�Cf��dңϵ�b�k����I��ty"Ҁ��U@b��'*9;��!Tt���φ3�R�ٳ��{a�^iա�fr�ob��y�.&�<V������X�ر쨰���ސ<�w�'hrpC������d��M���_�b����b��S�5�W�}�F�V��ң���/����~Q��i���"`�(	���hD���B�5i����p�۱�P�3��'�| }�F�ڈ��Wp ��>����)����y�:ȅ�R��5g3��BV�r�\�a�DG������T���y�.�#>�ꦂ@��/Ƴ��t�P�uo�ٻ�_k��Ag��ަ<�߷��6�^�E�T�#-t�B��M���9lm^�f�S��`�o0�Z�F���1���}����� b*7�r(q��0��@�g�wK�]|ӇȖ�:���5��'
�jR(]�8Mq#�k�Tl�8c�ۙZtؑu�9��dh!}y|�� ��p\��6m�R ۜ�
}/1;�g����>���I��(���jp��Ǒ��L����p�'�pR_�D1���x;8'f���Ï����c1α��/·w�"�}#��q���O�����_������[��1�����k��G�ѻ1@�Bk�K��:�<?qܜ���r��-���1�M󋃔�O�/V ��~)F���[���JF���f+Q��j�ͨ��L�&�;it�,�I��ԁ�M��
�`����g-�r�aD֔��#��]�B���@��R��I
�L���S�mԶ�K3�Rx�<��X���)&f�hʐ��э��C4Ox�-�'z�����T���I�5NNU֢s��c�m|��Q�e?�C;�����B�[pG��X�JZ���IT���zϵ��)��iTc���3�8r��B_�]��+Y��wbuPط����,Vp���Qyo�/ir�2��X���)�6��x@��tbVU����Z����&��Z�	�S��H��bՀ��.���nRkT�s�_o�_;��i'�%����0A�S�.�Lg�)�1���	�sk% L8���zI��$��I�۬)�?M��*ڧ��P��j�_I���4|G�2o�ɖ(T�<��x��w?��_��9��Q������£ �R2�~1^��*w�
g���2�=*L|�L��_�7[�g���Pbk����eq�o�[$F��p�v�M+�34�P-�M�q�C�����?{���i%�2A�����m��Z@$�C����F���'��E/��,�,���|���Θ�)y�#i���du܄��ق~�U���`�OS�Q��t�����]�}c�r���-�w@�d���)�%�������O5�"O��uc���3q��r���w�yY��,��TF�+�Z��{��<X�j��7�4+��B#ْ�	�*Ǝ.^gU�S>C�!ck��&����άI��c�9G�ܰ�S�9��+���fE�e�d;P.�`������k�Z��pz�Kђ���́k^>&���S�"K�_�H�->g0W�S)��7�|�{c��j-��&�g1N��et8z�|\���=��!#���rn�?��Gg���^�M^4������f�-f�T�S;���?��ܰ���E�3�q����El�1؄0�A��M���3݃�ù���e�[ �C�`e؏�q�5�b/��Ͽ?�M��A(��JMe>tH���"�h/J�]�Eg+^��Sy]y��?��?��.?[dEH����^V�ɣ0����U�α�;����� ��O)��b������r�,�bIE���r�5�	�T.��ph���p֭?�����ASNo4ʱ� ���v��e&�ڳ�B����Z�J�7�JP�ۢq�"���^�ac�M�|�T��9��^�~��7��m�:p�!�;e�u���S8ґg��?�|���C��<,���I���"}k���~��ϣO���^
x�������n�8Ǎ#�Z�b��{�\E)�:�3�00��[�4��J�cw� H�i}����Ğ�wv-0��@�Z�p�c/�r�FPS��9s|�h@?ģ�rX[�������5�1}��X&4�'A5Q�m6��K������u# m���]����l�k^0\Ɍ��{/j��Qr\��S/���9�c��l-���䧀��1��?;n&Tx�"Zז�-�͂�Sy�)�G�^Kx˛�p(:��ٌٯ�lS�c^�&x����<��@�iDc�ÓQ�됊���&� �M���Fкh��Ҟ�v+�����k��lZ5)�+���:)��D�ǭ�!�Qy1�P����v��x���r�'�j�U�*�(�i��{	8WH"H�K±!U�0�Q�>�}����@�~�����>��2��Ҝ(҄�C��\��ֵ��g��iUjA2[��x?�"�>B���6&ޛ�����LC�!�e��ϹT�~�Kgg+��@���V�����	~KT.3}A-������^�'��`O�㒋�w�̠����sב>����=]�{�
^v��)�~Ȱ�\yU���"(�g������s�u1\k�t�D
a_ ��B��աK3t��7))˥g�/��(�F2�n?gل��JM
W��[ _��I�־���H�V�Џ�	��J��>G[7�?�	���L��\-�R�����2�+"���L��6	�}�AIK)"PGPu3 LR9����\2OҺ!�*��e�'�8}�J��R� ��j���^Q�QN�V����H�7��+�儵�l-hU�P���T���w3��5�a<{�I�u^KlO�(�%�hzqb4"bv83A���~Oqh�EB�viPW�Σq#��
䍦�C��fE���~�~��wc����C�d	���ѧ�i��\Sʝ��B��b��o��q��2���SV1E����켫���d-�2�Jo����y���SYRq�8��k��(,��p�����Gu2b*�$�޹��^��#�U��U2!��=��1��������� ��;뮒W���T�3�.�m�>���D�ݡ����ϝLI�wg|(������I�r��UZy��3㶪���,H������n8RZ�0סq�Ez2n��Gi�s����S�h=C5�&��,��a<�k�U��
��CB�'0��"�,ip�����w�0gnw���<f�`�<m*�n9�����0��ʇ�I������x�\�	�ϟ���
�z�U�0I mb�Rƛ�+f,���Z��~UV�L��y�6�Q�+nB��JI��~�3���(߹`&���M"O�*h��v����]f�`�vN��K��%SYo� ��Y��O�.#"�7w*�%lS��p�/i���Ŋz��Iͷ�޺dn���@������Jƍǻ��mۉ�-�U��/%�)���,Uϩx�c< ���!W�c�6��!D� 4��η@Uo�k#v����-5��I7�p�� ��{I��^������8���b؁�6�MW�J�O=uG��Ԙi���D� ���s�Y�H�<z��PقA}{C����vM������+�g�"�������qy�5��i��d"b���Ը���r��W��TC�"����#��5��T�]��;���l���r��ɽx<�c��xW�9�ou�3c����C`��%��v@���av?n�`�i>DG�Es�z�Y���w�S�Y��r���X�qz*؂@����S�ҞdJ�E�7������A|d6@V��&Z@�a��<c0�V��lB<O�o����v���,�n�:����������H@#s&��%�X�3�ܱ?�T�^h%�߂Rw7��6�^ɦ��*g�Ex?\�}�.��A��l<��nMq�}Q�N�s`^.��Q`�&X�b���F.���xm�̈�D��&�1o�8R5�I%��:Q0j������y'km������gǪN��ZF��Q x��n�)Њ�Su��1,Z������!	d�sW��7�<��%�=�ױ�2�����~	 ���п4tw#�!�͡�o^�x���v�G|�8�I����TA�c��r=�S *��7����A!h*}�-�"���D�� ��d�}���5[���,�&TX�Б��Gx�)��<E"M��0+L9�C���M���A_��ZX���eXΣr[u��ƪ��Exo�d�ح����$�qL�wͨx#��1I����J�VRl�z�
0D���E ��3H0%�]��zMS�]��e����'�����6�5a�M(>���H�0�V���^��d��>�j��)�ћ@V��x��ā�09�Z�L[O�����ʆ�&��͐.Vh��a��Q�My�64�@L1m��������B`#��C�f�.?�����DN�
q�ȁ��]
w����̈�q����M}5�Z0�q���\�n�����Mr �!����=R����0�G�����
䯴��G!yq���hz6:q ���2��ʒ ��Ӧ��S'��\�1�:Pa����x��Hp-��YF��F��u?�2��4�͋d0��5 �`�^=_:6�}�N�i{+�H1C��\0mqv�ɼ��nIΝT<-�s=��[�u��m�*0�M���:Fn9ZL���V6�����arT�����/��PUȠ��p�����B�^�P-�Ah�3��@���HB��6Jf`n���reSR[��'�W�ۙ%�wa4(��+���a�&rU������w&fV���p�yQD[��!^�o��s��%���l_�UI���<�;<��h�lf��МW�
yR�|��n��I�H��(d���io����fy%��{=�y<Kf	X�j�3�g�k�3`�%̂�Ҟ��"X��~���yV��k���}׏�f�Ԗ�Tb��^�~�_���*�zvBNg	���1�ܝ����
-#�F��6�fs:^����:��f�Y	�!�d�����栌��('�nV� ƿP�(8��e�5�S:��d��1�p1!�f�ON�II�RC6o*X]��h������e��v�l<^�������U�J�F��G{|�j�Ԅ�B�l���ʔ� 88D��+ў>�'{߼�s��3b�zz�7��y����hD�r�Q�Q%D�T��Rl�����vR��'�4����
ɯ�qfz����(�5eY�1Ʀp����[ɜ�$	]9�p�zUg��N�#�2Ͳ�q�����%I�@ �Z��;Xaw�w��1�k���"ܖvU�����i�Ĝ�Vv{P����$�j�I��ظ�+W���̼e��� �y�Xy�,�P)e�(.Ϊ���x��6ͭ;g5黊>��F�E�wa���|?���{N;�bnM~sKUŀ�Ky߫k�0N�p�[��I�wF�|,�e�aL\��R����Z?�+�y�D�T������zhpsv^��d����F�*�~��N0B����U�}��>�������`��?lvqg��X4ꋑ+�a��X��f1��d%��#ׅ(�8���� ����xW�7z�Q]������7�.#��&�2�e_m@�f�������,��X|wМb1��6�7a���H���>�2Nd��2��?���O򘿜��PO#�QMTL�Pږ |x�Q�,��K�rUC�n$v����r�#�D3�ϗ>-���~�t]
@�����|�x����*@W�+Xj�5��҉KZ\���;Z�Er@Gɵ��W]�a��͙C����,(�z�5u-�������j�$Ԟ�Ϡ�)�I8"., ��i��w2!o��W>Ν_�>m7��H����o/e�����@7�&jX�R�03�������u�GC�0���{(�����Z��T�5����q�Úl�۬��l�.�|��������	�&��DU��,��f��	��^�{�u��n~/��-/�#��r�09��cW���C9(�����մ��44U[�TĤ
����ܭ�̷�@'�Z|�1Sf���'���n����U)D �}�	cLd��L��{���CG@9M�Б;"��Z��o�ɹa%z� �v?P�8�{c�TK]��׻W�Ce�G1�*��K�J��{Uz�1��*}B���F�!��A6}F�@���1`T#�Ĥk�a!�����k�_c3XF\v��� L��!��#�{�M�����8W��
�@���~[�<���1�4�{&��k��!m�6��je��Yy������/�`�I���(����s�7g[ց�+I�e�آ����mڌK�+}+՞��h�irA��g���|����O9:�Ӎ��*�-�-�L�@��L��H�N�tN�VG�}0jF��Uu�O�4s��]��۞�>F�������g�R���6:���������,̥X̨��2���A����k2#t��P�p�OO6��*h����ˌT���|{���qF����G����-�:������C��SāS	#ݥ���*�8�L�^#L��(L��<�F�G��m�3��\qF��)���I>r������t�-��g�r��<�Sw#afp(aN'A�oq-.
ޓػ+d	H���W-���Qa
'��v]��@�M�G?G��R�#��u44NX ��b��Oi��f�ћ6�L����� ���e�ڿ(
�{V�����)���m6R���ؠ%�X�9j�����|Ǯ�w'j��JD��KL�һj���3��|+���9�of`��.�H*�c�@���u##�vj���"]�*�/:%1;��f 
0z8��I+ҝ��˺��f��S��
�2 ���Ra�/��5��Bd�v��ѿ��J�4�L��T���ٻCk�ZT�Lp����몄	�gu���ã�F���@�������ɂ�E�K�XH�jK�넘���������H�wsi��$�l��]b9��]��S��X��(A6���@hH�k�.�~�I\to��M�H@� ��ڿ�R$\�t� ��N#�=&7չX�vT�e4�óe^V���\\nI���;��>����y�{T�e�����[�$���(�Y�U:\�}�;�LN����Xc��(Ζ;�=���e?n�������15]Fu�*�x�;���_���){h��\D̿k�?�K��%���3���XGHN��EQb]�����U�&~���n�(��L�]���[�̼�4�~�Z�h[�Yh.�샮�e �(����3�@.�J�=O���D?R,;��_ahG��̐e���r�U�:���z��{ޣ�a�x���_^ʳ�{2C��
�L���ВX���L��W�TA���âӿ���է����i�jDsZ�����6�7d!�cW�o�V�.5�T���d��>"�!�Wƽ4}��V���N�BI+�m���-�Ɲ#2	��q�!a���s������1�64�ZGrU��RL�	ϥ��跢e��O9�x��7���ۃ�/X���ܛ��;�х(9茍��37$����08ag�#�|y��=-�_����6�שּׁ����+v��"��1H�J�����>0%�l���
��6�iR��,S�ߵ��^`Bѳ>�B"�@����0P��*��xH���z2������b���G�O9)Nv0�Z�K*7_
���<lQ��^�(|R���Z;FA�iU��/�����c7 L+ͧuf�%>`<��=_�ɶ=�J�}�C�1�U�6!J�X��n�!gE�!,S�u��>e�b�"-A�%�9U��|�]?���9�(��a�I��I|��b\r�z�lA����f�Έ�g5�*�=x�?uo�CW�4��9�M��얝�6<��(D��CB�Kˆ�rLᰗ��0:/�}�C|�zTjn{�	�
��'�'��:�~Ek���"�����\���vI�v5���#]��$�?��v��k��u���nOA��'��?��A˶zi�*���Z:�%���T3�Ue�Cͭ��e��/�l��,����Ӛ�u��~���v��]��M{�M"c���˫F J>�Cw釞_�x#@F'i��Yb�a���u%L��n~&�*��h�VroV���y��J�p��p%��^+VX��	-���q��{����@F\_�T.���➋�I�F�։������|�@��� T$�.	)�.�-�Τ{�����t�[�Н���Pl�f.ʔjU�� �M'Y�;X�"R`�":6SU�ǊI%��<Dg(	K$��ȑ��n������ȯib���ø��7B!�nu~�?�����%v5	�E	V�"e��|F"Q��P�b�%�W@��aNI�|�����hh����&������r�e��1��;yG�m���t�͜�ۅ��,x��{+��m����6�/��˾���K��]7\ޫ+3f���ƲP���Y9���-���W��
 ­޳8}��w*t	oO`r6Z�Fĳ��6rQ��k"2g�K�q��3R��(�V['��͟c|�����>#~�{�^�� Z�*(:#���I���ƣ�R�Ѣi3���qv�vZ���K���	��[Ve8B1jG�:�-���dg0�˨�oԴL�(�Txn�}y��~��$1�qТ��C�7����_��V&3��u�kgĝ�V*��(�?ڌ�X/c�Mư3�pI�r=,v���c��ULo�cq�?���?��2�*rr�M)�|��H�~j���Lu��,ue��2�;�h�?���>a㚷/�b�L$E��R�}����<����,ݣ)�2A�+hP}'2�}p	��d`�r���qN�)�4H�0�]"UИ*@�n�\:y5W<˷C�F(���j�T�R�M�|�̽+�)�o������r�����h�	��)3�ޠ����ݺ�v�,�nY�n;��l�;��d����i��U��8�٭�C��'��@�9����F#�����B�): ����&�,�<���tz���&�	1���3��U��FN�GU�����hO�V�r�\���7�:��F�y��+K[�V2���+�c$���!@E�2^�HA�J{�*����Z��8ږ���`�&�����O/@+G[}��"���<4]��&q����,=����K����˴#cop�\x#�+,xS�����> ��e���w���/ZU��*U?w��Y�ef�p[��_��ݹ"� ��F�%�#�F7��nH���&�U��b�?J ���j��ѪI�cň�&BK����W��o�p7�p�^�X�����+̴e���&��?�l�]LOƬy�A�,�������cD�6�C�,�W;o�L7�F߀��8� ���I�>�ǩ��"�?On劺��d:�t��߅������ӓ�f5���ֿѼ��B	O�^K�*�avs��Z0��r+q7uvqQ���L|I�˃�Ć�JL�ց����5Nb�-�9MB�4p6�Av���3S��ICS�D�P��:�ZhWmG19�)��>�dj�|�x(�."�1B{%���6o���'�y������Ghu��k��c���U7��?�%D� �(X���N+���)��jY���^��-�@D�r�Lі�&��X�k���T|��shc��h`��MT������%~v��ǿ�N+6�V�J�y�?�n�6>~ߒ�������K"�`�a�#��Po(?����_�%u��x5��~��-�@�����aﭸ6���R.͎�6��s��@=�_U�cbF����������ˎۋ:�Y����aT�����l�˝H�I����V��|t����� �P�[��h���m86��������b�O����+���(�Y�����
G$�+e�����F���8���6����u"��ujHNg���I{g�?��3 ��}��e;T����(�h��VN�'vu���}T�U���ժ�	QoM���r��5
�hCe�zH���s�Kn&!A#n{�,䌺6����C���Fs�&��KO������Q����c\���U�P�#��"���h�P��gF�M�{?:P��Ɋ��jї��k����dh(��w w�����B��>�A��@%a��c2�bM8Ô�S���`��*\r�1�x���m0] ���LC&���3f�	��#���@c�@&�ƞ��y����D���3B?����`IO���U���0 2��$W8]�mR��P��M�!λ�7���7>[��w��&D��ﵤ�JA���X4\_��T��/��K�r�����6��z"�l�Fn�,��*	hkb���.͘%�r�6Q���	�����!�~-a��E���Cpb+���=�e���7M�:����T7xc��|��\~�A�F�<>���"@�3;k�Ϫ�(],���8)ۺ�E��]MOX~:�H��f���S�����,>sx���������&���/�����^3�:�\"�F�w��)�,���5pIc��x�b ��W}��8`�)Y�pw��6���Tf��gbsv��,�식?��`3��D�йg��|	_/�o�#)jO���hV�<�LW�zGĉ��m�b��ǎ�4N�ӷ����pfa���g�h�m����*��ܥ���[�<����������@R��C�uvv����͏ �"��b�;qз��+Z4����.
�N�#7������d�0[��iU�e0�����e���e�Ol\̰0f�j2�9�XX������D3~�oz�p6s�F/3D3�z?��o-����vD�?%�-$~�{%��*���&���S��9�of!�!��=N���V�Hˠ���U;J-x͵�ӡ��\���CD�	P\���gJ�=U�#mYCѸ�����m�FV4Su&���I���* ěw��33�Ea�����2���'����W��f*�����k��7zq{W�W4zbe�P�$��*,�5�ANYCȄI��[kP��#M�����b3��놪%ʭ� �\F�?�~B�[�e h��dƼ���'�:+Ծ�: �ɱ��ۏ��n;�"�Na���h��gi)�(PlaCs¢�����J�(�s1%���u:��gIR��K*����ͫ�C�m��t�b��U �+��$*�Uv��I(��n����{&�z;��NC�.���+�^��:�8MG>��̽$X<��r"].ħe�b�@h��>$�L����ȟS�=b�����3k!��ԸrMJV��})LcF�T3+D���k�o@�������Y������߈�0b���N]��ll�����5����h���nΰ^����s�`���	����O|)�Q&��ܷ���l�����4!�"��a�O&{B-�a��*�/�{��[CuJ�|�o�m!��Hb�>��sT{�<�:~m��MSK���l�l�ק$<��Rj�����t�:�k!r�w�7�
脯$��5���(����#�D���̿�H�vi�Xv�ך�����d�^�B��xV����ń,og���|f�u�=�z��hE|R�H��0t-��o��ׯ>�Z�7�#t��X��K5)ܸ���7�[:�*�eR�`ЅZ�E��aL�m�+{�G/	���@7��eV��!�01�c�(�7w�� ؖY��Ѕq��=��|��ND���O�J+����]jŝ���Ϛr�4��d��K��7������D�G��\�O��d���|,d5Ėh+3�2�����
x���>\)ҨH�~��OA��=�|������k�{D��Q�xC!�9"�!SӁ��|�s�+I��el��O-A�;n���0;cf[�n��&�B��d"L�f2xyQ9I#��=;vĆ�!R�+8���\U��d��%r��Dbǅs򦱧�d`��Rlh�D�a��}���l3�&<t��s�
h��煦M�{U�	gC3 �{�Z|6����X�Ο�mZ�go�\����c	�v���.����1+�,��uI��y��Ct�a^DԜc<�h� �6X�D����K�&W%ԙ>j���M��<`�,��>�<a��-�8�ww��/T��VJ�&��1U��O]ݬ?F���C��C�����]	d{c% ;b���ט������5�(����D=��h]:W◧�t��k�=u%H�R#H�R��j�m?I�|1%6����Hnm�dwxkSx]�J'.՝��~�+���h��.�lj��	@%
(Bm��sɪ�fA�hEm�?�����1�5����*�c�����yO��^�':�?�sH�Q�ڼ�:��-Q��J+�욤hv���5f���[��:H�����b���`���H2	f3V!��m��Y�����Yd.�����3Fq���Q[k��Cg��&��\CH�^����X���+�mylƅ��>�����Ĵx4�IJЉ��`E��XJ�C��A/� �E��/�8�w}��������Z�&|ID�25�Lb�|@n�@�δ�T�� ���G�zr��љ��J�(^�m�V��H�9��S���x�m��Dj�\���B�E�=��i��`2���:��0�G���G�\Ԙ`����4�W�b1���ݱ�B^�7j�=�]����kL�P��1����Lc_�ϺrBC�"�,�Y&���!��Nw	Qj�4��E�ؑ%AM��76�= �;j3苻����Hc$	�V�����@�q����$����+�X������i���� �5w����^c`�aDl����0\��KN����h��C���_  ��S�i0�����]S��-���"2�)_�k�h�t;���$��븋���=�������E����
?�Vʄ�!�v=�CJ�?pQ�Xw Ǫ�诲6��5�Ͼo	��a�Ԝ���{M"��T��6�e�&k<�	�4$�_-μ��p8������u�ħ8���=���s��+�g��js:�Xځ�?:4y~��eɪ�
3�L��1ԟ�Z1L��Sybq���n���}��ꁾY��Y��;<n��3e�C���xk<C$�I�GV޹���a���ӆ�A׶�8�{o�|�$��U����l!�$ё`��th���T
��=��tR�9	�����ߗo�p��ե�h�� ��حq	`��{px��lJ�[�����gp���~��F��)~]����~-1�k<몣y^K�6�@�c'ڞ:�z�
��_�)��[?9�Ò�&������&$�"-���m��Ձ0<��6S�h��v�&LCa����������S!�G�i�s�����i�\� G�1�)JM�e���C�D���o^��ޏF��='(}�|�r� �������]��J��.������.)�fW�c�!=�ֲd�2�j�;i�q�8��LoIZ����Q�^������D�
���i�U�������!�y,�	8�CxҲ#Os>6��[��%JH�@oT���13}�6�� �m�d��ґƤ|�
-�7�s'^'��vI?�{�~$R$���R}����;X�MPyR �p�k�d�	�KYs�Cv�n�����}�v�+�ϯ���ѹ�ԭH�[��I�<D��0噵����$8�Ω�<M)1M��)��ET�(���X�ϻ,�[���(X'xJC*���l�ш�B90��E7�:Yh�{�`@+ف��a�"A���f�fe�΀�p�|���׸:�%[�����3�(�͌U���̢و���.��I�
�(�ģxC<(�$K錯"��l+?���"� �r-9Gt]d_������&�'KbO�]V����0�#�ԊJg��sQ�V΂�T����@���C�X|�����R�ƹ�`8�Qۢlq�!
P(�)��Ϧ:Sa�8������cǾc���B�|e������Pҧ�kq�'���W�%u�����nd��v�����Y޿l��m辨Rj��)����Y��\��R<�r�-p�N�>
"�_{��xx��?�u��5C�r_��r�Ѷ��ߍ�?iEk�Q�$�ݴ�42t���������W�&Pa�n�\7��O67�t,���l�!d��k���,�Zd��wc������)`���ʹ7҂&�|�����r
8�Ǣ���%���e?��h�Jx[�|�ҷ\ϒ`�*�#����o��/����+]
h��a_�i.��*G,��O��n��F���e�S;Ϥ3�|ALe�Wao��fU��[�����7���O�O	|�W������{w�k�D��<�̣+9H�����L��E�/��7#�[�I�o�ЉF�!�Q&���!��#^�8�v��s=h6h��4#3D�jv�ut(bN�L���w[�q&��ĝ���9����,�0�M��ы��8��k���ݝF�%(ФxZ�P��t���$��aE���Ig��j9iur�y�#j�՚� z�R�SU1 }���sX��m��:�A�Ǚ��:h
��H�v����e�1����[�B�v=������Fy��x��X�8��W����<ٮ 0�cd�f<$ѯ�"%X�=o1"�l2�G�DI.�1#;g����g(���G�Tuuex���q�#��%z�ga;�q�����S"��1 ��⮠��ɉN8qœo��n2]�wRf#)��~H��$�*c�G
���Ct���9�.��/�7e����Q*�9S="Y���C�$�"f:CA�aȹ��j�ؗ�?|�X�wF�D�����xsn
� ����cy�������]�K�w.��F�a��b��N���۱��ѭ�c�8�O�|��m�M�Uq(���b����K��;����n8��F�<����'As�gǸ;��q�ozo�\�_uSĨu�:��_�0*��Lz%�F�@���F0n9��{��M�R�m{����������5�/��J�g�a^�ebF�vK��I3���z9`�5�Oe���8y'�D��ZLэ�Y�jBA��s��I��-�F�<�U��H��Vd��?��83՘'�˒� )�u<�6�d���]���00�.���fk��<�ȕ�ѩL��z�{��2�!�k_��ϟ:�,;������>0
V��?:��a����f���/:��^�@ xY;gI�@��J���9�TE@Y���.�~�7��P�`N2��wl�%��	��:e������r��-:U�	A�F@hU)膷����b���w܄�0q�=�x���l�m(Z�0�+�����Q߶���/$t���� K�����X��a���uN�uUA�e�Sj�Ē?ٶq���{ZJ�}�-���]wf;����v���8�Y;~��{O���a���9 JZ�G� ��v����7+7�f=��+|�r>�ʹ��3ˡ�*z��r��tּ�uf�ω7Pu�G1���Ũn$�@!��O�B/��mWJIg#�Lظ@�J<xt*���/M����H�Qs+��H[?��!��f{�f�1��ś�d�.;�*n���=?~E�J@UI!f����$��������Nc��i�HV�oǏu���	 ��W4�߶O}�����;����9@^Uh�h�$ލ�MU��W,��J�u�[��.�a��2�S`W����!�[����(�I��C�1L�����,CV��Mc����{�����^���'B^dh	<F���[
[1?(k4iM|�Q��;��8���,��r�3g;�&�w��X�������W�H��_8�uF9���L�2IaVZ��k�)���{�NZd������MX�Y��.l<�4�=�\/�ǘ�K�y��&!��nzA8��-[�`Ț��6��<�×Z�ؾuR�`
��N-%p���R���4���1��f�ܐ�i��<Wl���{�=T��(D�opΣ���Vj��5x�˭���U�	O�ˤ��DX��+�4�i�9�+�|��l{	~�������m6at��ŏh'1�L2���I��e�b���\Y��ƚd�^���~��.�mm@�a�Ȝ#��A^�u��%8}&���C�Gb���%srQ�Kk�JCгB��41����|�rJ��R]�wӔzy]��bƴ��{'@��b�
"T�5ep�s�\ĩҧ8,�s9�0(뢑�%��f2#���>Uiy�*��|��g���~�\�p_�A� R�M��ʦ �y�ӆp��z�ߍ"�l��E\Ɂ�WB=2�!3�3�(;�C3�1� m�� u'q���7�*��Ɗ0��
�<�!"=�2�;@����o��c��igGH85.�37���6���F��;6Kƌ-���T�,�v��q
m���G<�jg뿀�Fw��V�B����i
7�A�B�U��h�k�������Ñ���i���I@�[*X� 1�����Jޓ9u5d/))��-�i���J�V�6�FB{�n;\)B��noƺ.� <8����p�@z$���Noj�KË,�� �2/�����W��YcZ��1��k"����T��Ċ�����
��;��o�c%m���|�
֩�¬��07�Wd��l�K�W�ER�Ł��۩��w��ٯ�kn�Yh88o$��}8�(P�����Z)��j��e[=(,�Z��Xkr+RC�Fj�
��.���ʷJ��l�A6�.y'*�f�)����K�1q�j�����G���חRSpn����s���O5�Ug�ΞKǵ5�w���pt�Sv�ynW��i>>�����R��3�z_#�7��I�����N�EE'B�&�X����C*��B��[�҂�[q��/��۰�S|�4�nD�[4P��^=:�����i9�Զ]��uM ��F��Xh�����y>:)�9�Y�gVZ���gGir�BM��S%q$��5���2���vw.��R�סi����:e/�Vf��H"�.�e��'DV��$��.i� !�-�`M�6jG"�%kR��$��f�Q��WN���	@Y�$ܑ%5�xN菴ZY��AW�Z.e�*ō�&�bB�o��I�D&1U��N��ⲷ��3�E{�'�?u\�"l$���@�u�Y2���Ζ>h��t�ߜ���Qoy�i�P\�r���ϊ'a��e�%�E�����Hb(fg�me�����(�y��Fܩ0�wT8~ ȌL��4�t�L \}��R�L���`��̝_�[����%��u�b9d�����DF$�辇�*�IU.  �n���@��d���0uX]*��Q;���n\��^|<��m��$��d2d#������?p8�/�,�8UD�Jy(6["�.sX���O.)��R�(��#��u�@$���f	�YP�x��g�wo�B�A�K�:�U~��S��.hכ�r�r����&ʬ�39��n�z���M�;�����ZO�����c,�VZ�Um��H
гɠ�K1��ك$��Lo8�\x�g��zŮ��݄%o-�N�֙�U��{̐�v���CA�z�1��p�������dQ��6\�*���\�[~�I���/Ǵ�SY�ո�ej���b��Eխ݉g$���ԣ$6�Z�6���r#�᪕ϒ�=�]�ނ<���%���Jٍj+�C�=P/27��6��dcl,$�ّ!��I^�Po~�j���? ��d��'�F�fi|'��̹�hxW���8��K���k.�jh6-��W<6͂L��Ѷ'����0h�~�C�[��(�_6c�u}B/�6K�\5�ۅV�*�B߆"�T��h>~t"��җC�|i���P[�]���̕؅��p����q �MF���Gx|*�U�,٪�Pm�w�4o�u���C��8;Hw��*@�g���«��ǅ�d2`Q��t)��V+���>�gxZ��p�:c:��-�H��Zmj>)��xL��ޛSA=��V��@[��eI���ag���"�sM�_��l(�D��ܢ!�з�3��ۡ��X��џ�*.��:}:������1���{j����G�)Ԃq�Ɯ��b��;��BF���[`V�^,���)����Ҍ��Y���RRg�7�:��^gc�Y<>�"x��8��d�}_C�`w䨶D�瓪]Y�5��7�H�o$B�!7���V��2���dP�x}(vX/���3S�A�*"]j#�.������Z�/�՘�p�����#�I& ��`�X�S�ҷS��t������#��V���ois~W�9����;[~� G~H����ԀF�j)dkԈW5G�A��#/Izn��&�O�U&����Q�+�4��2=8��@SCs]{�\�&_o�㭮����i��=�"�rǄ�3�7"M[��*}�@)�u�mkk*<�4I/Cw����n�gM; Z�#%f��ߺ7 ����J��}^Y%#~���a+>z�vB� �J�y�emj��I�WPrcj�g��A�I�fw/���hI1A�.�	ź�����ܨʾ���Ypօ$8N�N���X����^�^� 5�P_�:�@����6<���g_�"���U��mm�-���a�a�J��ڝD{ނ)M־��%����c��nJ��"K�|�Y ١-72�k��%����B��RD}3	m/�W��Ѽ���v5技�.g��8,���	�C�����#yS��w�oI�q4�lR �F�T� ��wިV�-ǜ����4���0�?�ϩ���	��閎~ >BQQ�c�d� {Eb�k�A�
<T��R>� �\N� �tu��ϥ���Em�)�@��fV�	���x�z����Z@��K>�7t0��2s�)^�
�O���?p��������/���[�vU[��S�'W�	Ryʏ�(`��G�h�g��$<9i�iTATU������."��l�,!�e�}$}��0ش!����RV�_��Bi��,�5�������z����nNH�!��J4���K�iNʹ�,W{;�c�|�P��/_�l�"�ЎK�^�2���c���sG��פ-H<`�H��d� ���0G!Cb�T�iHNu��N(�r�_B��m��7�"��1$�)�iU�(�=4{p�'���Q'J���_Qd1��4a��Z���GP��0����p�fh��ؚ�@Є,��M�>:h���"מ5{�R���m�n�K��h���U5~���//�Ϥx�|���h��B�>E�ׄa�7m=5ԛ�8Y�"*�n�v�!��rN�7u=3����N-}�Q$�THk3C�w9�ȸ��6��a)��r�w��٦�
��+��ևX�v�Wr���*�ח�`��)%���e�Rt۾A�[R�u�N��'u��R�:�-6`C�gj��P�7�8�<�e�S9�(��o��|K������Z�^�xW���`�K�(&l3��i�U��z���k�<�̞��{��Шom�V@���7/*�w��?�ѡ[�F=�n�#�5*D��!J{�$թ#<���͡�����Ϥ���r�F����xNiЧҐ:���K��@�����l�j����v36�r���QFFzC|<w��4RTS���4t9��I�l̎��*��3�Zե��r�^ �_r[���%�	�.E0f;�NPgP��Ё\ k�#Y�*�ٴ~xb�Ñ���i*�I���Cw�
M�CxbC�t���+�!����A�8̸ʭ�xqUșT�CO9n���bA���kl��Xҡ���@":X=�J��F>��f�z �	<w_E/�Gۚ}[�7I>*G��Xd�F�����6��̼A9�����o�G���/U�两��`4��Al{P��vF���T_�M���n��ن3�#2���hp*�6����j7G#^�D�T�j��ә�nʡWϫ�l332m�d! H��ݹ�7}_��Ƣ�*p���t�yIѳ�2�#W��{������?�Iv����A�͕)�a̬��m�Z���_lm��P^�IE��WG�z��:f�ɍ��:ƍ-
�s�d�����'lrd�7�T�̘߮J�����q��Y�,F��ح3,U�Ӂ߫���� �K�����H�;��Nu
gJF�L �8���w9��Z�r|]�Y�H?�S{O�|
�e���$�"�T+�?&�<=���7'z�6�'�'�`-=t�x���F%��I��MZ�K��m��@1%���Z�AB�TNT��ʂͩ����E-�v�uOe]4���V�.��������c�������|�f��rn���z�6އ�O��iD��`]��Rc&�-�O�AS����5���q+)rT���P��RjE�����&ܿËW���y��q'�دa|e6��Q�������M���o�Lf	���<H��:���i�� ��ݐ�� �59����;y:��E��@��2�TE}E���|�����΢��*w~�D������%�C �:*Sq̤z� r=&��Y3A=�(���%b.�b�I��	+\���su ��;^��ǖ��bH����Z�Q��`���	�,0{��+R4ً�?���4�cθ��x�{k�:�>P%�KQ>Z�Id�M2�S�������1���HLFCȿ���Da��N�>���밊��ˢ*|
ћ�G�"X�H���AՑ%^�����mW����c�z�
�L�4���3m_�m'r×(��l�*�7����F?���*�&i�sd��at�G��@aWa�R|N{d�V�t	�tQ#����},�-��y �'i���zen�ưg3ٞY��[�zK8��%YU,e�<�Y��z�-X��ĥ�A�S�� ͋�x=�B�#�������m7Z]@�k�G�_�G�T�{ni�x�8��0��[�| ��������P� �ځ[ڎu�ע�����=e֥q��fp4��9e	���_O4�z����!�6��Z
�S��@#���D�3�-�����Co23��(�c�P�~�3�����Ҧ��h��D�8==㾢�z3y�%��i�@�q�Rm(v5�WDW`ep)��n7�4ֺ���H�$-%^�+_"�ǥ|	�E�W�4�,-zW��� �պ�95�u+�4�#R�����M�/�ٱ VY�I���G�R�ME�غ$�`���N���$4��l��\3�tC�` �gh��E�p�����4����S�/�o�#��D[ׇ�J���>���j���J�5g�?M��h�00�v��T�t$9ٟ�(�s���O�v>q8���rEPM�$Imt�f7�('~tbj����C3�X2��茐�$z��Ojq{wE:��9w�^�56`2�hp�-�G�s"��=�~:��s}�w�4k�/@G����M�"|����[��ә-�ɹ�(sBH�Y��RL��,��c'��gd��^�H~v���9v:�L���d�c�����ޝ��<z�e�8h���_=0�i6Yt���bv`Kkg��%��<(Y�e��Jc�T�<�=�����N~[Ym4�{�}8���v���n�l�J���Wmlp
����Y@�&�b�b�:��r�$�A�!�Γ�EH��)ل��W������9���z���M�x��r9#�8G���U3/��[��g#ؔ�u�=p�U������N#��^�&�
5뗷�d �"��jHK������(0[[�EۧDb��Ix� �,�%�*�g��mA f��W�`]����<�ku�nW�N��� '��y��E��[�ҭ���Y��ܞ��B��	A�1ǓFh�{��~�!�M��\��͏���g�6a��G�˯�Z���u�'B�:ZY�(C2���];�籕��5^2�Jl&�co[�;��ڣL��Q8�\�\���XHNJ�Q ��젌�ѸWÍmAsg�j�ăҊ�;���*\���t�{�b/GZ����Ӥ[d��J�S���B(�[�v�	���Ukٟ�-�8E�t�]Ÿ7[Aw�=�E}�FKu�͂��1�����I�e�?,K���&�e��OT��\o��R�D\�6���.��]�Ѕl��Z�z�Zr88�b�	��k��{�YŶ"=R���|%|���,yK�	�<m�O{B�����zu���L�4K4xQ���+���!�+�XV:IC��[h"�����`��V�e,d���df8��*W�����͚p��=���xʆ�WWR#�x��T��ѱ��j�?�;Xݺ�k";�d����yBgݓZ��L���[�?E��KT�� �FS�eDL�c��$�_L=l�+L�p`�ٟ�{s;�;W-i�.�Kj��Ƶ���v&�|Y�_
�p�m VE�,|��f�9�e�W \3���T�N up��#a�K����M3�cU��?*xhό����K-vkJ�mW$`����z�;=�E�L�$�Ԕ����.���SI�@�����aO%�
>tj�`e�����\H+j�H�~	�յ`��6A���ЏK$�Nl�3�}��2���i9mĉ�<���d�|t�1hD���i�0�`W�2��$+g���
u�G����1$nx �?`Ӏ
_���Ko�9�)�{�@�$ ��+2��l�岡=�Ζ�,��z{� �YIB1����R�TZ��0Q�Т���1�z>�@�T_�L
oso>'4S_�a�f�H0w+�z��'EڛJ^�Pw�ǐ3a���5 0ߦ�`��ƜLf9%W W7�|OFW��ϫ���5�ȣ�(<��i w$�l�k��p�/�#F@�H�k��(�j��߂�rxU�ǿ�/���Ȱ�Mx�ޡꧾ����B.�[1�W�������V�Ui�" �B�^���~�#2�|+�,+H�44@��C�h�#�xg(gV�:|�N�"���8�+4���MJ����������Ot=����6V��ٝ[!��J9ҶZ'!Ƀ5`tQ�i{	ը{��f�IՊ���c,�h�z�^@�(�Znk[�0�����C0������Q�^i���� Ǆ�T9ԏ�o?�hИFY�	��|���xM��;SS�rT�nAwj�yÐ���8TTi�����M��c6�U�����$��"��%{EƝ��T��^s�=W_��?����ƹ�$���;rm͌���k�t���r�!^����҆���Y���3mef|���!��1p6�x�,��y��/urj-��fKw���0��>��R.���͐M�∃Z�v)�?��ӅE`�
�ԦxS����eB/:�$I�|���Fv�
 ��О�3��!J���B��"���1d)�Lv�<�v�\�VX��`m�Յl4��0���>n��X��n��ϋi�P����k �e��&8�(�8�>Ox�I�\}�:t�6��~JjŇt;N*��C7w�&3�G�=(��\>e��Zg���mA�#�Ç�ZTaMS�$����9�d��Ym��:�*�J �ėe� �k�@��@ �u�:��D� 򔕲��BK���V�6%�1��	�5΁!'C$������+��~��p��u���$����h1�^��\�%���1.W���R�?.\���6ߚO#!N.;�&X5`�G1*�)���ި�����+�\�9���q���V�*ă �2N`D����	�
Y���)�;��K]6Ͼ��X��l;�W�ѵ�/�
��G��Pm&vN��2�d�9�3�g���fW9�Fء�Z�ka�;�[�Ǻ��Ω.�m0}�*���e���:�E��'������г�Pxu�OI&����=�Cvl�;��R���vNCW�|[*Zj���4oe3]����U��@��y�	�T��l	�U��CJ���7�	�xY�e4��L5�7�]m�G����7����XȤ�\}4��N�qXr�V�PYW����k�_�y h�'>���w��Co['5cc����q	x�����D��>����J�8�V]�(jN�Z%z�W,P�ԧ�d3�d��m&���������6Qi���	����N�">���
&��]���&��(�No��SX.��frhXـ'5C����6w�U�
.2c��j »8j?�M��J�xJ��<�8�{�.���1�{���j(��;H�Lg3y�Ǌ{_cu����]��y.�)^���e	w�n�#��S������!�|Oa�uN�wI��Y�Ҋ����)H���ň��4d�-�>�-I���T���.�_3�Ǜ罫ÕrC6���;sjZU��:�����
�H���T��������j#���}BC�mfXu���vN�M�v6��>�u�����|�T,�}�����6������^aj�Sz,�G�TE�k�O|h�6����8��5e6�L��f!S�p0�k�X�[jF?�#}��qz���1�Dv�M��y�Ȣt��I:��_R�ܩ�o�R����Lt(�u>�UD!���A(���o�0#��4F0�2A���-�g�Z�cC����v����{ �e�ز���"�$�D�%]Ȳ�_X��s�'�k^9���5�->���^�g;Rq�F`_�E��Uv�g���&f���b��0�5���f�q���g`��{��b����a����Tr$i�5`������֮o����: K?�o�\�]Dz@d�M�Y ��Yd$��dQ�(\"��Q�mz�6�u��ؿ�k��E(#gE�����tk�/�!&<��)��'�v�^�$'��д����|n��v�>�O�z����@ؾ���f)���0��K�_"�kwc�D}���L"��4�l}��pW�WC[�|�B
���V(�A������o#XSǷ#he�h�b3�R���]�f��z�r�lO��!^��� v@�@�&Ay\\r�9G��I�mX�4 I�t��Qi��c�d��r{�7��{����}:�׎Ő7��ЪB�x�ds:��a�B����#��ւ�2�	4M��2���{|�|��nP-�b$x!�ႌa�~>s	��W��+N��Hw	�h�1'�Z�uL���N�I���g���ѠY��-xvk�tb����r�o��գZh��@h4܀��X7/��:VH��s�o*�#Z�B�7�jd=��6Z��w�@��&S7t�9�����)�$tj˜����GBq=栮7�N���o�B`ޝ��(���(7`���l��Y<�H֑��J�IT�N#��v��3z�n9Cv㰊���05Ͼ�mZP�_'kq����F�#q�o�\������X��M2E���JEb/�9V��Uh눇Jm������d�vY�^ha0��hk�B��'Xz�`��h� #w��E��kD�u����wAT�z]�� �KU,�f�q�ٴ�c�/�_Ӵ��7�0��j����W^ܓÌC���^�f�1
�Ur�\��SgC��P��f޴�w��oD �\x�;���:X�e���i�Z�:
-Ys��W�}'�Fa����wt��ww�YJ��q�o'v�78nT}s�Pw�\�DA�g&&��9iŁ��B#�a��_o��l���n�6�����Nbd��;�A�O��]�VB�K�����z��9)� ���\8yǜ�g���R����+�YB��0w�!NUfds,��P�!����P��)��t ���/�~䨧.��G{�[�n 	��( 2��@%�V/ߤ�G��o���䫐!�ҳd���ρ�>�c"��/	�^l�d�[�1S��wf=W]K&c� �7" �;�?ʩB��T�L%�NaOu����~�Z��=�����{�����{?v�|&�Y4!ȕD>�lx���][��(+%��w�����mf$>ƃ؈���<�ZY�٥o%O��_����YS_),l�{��ڠ���Cl/��!��)Y���G�~Ƭ�����5i�D����G�I�\��`��y���Ħ�
.��eK�:�%}H�T�m"{߰�l�v�G6��[�Bx*��݈�u�t�ߚo� R"����7/�(w��E�̅5���f�/��Dc�	~!�?[ ��ky���6�O5�&z(�n�q��J�/�8KMyaEh�Yn��~��P��������Q>F~P�ԕt�����.c��d�ӳ��J��mr�bJ�v����3�����q��C�јUW	���CW<��R^V�'C"��]��?�/zu%y?�p�?���]<��;v���_Q�:��H({u��Z�J��E�?�{k�a2�xD�ħF���?<�
�O-4�������෽&�Ёݲ�E
6���?ڲeK����^��@��o
{v�й﹵���>�!�Bb I�)4MA���ԉ�AN�=h~I' Ov��A�1��.�0,����z�q���;+ ���>��%/;ּ��i�O~�#E>5��&#ĽqP�'����#�2�d�#�ᙐ���*�ǕV��-�mU)y��a8�ŵ�s���."�]�����O0���� 8� �4T�����%�+�,���#˔1k���X�/�� �V�k�7`�h��0x/��J#=�d�["s�/�{�%��HH�˳�+�']��S�B�Z��>����C1۳�<Y]_?[QS�n E ?����_�8�A�V|Nm�[�0��?;
Plb��+����:�+S�TtȈ���9D[�esx|�W�;���E����`/�^3b�-B��jhG���s��P��Xm��S�3���W�S����A6�z$k�@�(t1�����wd�ȕ؉�t8��Eja�K���jXVq�^���Chk���D�����l��)�5%��@���j?+0��[��?u�g�SV���U&��ߦ`���,3�đ�ޔ�-{�ջ��.kv������2 KU�B�������X�4��@8��TC�����C��2�*紅��8��Q�	 ���7�S"��Ɋ���[���*ȥ����!2V
�~���2Ĥу�Z�Y��@�V�.4��H�� =�ա�f��}ե�np���`!�-�;8V� ��:	Z	�)R�ܿ�:K]�(���t�U9�D�[%����<b��R;�6�ڦ��>��k���ޥ;(���~���Ϯ;�rI����$\ 6Y��.�$����/Q���`QQc�����=� g�n���s\�^�KdK�4�Q�M��!�>�IQqJ��c�B,��а0�`���?/e��J��=�����c5J���"��#��$���k�bs�$��@��~�`�8<P�����Uܢ�❘w�XM�N�A�$0޳؀�(����G�O�� �ݲn�ə�Fy��Ӗ�U���R����C;�kk�����q0C3��;w�.�c4<�'5N�Ј<��4��q¦y|���a=yߛ$~���t�/�`�h�ȡ0�'c�N� �2UXA�K���S���RT�����o�3�!���S�h��+�/����If$����1[;���9��//tߕ�v�n;
|�dJ��"L$2p������9����Rb�x��uq��h�c��,&Q���q�x��W��.|���9m�;���uZ��/�=u������ܫ��~�v�'�J7�cQ���`��f{�ɩ���%��w��M��T?�	"&r���|6�g]����W�{�T��)���'�}�T�W�K�a�ܲ��I�^
�S�.��ãW:>r�o �����?�
m�X�`�<���b(���g$�i�����3�� ����W�n|�(�g�Z߬ �W������ɇp[kT�ػ���)��^)�J��s3o���i���:���B�`���y���T��r�M�zmt��0���B!jx�`��]��M	r���� ���i_������dy��l�cUZ���#�芇fwP��e��a#�*���z��3C�Y\ ��u��h�ū'Y�Q!-@Rr����!e��f���8���G�6�Ly��P5OJ5�!)���a�!	W�������8����r
V��ӓN0��U���V�%š���b�EY�M!�z� ���n�/ d4kf����%U��c!�Ɏ6����ΰ���c��e���#���`�t����c��g��1��A�٨�
2i� �-Za�ެ�l�p�?���d��Σ��_�gK�Dȓ(�H �(����^�����=�Я�}�݄��C�ɳL����'U�q��٢W��IL�q-��X֧ ���N��{Dd�vi��kّ��=f궁�/4z��6n���Ώ���V�SB'n<*�n�+�#^yJ.h@QjI���t�u���ܙ��y��kSF 4d����	�e��*�zW�o~�}\��\ި�����b�I��ޝ�:��Žs�mF˕Gޠ�Ƴ�Qeq�Q�<�<(�b�����=�����Ts�%W�S�#�����s���G����������t�$en/��o2Z�����%d�4)����	o7���*��Ыʰ���h�~b�,R�f�6Ϋ���d�O<��i��6��"]��ȓ!�>	�S4�s�)�J0CĮz�va�DÑ� G���Z;��x��D��3s�����­���L[E@h�+�%�P2��[����G��+ogE�2�;Dڪ�'���g�i��/j��v�X�>�/�4}���cN
�f�y�Oq�s^Ǻ ��z�"e�Wp�^���J]�h��������dQ�������'���yL\;�ɢ��J�݉y�a�!�Kq=$��}0�X�iANY]_���M���6�b1zS�r�Ѯ�����	\+'�qۈ"J-1�t	6� a7�}hk�;���^�� ��WZ����C���_�������_�B�&��o�sZ���G�Tԑ�(��@��!�s.�Z�ֆ�)�Zh,����e�vi'�Xf.���>��R4��F���<2���8>�FV�Jlh*������9���o���y� ��DY���T����� �;^H��h��9!�X�\�`�x���.�5��+X59�cr��n-2�1:�y��m�6�ʄ9�������aW�d���B��a��s���N#�лkrP��cޤ�6뻚e�\o�p�r�P�j\�g�:)F��V6fx��,��
���B�!���
�=��K6|,�©�V5�O� ��+��?8��|"��Ůظ���ә0~��l��g�y�dh���e|�&!�6��3V��*�$3�m�\����W�oo��1^��+��2��L8���U]�V�O\�H�md�I��U��5����v��@#M�F��@���-��ŉ�hrT�l,j}Qgӿ$���}�pْ�r����VH.e)?��a�0#���六���H�N������4�Ȯ���vJi_�u�&7��f�c �~<�YK(�O�H+lo�+|�Yk�/����C�w���L̏�{n��+)�,p�ي<�&����Z���L������h�<*N�sEA�0���M��Gs6H|���v>��o��P
��[�Jk��xՎ�2���f/a�����mؒ�I��ۤ�%�65�-�O'����d=��t�2��)qnN+�r�PZ���z^�ݒβM��X�ֿ�V�5}���E5�����W>И�#�d�b���z�y؅�7��7���w�U��lk�F�	B�l����)�����ց�YiB� {y�N�u��Mf�%ne��lܼ�?�gH90�A<�	�>�e�$����L����8�j��-�B ����T�WX�������Ng�0���u>M��ru�)�<��ߥ*�Dk��g��utމFhp���A�gB��d��I�FA�ɔ�Ј^���|4J��Ę�af�
&!i�@��;ۤf5�ijHʩ8����s��#�':
e���4�sW!�Ƚ���ˏ#� ����x����ꥣB5B��$�*�N{ɛ��g1^��ڋqk	FM	>JN��_�R�+_$��C���>���|�K���a�%�ϓp� �{f�����F�(a�u�M��*-�l�YmL�����᳃�[oXK���+Bv��UBT�}r����H?ɾ��b�7Թ�Ow��Y��s����Cp�=Ɨ���tI��V���P��	W�*w�֦�!��&�?��Z*��b竎Bad^\Um Y5D���<�i39�s��H�W����NiY�GݝR6&ݤK��jnY�;�����Vt�����V@ >!'6�]��ngg`N�����s�i��,V��4��&E����/�\��P�(��P��ݘ���G5�U4�ƕS���뿠p���KHn�ȫ$�Po?���1�@�L��=���� �D�F԰
a�� Ϳy���`���Zs�H�Y`��}��1YJ|P���&HJ�;�D���Ė�(U�Ĩ&�J�1R�n� �_��l;S�'L����Ύd����ߙ(���$��1�f�=����Q, ��z��kL��e�ֻp�	q��1�i�(�s���U4=K4gƛ ��Kk!۠�";�z�n֢�$�0�,'0̈́���, ���	fA�I��!Z���k�
�x"^��@��T�Q��=6,�����,���c ��� $!K����Q�Nmۛ�/u�Y�\IaK�����ԍ瘟���鉥t:�2I*��	[�O���݊e��y�hʡ�m7Ze����� �x�[��WN�F�4�Y�����rm��fj��\�&K��Y�2��W�G���<�}�YK�
�h�0�����]'X���'��ສ@�G�����CwNT%��~p�GI�ҙ}DQ��`�o��?pOb��Z�i�@��y	�[TL��dv&�5�%��������W�8�/]
��(y!H�K(m:G$�e27A39	`�M��>̀�;��(R�b�7�DFڛ_�<����K�O��;��\�K:3�cp��p@�o��Yu�T�\B���s��}s��A�ۯ��%�'��T�D6U�2���h���|�����V�@��6�V9�c�+­��t���e���>��5�R3�^�8q�[�j,m�|_�4K@�����%ݵ�mJ�U��N&_�
q����,�Y�%	� �}Z�	��[%�+��	0�������P��p��G�hY݉@RU�����z�'{�����C��hC�0�*UL��r=Z ��Q
��	q%�CP��F�"e�A�V�w�/�����T�ɉ���<���Uk�����p#��������?Y)^�<��^��:�GT���!�� ��Y7r̘of@������ ?���)�=�k�N�^a��Z$��k�G����D3�9�@�`�/ ��=��ݗ�T����R\1�r����o��v^�6
]&��G^���;k'UF�A��;��FQy� ���}n��������Y�62��~|ȇ�ꋟ;�3`��A[L�OT
���]����F�&�bM���C�D��3��i!�e����tl?u	������$i��[�`�Q���B��E�)2xj�ĥ�u�Y�k�8�����)��zۖ�v���?�؟���m��rHT$�`C�d�{\J�j��6�w^�NE���X���2��P��н��_^BWh~5�Fޗ�2�Qf��>0$�׶-޽w�@���kؚ�Q��5+=�����x�d$��d�ʄzNyT�Ƹ!�ta���m?ۦ��Ew7��Vm���M�&`H���
x��/���C|�J�|�=�K�d����h���ƍ��J��Ù?�Ι���i�'���|���q ���o\�N�M0���w�T$̶�i�����4��zʥ��&�x���T�R'��WL *Y+D<�/5V�6�%}����DJ���{Xmq��0�|�ͮS��dv��l�����t�$�㌆�y�����2�zj�{�̈�^_uU����9$�+��;у�g�KH��O	{��J+����d�&c�(�lRO��K�ק��*���{��߀>!Ч-�/].=��t�D�b�V<lro������ġu��n�o�D	}&*^�L�>���t�̟;�3�X�S�_��A�8���1�NƼER:�V�r��=@*x�ޡ:��:��ZxWJG!�aq,!��#�.q#��;mJ�v�ԸA!�4��ײr!sC�YHӪ�wU! ��,=�w�k:�<D5c����6 ���<�d����D�>�$��<Nɛ��5��OX(��8G��,�%��HT�Չh�SՀ-��cT4Nם�t7ˇ�������l�	]cY-c	to"��=��[?ٌV��xd�s�2�v�"�G��KU���p��;P���6I��Hg9;W��[������ĎvP��|���e���^��)몪WP2ax���Y5d���};�9�̇z����)~2 �S���Z�*i�4���N�UV�Rs����ͤH���R�eǮ����5��p)�7�Z\�ݭ�M���M1������R���r�E�;�.s����8	Ʃx�?��������^Z��6 �*�Fr�������j�+�|Nk���J9u6����ey$4�6 7p������ŗ���-f,�Qlz�{�Z��6�.���Vh�~��#~�s>?\̜�3�קƪǤ���������$p6l������Ѽ@�#	�Y5|cF����Yih��G\M��F�s�L8�̬t�lN�Z��l�|��L�?�Z���n�q��D�:�*�d�|p@���3��f����j2��ÑP 3	U-��dYS�X�U�:��%��sh��	|�v� �$$��k����M���$��_�lOq�}P٠
H[����	Ep0�(�r���{�W������M���L��X4�P�m�^qED��yM6���*�}�so|�r�7�h�'{˵E�o 	�i�	A�䨛�t��9Ҿ/�U��!��p��ad���@̖EYu(�F�PXO�۰Ӯ�����W�Iw�	�w:���X��A;|r���˒�oM�/E4�����Zy|���"o}2s��d1a�t%�_��0F�ҷ�*<C��f�|���!�d"n%<�ԭ�_��¿�l�7��FW�<#��j��IK.�F�� :��ㅂ��y콎��Z���lJ0g���~)Z�:�K�7
�0nq�e?�	|Za�Ȯ����Q7��~� _������6^訁���`+���z�x�����|�a���IS%���S��*�Y��\Î�ň*�nV*O�e�����ck[�u��� ����l�? :�G�E٣kY���-P;�D����� o�?�'S$��|��g�p�cP��a�gY*W��d���
$pH���bǐwMZfC�)5�<�ۤ��w����h13���k�;���`�~����^���/�f$}��	��:�UH^%n�f��5�)*ҙ��9ů���Vj_��Q�T�����e	�
���$ēL���E�Jo�*F��D�+�S	���-�#���~;޿q�bY��7{�p�.�^�h�g۠��J d�"%��fh�$92��_ҁt������Bz=�rbH�a!�Awh�U
"<1T�Wu�j�&��톞gA���#���n�':P��r�8?p��K�-�ݬ�tWG����7�Ώ�����CDڂǭ��A���_�uB��簍�'Ϻrq�{2I�2F>���p�;)�T�} ⌾���#���w ��r/��6yy�8� #�wYn�v`�[@I�8H�ܺ����o��N�j���Q;�-d���1���ڧ�?hsY �A�b�"�E�>8���@�G���f�p�C�bߣ�B|�rB����o����'~u�kX��c�	��X��;,φz˨A5���p��U�7"C�T���o�� l���$�~�
0�jZ�ge�1�u���XM?�P�a�t����u���h+p�<�Ҷ�`Q���4ve�a|����!�~.�?��� u�����6���@�x�e�P!)�?�\���;��]���~����АK���;q�[��bזH��p�������!l�m���cRp�|�!����m��ݪ��V|sj;�]�Q�ۮ�+զ�.ٹ�i�j�]�W�-@�e�,��m5>~ڍ��9#��� ���1KDl����%�ä��7���c�FS�#�#�ŀQ���1a��>%�N����/�Ɋ��Z��h>*��Q7��aN��1�3 �_�m̌�x'�� I����e��L/��>�
��3�p� ��`��b���6����C�xs
�Fr{��^���8,qoϦ&��4 �Y �O/]�ڐy�f�	 j�$zޜ�h��m�u�R"0���k j#hQ���P�� 6�NA���-��gj��Dx�*l۞S}�=��q����޷�LET���v�d��1�sF0���&?�Ţue��u?�?��*��M��ٓ��q��΍�J��^�^���Z�g��}?djM��<B������ş�#:U.��o�.p:#� �os�F���~��e=)c(�`���*Xv�/�<������h��O:����vb��%L��[�HLT'Ŋe��n��U�U3i�}I�Me�>�̋P] މܖ�DY�6wiֱ���Cn� ��4�x�+5XO�(�C����.�R�gc��n���F����lm��/���p��o�������;�����eP��{!��ݏE�$��ҿ�a8�T�:�+�Os룂���]r�K@�k�t�A����羪g�&�t��7Ť��e�"e>��\���L���)[	��r4���aN&�p�	YL%��1�+��=�rJ=W)93+����>�E��{ź��SkAPF�(�Y�d	�ai���G�^ҢFj�\��Z@�R7A8p���n'�D?Q;M��������_���[敖�a���_	��[b��By�S���g^��ϯIr� �f˾���Q���I$�e�M+AgX�~a+��m$�����C)L�_0��i��FD_]�bT� +u�W��P1ELy��|�����DT(���c0��@��3@8����9�hj��j��0��!����� �Hu)əM�N?,Hk'�F�MQ�G��Q��u�n-�#� n�.e���f����G�-{���S)���g���G��|Gi��3و��G�%i������b�Xl2�m2�+�*��]���}!0�%C��؁+��!E��F4���X����p�[�r�x�jsf�g���*e��d��0Eӑ��U�749����g3�	
��
�묛Xv��p�oE!����:����Ŧ6h�br4��q�-�K�Ab���ƟD�W�-"�	��A/����[�yLE_�cM�>�Zl����Qr�[-SX�2O��?���N`b?�I/���_�-�p ��s�MB���� �ץc[�Ț�qRa��&�U���2���6I�FEQ��:ҒyV.�=QO�n��[��bdo��Z��J��<�$�~=�~����D��nNi  _�a�r�w�
D���(��1����8n-�#m�|k'�O 0Zp���^��(���J�z����>�:vGo!�D�bw��:A�����P�c��,�2��ԨBÅ�>j��D:�|�}�[Tҵ>Q�6Z+�?�k� (�����W���[���"������=���:"���~�"�9ұ7��(��\�)%B�?�EJ�CQ�� ^8A,�1����E~4�8�_D(�x����AXH�N�r[$�/~\4A�zc%�������_��Z*5Z���\�v;��fMz?���~��u!�p��]\{ w �C�#~8=����ᒀyxx�別D�6��Cfz��UD5}�c�.��Z���>�=\�)8\�fZf`�^+@c^�U����+,_Ľ��'�b��k�|�m�Oj܍��Y@�g)��ڄ���SDE�:��S_]ݚ������^�4V��9��㼀�3�>[X:�<�f��ڂ, @���Z]WgΨ/��lų¶Ё�tq��h���Z����P������y2���G� �7�nz�l;S����A<��k� d�t��J"�}�����mW�V�#ӢW�m���_	tDY�+������J�����H��"�\�k���d�yt�Yuh#�Eb�,�
��5
�9y���> m�u�V!��^Z�WS�y�^�v�b���6�X�v��c��H����*�L^�>4{e��� ���b>�I�?TcNg�$��iy��m��`��?�=+PXx��.�����ޙR��C�G��>#�ޘH_gSԊ��#�o�;���R�Ϙ	�힀���B� ��@�I ��!��p
a������6!F�x�$Q�{{�7%��0�rcl*+!&�����u�L�~; &�<]��Jxw�}!��n���O�N�����U�!��Tt0g��x��~X�<#�]-娬��_^�2���bPU��}���lO�Fu�L���je��4_{�8��j9��Ԙ���$�.��}�Q���`��j�$5� F;Y ����+b�g}J�t��^h�2[ĠŎ8���rD^�:�%��S�b�M	9h�8�3��9�:$j�X�(
�_%6Q��"�Z�㙠:��"]�����7�(�1[��,�7��L:7�l��X��x��i��!�l�<돮�:�@�#����R����|�G���K㍛N������r"���*N�7_��<�# ��}LY���!r�>ƙ9�����߫�e�5�ZP�}hX_n�V���v�	�����%Ó�>��S�s�(���T}�jm�����)J]��r��Yy,����ov^��I��O�A;��AY�~���k���f�Y(/�0�{1�lE8>~+�c���(�D�ުV�c��m��[�sI뤜MT)J�
���wf}�X�q��U��7� _�,���.��`�غ�{Cq��$�W,>�d#Uj�	���#$��a|I��3k=���2r��Ƅ^5U:�eC "��
���b����,�6w�d���	n�.�̸t'��+$���K4Aal,��	�h�;��)�c��p�g�'n�2��3^�㔽�����lHg���vLh	�v%�ز+)�|m�ݣ�y���ZZG��oC��jj�X[��\M��[_p&� y����n�����qO�'��)a�!3��?`t5ޢԊ�yy>"��EkR&-�Md_�e��K� '\ۑ���k�ݒֿp�����bU��W}��+��>4��o�k��{�p�:�W�����z�`��Q(R�o���I�v*�O<_ �&줵��k�?�29[�L)(�q�0��<����l�eh{����������6�5���/M�x�H��񒙴n����D�:|Aɉ>b�����9�n��O�G`�.< Ҙ��-ha*���7����=8|�յ�u��h�i��DM,a-C��~���l�X�k,�����Jʤ�P�P�\U�y�UĆ�$VagvU��f|��������7 �"��X�U�n��V��y�[���g�j<��؏Ӆ,@�����^u�f�G6z��<���w#W���-��s�l�p�\2��uN�@���<�.u����$��1ג(^knE�Tw%�3�[��j ����=E��Ti��j(���X-�	�n���!2�_d����?kH�ȵ!r�n�X1ۑ�vPe5gt������!�>̇���&����z捹����/E}�i���#�]���p�)�L�ҙ�\}��Y�Z�c"v?��?
��r�1���oZ�r�����&6�'腵P�5��һV�hm�f�sYp�Y��e40��]C4��:��<ڷ�*���.ώWo3�M����s�� ��K��4�H�G#x��s�����U,���l��I�):<t�^���Q�x&,�̮�h�4�B([�X����B�Hm�L��Բ��~�NފR$��&��ٌ]��@�V~�X���ci���Qݼ"�ly\t٠ �Bs���C��C���އ�k�O����n��Y�mB�L��n��+���Êp���b�"T%��Nzl�[�\`I���ck����X����RA��K\����g���w�5+�+�	�ڮ���ϒ��
�$������K���?C�yD�ߔY�t�jG�l����-\�6�]��kJ� /~݌	XQ���P�<��a?'Np���_��xb�����IW�"��d�4'΂H��s;(��Qq˅T�س�s#1 ȯ�B,ҽ�K+ε���
|�V����-ȸN6R�e����o�fj��ܔ^���t�w�^�߹2�ҍ����|[�����"�������o\�g�^2rmI9Uْ��trj��J!Xg�
KG��rVj^ŗ�����#����gN��SJ�tk��w?��~xT��L�Ѝ��f�Y#\A����<Z��:��w5|�������h��-�R	D��HuR];��4�E?r�m�{��sh����-�R�&���$
`�_d�G��Hs[۽�� ��jZE(H[?�Wzv���ev��q=s���.!)��	3b ���\ $

��w�u��"2cl2�h����;ބ���p�"KwGp�~�<qh��� J��+,Fw�#������
�� �r�&KW`��͖���8XR�FC#���zΜ��*4����o
�|]��Z�ۤ�]��^�ʘ��S��U���(H}�n�� *�7U9��m�^��c]i�96��!�E�'��<78e;a���u��������<�׺�G�+���{�,6SD��B��)~D�_#�ZT��É_�n[�lt��sg����Z#^��k�.��HX9-P����v�+��L:��	]A��9�*'��1�������9ٯ�ײ�v�������$�A�h.*��_����J�5)���"`���G+,�j(�E��������֪����&K �>�QJ?�M^�Q�!
�W�2���R�4Q��I� F%\���4�hx佄�W�-`ف�7V�;��4 ����7��Y��(����;R-=X�y�L�S����үǹ��7ye�i?�p}�'A�M�?��b��G6���}R��}��<�\���Y�"�:[���a�l�c|�Q�G�h�yf���6�̓`��Q��#����| ��D\(>t�ڵ�~�����u@f/��C*ig!���t��c4�&�1zY�)���^Ii����j�lݥi�Gv��ܼ:��qKrZ`�p��/�*�r�W��r�� 3�I1"](pNf�E�7��nqn�5�B��(Kڟ��{1��Hҡ^>���C3,C.��7�ۖ�K;������if6?�h��{bS����׃��/n��^��x�0T"ƨqB ��0��<���zy��b W>�#�^����Gآi��b��9y���� ��%]a�b-��`�sL��|;OH�BM\a>�jJ�
L���i��b�91���vbt?,�F�:�Dt�����n�����eۃ��
|���ŵ&)�S��-�a�������]��.�%�3�tl��J�~WT�Q'����xң�@�5Ԑ��Ȳ��O�^�-
4�-�7M=�p�\�ԧ�O�%�ػ$+Rnvi�8B�_`�J������lM���ӂS���hmOb��(�`� Pg���Fv+h4�A���zk�X�W6�WT�����?�Ϩ��v�V
���}�Pֆ��\5���=;~�f�]l����{�2����3�a�}��Έj��H����E.k���-�������L�Z�э�8Zzs��Oߨ�y��ԋ���x�0m:v�c�O�z�ߨ\�����w�O{�C��}�>l���r^��H_ I5e�FHYO_�J��0\�8Θ�e4�A�ODU�[P|J��qs��4��Mf
H��.��~��-�I}NqU-%2)[��ek� �a�{�P*�}�q���ڔ�%�M�CW���#���HA�c��&�ɶ�t"��#���;49m3�[ vw/�PC�^�N� ���g�!k��R�z��)7��Ek����H]�N�z�&������x$��{e��As*�)���;'�R���w�b�l{J�KW��D��"���݅��|�w��kHA�d�I�:��qm�G����=���(����Ahnc�h��k+��R}2���x�f�6  �t�+����epV����?�{�� =��,t���c¥�⮜�K?��o*��i� �ذ�M���1���2# U�f�����蚂RU�E� R/I2�n?T,��������Ef�����҅��M�1�ih�p�~7������xw��nٹkú`���	OP�'k�uyfBFt3�T��3M�~u0i�:��W,=o�H�xs�ȭ�Wj^�[F��ܚ��ץ�7�I�R�j��lB�E�P1��GTV˰�(×���&{�w$Z�]8s����ђ�u4-��X�O�?�3	�	�i4�\����]�3f���� Q��uMN�y��16z���ܱVb
�=��g����;�D���W�n�6�o��8� ҙ��w[{�6i��0%�C^<J��'7B�X�E��k��A-�<�s:=�z�1y8�&)�$G8�|�dtH, Csc%�wS�9�%G ݷ5�{����ܺ�� t�Go�	�1t� �|S��1�r#[b0�Ryb���A��i��[M@i������Kv�Y-E:�X!hw��~~�����lˁ�!ӲrlC;���#�+.M$��Xί�/��VɅ� ?E2��h��	v�����bx�Ȕ_���C.�_�V��`Xa�Sqj�����T��v70<kΏh�����Ԣ?�i�hC�j=`n��\i�W�G��R3�꼚R���1A����Y*9�d$�W��ݐ����]�ɒ��-�9pn��j]��k��im�2&ó��mq+�F|�~� �,%�|��$�<%�p�4r��V�Gjoĭ��]mT�����K�tm`�}�Q�\���fX��;E��<�%9�(h��m@�7�	�!�c#��^ڷ0��xTieem�ڽ�}mVZ�'�RЃ��t��a(�������rs;�5\$�0�7��3vQ��#��ru�|"�UU��TS�I�3 �	
�нb�ַv�pm����^c�a$e�_��aJVx�B�j��-����' ���� +w߅�#7���*B*��Naʎ�A��I+ؽbi���4���L���1��*_�x�G�E�,�ہ�0����H�썡x�<"E�M�Y���w��%�������:9lsBQŻt��ͮs"l�R�o�.!ՈB�#�4'���:��ӟC�L��a!�
�.yNw�Å�;��홣�FR�At:|R���iڂ�uz����}�����AZa��B�갤�E�� �0D�θ4z|�:���>��q���T_l�&X�R;���N�!#���8�kx��O��i2�w��sY �&o���⭝�^Y�2K�K����:�v�O�YNh!�na��>�W�)LD�|����L2y�O9$xo�|�;K�&O��9l�|Kt�T6E����ys:��������¿	c��߫�CS���7ѽO��GZؒ�M�(ق���Q|�+���TԈt��o6�����N���1&��~	L����07�%�Tp�x�@�%"�b��� �A��g�PZ�����liS��j�-c�:�t�½���ދ!��W9�R���\�a��m��a�+2����]���.)#v�MwԬkM��6�����Ѝ��>w4�	����@��:�.�����%���zfT���r�q � {A�G�Y`�r=n~��~������\I��z UH�mb-���QI��/����E{�܌7b�J��Z��9KS~ԟ���V֔{�w��;w�TV2U�x�9X�U�Q��c,�!}ã�J�ݿc~/�{�!P�VU�����*ۡJ��$�uU�5v�lJB����=�k_��+�p�^FNڹ)�z[M?a?��u�������1rjz�ǲ��C9�j�cy�K�M�^4N�֞��8��Q��s�r���m-N<��x�l
[����6t��M��2���ǩ�V|W�U5h1�	
%mGX�V����E*�s'How?�w�s���O�T��(����P6_W���x�����ھ� ����N!�X��k�5$D�y0��m��>�KM'����V����\��޺z�Mǯ\"���=�Dpkũf�*j�\���ژ?7{�I�'��K<SC��&V��氥��b#,����1:�d�I�~�z*�*PZ�}�]cJHA�pC�0�@Y���y�	N�V�1�Q��Ýj��(�%�����6(42�00�]^#ܿ�<@�D�G��{3��Ej���z�0��� ܏$}��gu�pW�jW�;���5�X�Ipf���Er��Q�Ȉ��-8�67Q�ϣ&�b�u�F+;~��?l(:V*1|)!��:x2����b���`H� 4Ċ� �������?u>������Mj5���T뚌��c8R	?�"�� ���m�*GlwnT���r!rP`:Z���ŕعֳA� H�xN|��o��f��I�po΅)WC�C9u2Ы;�2�a��q� ��e��������T0|0�h�$��ӯ��h�*%��bB��.sj���W��@��	�	^;�68�ƪ�sZCũ$�M�H��k�q��{��Fi�6/ ���+��{��\bѫ\�	�8��-�瞩��0�p��U�]��R$�oL:�``��83�(��H�<Wv��Yc��N+d���B�D7[
;�9��K���EŵZC<�.	�~�ꂡ�mY
4;�����c���R�
��ѵ�Y2.�k��DڒO�0�2{�-ի��c�)��7���vGH��V�qL3e1ev�D�A��cb�s͆vE��%6
7a��vv��h#�*��j��tݺk����O�t;�����T��]:nu�h�"�q���-�q|�b�*�m{r�p����nf�����JB�Xoe�CxVM�s����"�e�Z�`P/�;	���]*J�P���|w�*�[�l�S��i��+ͥ�ap�T�AZ�qd�U]���G�v\ b"�ܻ�"��M���S**-���v��P��E�~1	W����͇Ǔ����P2zH���������N����KY ��o]��u�؍ݯK���fc(��c$�2+	�v�%�5��Je���1C�2��}S<+�}���>j�Uc0m���r�!���F|61�zY� 5\Qi������C�o�w�
Eb��H�sb����!�B硫D��N�R����:	�yh�= ���VQL�5޻�9V��J��dn2���3�\�ǵ+}����!M8�x��֜�8E�\�����I	�bo�n�kU8�ʄ��,|r� ��4ܮ�|e���Q�P1���^�A��,�xk�@e@�4Fu6Om��xi��a{f��Q����UG��+g�&��mKi�QӑVѮ�n QV}4;S��M`��_
+	�ĵ��li5�"��KFmkU��m0a��)4�}��I��? ��-\L-�X��vy���Cg�z�mMs���5�Y�Q��E�M�(����?���w����H�S�F3��
��O>����?D���Y��_�ڋF�&�Plp�p���f�;jJ�ԯ�B���� ?D�������iN���~���UA:=L��ҫ آ�%�	pn�Mo�l�"��yU=�_gn�����g� �O٣�O�W�N����a���8ʆ�`��Ií{����$2�ʠ�����dP9.����et�rN�������o��{/�@�X�����oR�s2�Rր��(vb�Z�+�^�ܮQ��, _��d똨9��s�0BQU����p(�ZC�RE``$I����t�|���z;U��z�v3n�GG/TUM@	"%�ڪ��J<qIMq[��-��;��W�tUy��]$�2�]R[��/"}�����r�ڎ���m꣰�T���.ܰ�a/��y���z�u��a�R�����Jx�"{c��e`g���O�HBa�v���U\����)G��K6 <���V�
�{���*�̕E�7A�s^?]#����<���E����[/�8�X#2��͗ؕ����O6M��j�����6͒��E
����Ǯ�/��A�'�Uʇ��F�Nn�]{�s1���IJ<��M����Ə��f��#"���Q�L�����K�{�t��[0��W����SN�k���O:�r�[tk�3<h�'ߌ!Lh9��EX��z�kԩ�O�L�q�����m�P��C�� �?����Ļ��wQ�&���$�H�.,�49�<�0��P�S D0����`^�R�	��(Ŷ<���u�Ckq���D5��΄{م�s��+�E��7ci8����9�j�v�Dm��pJ��?��a�#���{�Xo� X)�ܦC���}Z".}H��&T	�Qs�g�˥�Q�ohA���i|h�ћyB��N�<Br�ca���t��yT�L�4DaQf�������a1�a��&�U����CU}��1uF�ힷ�ǐK��:��z���jx����c����R�9��r�<�]A�#-pc�W�����*D�@ ����=1���wz��S��-��F%S�^(`��U����$AFH$y��������難����ҿG{t}�zeX�F��0p�]�N�b��=��?S��O�,D�;�y���H=��R�O;�O���*h���Wϯ��fJk�l��R�j'_<,�G?Eq-m�W+�h�1e�d�����8f����R���Ѐ��ܸ�Z��8�A�_������Đ-�ak�M��Oj �24�7��&� �=T�7I<V��-
�p�u��v���-T�GX��r���R�xBA@J<Vo�5���� �� ��{x���-◾ۀ��	�����ջ
%�=d	N��yU)�w4�B�]��K���CX-=��B��~���t\Z��)���S?l1|_�ujv�Kqղ>�/��8|�Q�wiG/���q�!�/Y�?K<��T�f�M����us�i��Qq9�&˩wo���g���l�����O$�G�\lb��P�h�7��V�H*�u�[W
�U�p/���,(~WY��]:qۆ�6��5J,�22�tsxʷ��G��.��e����BD����Ak�(I��}�^Aك./�������*k��&��:~@{�%�,�톇�,s�t�!;~�o�m�^������R��S�q{?��RnI�؀tE�<�ў�{���� �Q�H��h���E��'���9��'�6�X�IT���Jww����d@���z����X�U�8s����V�.�������v�����>Zs�]K �;�_1�>�w(i�2&��i�Al�/;2�R�Q+#C8#'�$���5&X;#?���d ,tC�Y�S�|���t%oQ.����� `�eXP���1*�[���-^�����L�`v�7,������)�rK�ߜ������E�=�"�(��S��l���T��V�|!����̮rt	�i�w��#1�lSⵉ,!��0V���j���B�ڒ�@�)l��Ns�+H�9P��iȼ�(煗y_�����F���![��"\�pv�$3{rB�t^$�R�}zX���AG8�#�A���Z^J�����dw�4q���������\ k�n���ߓg�Tx5�X�������t�ЙNڦ�,��I���a��K#s�J�;M�(HhG0k6��^���R������\��ƅ�1�/����=�x��f�U���ʵ�a��e�����d���1�6(��!D�ߙJ���*�4�L�Tǖ����w5b��X�{�g��=�{��&�]��o�I֭��o.��LH{JF�����d�NB�\&T^6���{����I ^yr�]9��`����Y�6�nBm��s�\(�����4��C��>}Ën�w�_���n|�0�Ch��I3�bP�$���˵H!0\?@�jW��f�g,��aɃ÷*�C-�r=�c�u*6��x��B�"Z��`,^A< ݘ���%T��U�'���f�������y��׼U�0Ty8!�.��#��l[��ݞ��Z{��Ϭ��u�7W����b$m��$���3.۸�(�($��t�q�h���w@���~��7ye��+��Ѱg˔�{�O�RCO� �ܞ���aA�P�����7Q\X])Ģ�UQ����k������~�Rb�&"Xt�U��I5$)�y����
y�<`k���ppmlrYl�'�AX_���]�̽I�E���ߖeJ���EB�]'�Þh�'�8-ï�@����nz|��R2��|:.�Ă ����
m�
ޤ`$,�ZS�x�����0�\��ASU�6
�A�fm �rȞ�2�����cp&�h�9�ރ��_СC𾫝���q��ሑ�$n��i��{U�6�H>C�ܸP[&�i����e<l�۱�/j��+��?x��w�|bG����7��s��@ի$��Y1��I��5�_���o���'�ܽk`!B>�i�����]�(���M�ȶi��5R�>D	�
��o|����#]G����%rj�c�ڗ�/?�{��w<��i���{�����H�W]��)��?1&�Pci7�\N�5\Q�h��YY�ҖO����wD7Z�ޤ��Co��\�fĸ��`�w1=�s�����Um��	�#�4H˓h-֕��M-,Ҥ�_i^Ų��{e.��2�d���@K���T|`��@n3�,�=��!7N�x�d2xRK�jM����(d5~��P�*h�R����z���)�1,�K%�*�V��R�s*��II�`�OOK�m� ��\�É$0��(��vX��J$y�J~��_ ��#Q�#Ў��d��`�]��vcQ-�|���=��3O���@o���R`��>ѫpq�o0���nf��y���]�r2����婏QzY�Ĵ�������<$9Z��&(؂�}�IN��`4�~������5K��U﭂����<TT]��A7�_S�y۠��9���]�7{͸�»W�rN8�ȝ~,YۧͲ�����v�t.��1@]B�q�3J̋���b��b�����ڵ�EN��"�e;_���:hѶգ@�������X�~����xX�Y{�	>��y%�2:��Y������5J��inoW�gQ���K߀|��O�Vv��]��{���4$��*�E:x�R�Usn�C}�2F>`Y�ت�2M�Y�X�`NKǻ7�tSLg��3��T�0`�Q�`��PO�g�J���R�����[��<I~09&Vb����sN1�|�W)�:A��=��f����=��1$���s�B{�k�����d���n�ew��oٶn�`��Φg���\j��i�n� ���wA���<4�]�7��=8ԭPIz.x��t'm��pB������ �W�*<�8�F�ߗB\�o�5:����9`����_�OL�\�Ywf�t·�F4�;7�a�!ʡ33����D\�
&,� s"d����)����X:_s�g�֪٧5�N�<%�����X��js6i�=8�C7�����5�AiB&����n�	�r�S
te���g�������[��gkJy�������7u��El�ɷ�_n‥����@D��/������ᑋ�j�R����3�{�u ,�E-a+����W��_��؋(vl�Q���Z�^��~��C��:af����i�d�U�Y4��^2����O}��wr�2��8��(͈���t*H��8��w2�L�0����/�~�Lt�醙��[N�$�1:7%���� U�l@@�>p�����D<re����-�ޕ�n)��b�I.��2m�Y��dkcZ̔,��ɢ�햴� ?g��`���d��o�E��G�f͈���yg�>�I�������'��	's��Q�4ʽ�vs��z�c���U�� e�l��j��$4����
��l�nf^������l|B�n��6�X�i�z��h���3���KRZ��C�B\�k��d[��Ə��I�H�7��Z�U�x�a}��\wT����i�5�?X��~B�ǩ��"�S��~ ?�~��i��l�>j-)���~,T�*I�6��&�����\Ҳ����ԓ}��M�y٢����E*tO�mIl�A�0�:\S����/�t�ñ��ը�����R��U�O����X�<7 ,Tמ�f:GE�֚�X�:<!�;;k �=4�_�yvTQ�A�F9�s�o�X���bC" .D�G@��ư�"��U�%���b�y��.�ZT�8p64J�$���<�&�GJI#�ʺ �u}��V9��tmC(�@c۷�Ī�����u|��m^t0�:�N-����t�����_ͳ�{5a�
(B]��ދ��C�ݔ��p�H\h_����л�f����� �&�Ckm��H�iu.
37���
f�kUF��$`7�ȀCg�T��FA�jS<�qŀ�g�*�׌X��;��Vs���9��U��!�ӄ
A'���(|�f�+���76ߝ(_���9X���:����D��Z��~$�,X˺�M����%��RAaOmf�k�3�x<b.����7�V�x4���v��	-���d�O�:5�C��|z~�1���=�Q�N(�[r��������~�{㫵��ӈn�g��f���WoH�|�R��蒌B�c�'w7X�]�]d��dh�I7H��j�_9:LN��J�'9霌p�Me5����P�K{�K��SJ���t���5���w�v�l�pV�bִ-��	�5�#R0]�4
�z�4��2
�xJ�_��]WpI���	��1�%7ȴ�
�&�?��'_�0��!9�
��7.^N�o"e�����؈������l�e�U����Wߪ[��Z�ƕ�W�p{��N���IЌlq���_��������yA����b��W�}�_�hS������ф�����E��Q��Pc�DJݢ���ׂ%f��	��@�5\,�(���$Xz��e؋o�x#��J�!��(�ۙuR<����J��M���	:"B�RvW-�$�z�(����_il��z��Hy��TrBgBm� [��[3(W���h:�E*H��d����s۬�oƕ��J�E�/��;��*��:s0��s����6��_�c�� ��z ��ːL�=/v��67���{G��*����0�<�p��XI)��R��R�2��q|f=��'�
�r1YKS�̪1|�E���_q����>�1E5ׄ�L���%���� �
F�qM�6saӢ��MN#�w����އ]p�C��sE�Tt��)��8�*��Y�)�q��<H=�>�2�k�U�&��Y|,�B\=���i�n8�k�Yҟp� �1UEip��'͕�u�� ��qY��V�hS)~rBeV���vd���ҝ����Y��L[-OE�o,�?��q�Xut's[�<���£SO���[�2M�JceL�+���+��$_b�������u*��������X~��$^����T�Wx۔�RK�f^�2PH���adǶ����M�
�:��� W�Z�Ȩي��l��eow)�P��R�m�� 6\ÌI�E�!X§	�.��W��]{��LMc�P�y*�'�U������g9""�
9���Lo�#��̓���7�j��p�=�_�4�@b��ˏ�5G-�#�u(��uT~�I��_S��9Q�OX ˞���G oW��;�{�q@n^���<���������s�7*0�<�'!A�1�r�|`��f�'(�����Ѿl�l՘~�Co�:�γ��t�3= }+Ͱ�!�ņ �LB4��>��F��#�2b��|�(c7K��,����`��U+R�Au,�jȇ���R�����]k(�w����ʍ�>Z���
)�!��PR9�eC#�/:_~�!>}F���2)��H�V~�G�}-4��U"���~sf�7�>%���a��"���,Úp-���S7.g�kxO�\r���I҆�������?"�@ah�^O���7��w!�M��|&7))�
�~1$0��iC_^���^��v�$�A>�mgk|r0JP1Qmx|<)��r�aD�;Ka��=����zD����YҎ#�
fc�9���!���S��:�kH>8�o<����?���h'<��\-|G��B�v���]ظ�_�^c3�<J'�"�7��KD&B�:��[�Cդ�wi4���������\B~X���9]v�Kb�O�$EZL#�{�����ٲ ��+5�O���]�i �]򮌰�����=c�;b���kp�r��Ş�&��9Ι������o9����,���֥�;�d��텬�ld�JҨ7jց=��&}}�c���y�M��/�B�o���Km�Gb��]O�b�i��2�̟�69������]�b:���,�o��bn8�g�u\�A�G�h�聸�a��j�ǖ�f��J��o�k�"�߅�ԘuG�=9��FKAB�o�JsLj��'�.{c���-���mC�HVE�=�%��⃼h���u	�_�^�WR�0B2	IvGo��
k��nM�:�h��*`)�]�)�7�Xo[CΈ	�ċ���Zl��vt��Ao팁R(���`�2 ��{����/,Z���p��u�x�Jz���8*��ᓀ�N�]H��iD���*s�y����匒�9�����$�=�Y���~=�7D��Kj�H�2~Z����v�Z^�#��Dq�_	�`u�ApG�����b1q�$���t��u��*q�U;OrD ����̻(���^@�~)��/c�s�eS�iS�H��g�m�v������_�y��6�
����+B�5�^;���<ʥ.��j�3\3X�r�DI���F�����e��XD�<�[K���[E�]��r-x��f3�?%�z�G}���q�i�Ǔ�j6�0��g2��U�M�
l��k���{@�}~~�F[z�5F�tOgC����(Cp�; �ށ��=mW]U�Ź�e���&ς��lU>�ё�*�:̹� �G��_���2(��K�fe�(�~c�}�~4K�����d��"��4)��&/C<��} �'DM�G��i1�o"���h���%sw5N�-�yUh<: ��?!��vD-�`;iEn}�1k��&`����Xp�]^�ص���.���o�P<Sy��n\��¼�i�9��q����0�Vĵ`3�d졟 ���t�A|'�^~����ְ���� �h�j���9�l*++9���+��َ�d(3�U���=��
��8�k^�j����p}�Z�4��bv��0���u���}B�<�k�SP$�*A��7�I]���-J �.M��n�v0���ޒ6��+��>��wVG�l����Gg\�,�o��%�ƪ��r��TȊ�k0��,z���^{|7�0�W����E�Q�[۞	�����t���4�dT>�Ę��	���V�Q/ ���0h?���rɎ�SmL������5A�EAH�컢�n�)S�.W*���%"�}�����S�١N�k��u��z�����[������Z��X6���5�]�(op �N<�k��H���V�=�w�G|}j(��$�%m��%�QY22�S9+*_�m�G�H���-+0��W���6�~Q�O�o֪������넾�O�7�2�gD.4�n9��A��)۶<�l5��5�+�7wڀ��~-95
\}ܾHʿ��E��]�g,=�`��b��i�}^����p[���A�"�h�x0���t����+0F hYlo��c��u��Yq,Ĳ��-�):�%�O\�Ns-��`ez)=�E�k�1�t�L��0�?UM�(U�#g�5����݄'�}���P�&��Y5'�0�s�./��y�X.J
H�[C
�շ��c��n�d��rë�!�Z/��3�}�vj����=��n�^�����W��E��F�9�+���Q���E!��Ɩ.��J\��6x�|�WD�ntm.�4����qw]!%�e�E}��m���n��G�i��s�ӂD`�O}
Pȿ�GVSEC~+$}Ԝc�<�o�/C?�RoY���%S!t2AV��a�Ra>Q�m����L���hRK�>��^si�����1�g_�A_[��O(i�����`ײjJ�d@����h�Z��-*�)�%!fN��I�\�3���Y�
��H�A��xI���ý��8C�4��<dC�)�гSF�Ѽ�`E��1�C�|�c�"��A���hs�g���E`�,L�^Ӹ]�sE����%y��r�Zk��_�9�ҿUZ̫���uA�����I:�q�`��[Sև(|�G�2����찺�'Vi�oT�3�h�|1��_��AG��xU�ao�!#�����Ts��H&�d֊h�#|Ă�/,���/޵f� z���#����Bf1�of�$�xc��"dn �-7��\�܆�&/8�}�#�� Hds ��:h�e�Z.��Z���;ũ}v*�3�b�y�D�
r�/��#������=�[`���ӯܮNy�񿴵ЎN����є�H�91\������\~ �tj1r�i��#��#И�l`a�����\��u!��0�
I��I2��k$��V��� .��r����M����K�-�`@.�7�YUm��ESs�k�����&^59���n���}��fF��]1��#�գ��BͿa(Xc�f/�v��}��Zi���J�n�a�=�����du"S
�$����2U3x�p97��<�(��:�l��g�#?3�=%����tw͚d�3��u��ѦZ[���I��&��
�N9��Ϭ��%���������jA_X7;�J(�!�r+�y�q7�S��RvJ�v��4�N:���bMu�S6M�{��%ww;S�^}�̀���`F��b;�QýM鬇h�#i����5z]��ݼY�Bh�M�w]���.�9��`��iח��WA�s0���4� �	�[4��E_���ڸ#I�{��i�<�����Y�P��q�z��d���76������}C����@��vZIa�ԥ5�%ҐgZ+��L�.	�G�'���,�m��k�)U?�j�l�g	e��9�T�Թ�F�syݒ�0Y hvB`��<�O�LX����$��L����JX�֑��z4���9��L�oI��WNyL�����'�����3���I5������b��H�%
-}a�~�n%�!*�eF�#т�����e, ����_�8ѭY�<��D턾���Ҧ�P_��h[eX�Ԁ��%�bƀ�Kjz^��q�|؞l��.��
Za[�����|{;�%nO�g�dL�+oDA)�j����{T�=i!�E�Wʱ�s�G���9m�D�^XpN�� چ��7gL2�۽�1�Y2	>sr;��&���٫�����{��ܮ�Y�٪���]z'؂Υ���^h3?YVV���`��8��TW�VMON-�ɉ��.�S�ξ��Hkh��;��i_�4�=�e�s �y=�X��(����}�Ե���X=�n���S6�]��W���lH8�Ѫ�ع�:z˻����[V.r��ޏ]�w8R��0�xe�����x�_|��-#b&���|JA�����֫��jZ١� ���$(l,[ΘE��5��ܬ��m��AR�3����>z�R�Q�Go� ��*J��&vi�X$;��B��O�X�S$�zv�������H�b��i.��*DZVN� ZS8|H;v�"�Q�1���hrFé����)Q�N�*��?fIb<�3�[��0E>:��.w��)\;?��߾�|��"��FfyZ{p��#zoo��*�:tXTw*�v�=���S�~h�c���|no)��R�?3�o�5r��ZZ+e�[J���Ҕ�ϛ~$��h�jy��(��#vש��=ɐd���ݖ|�Ѝ�pP�RRu�b�H�Sx�Ee	.�B3��6����,���N$�y!�ܝɟ�W���5'�U]m��)�u���Eh�R����D�[��Ƀ]���bC;�LL����Ա�̎��j"���S�/j�I%��~ke��H����X�0��k��Y��+�)N��Oɖ�o|fx
�&�ۅR��1�'�W�w!�k�mV�π�R^Ή�?�y���e��y�G�vN���*�]�	a�d>����*�5�H��J�O��!)���z��5�GqoJ��,�b�iJ��e]q�w��g����f�������t:"�FI��������%���<7� �Ni�%M�<�
�z��3m	�Iq'xX7�3��G�ң�9n�Ю�פ��������V�(��q&��*;F��2Kc�>���z�n�lN1�G.PeCM�Mb����EĮ��0�6^Qw���]r���_|}��ڹ�@=�'ω�))��X �e[�jcu~��?���{WJL�7����R�w������ߍ:]����I�A��:������0���e���pU�6Wꬸ�~FR�)A'M���e�M��G�A���>������xW�����]$[Amm����zj�4�g��w��H�y"j��ؽ�G{���6z�*���l��0��H������Ay=�@��eg$��	q�)��+iL�#�Lg���6�|��ѭ�`�B��9H:H�(��N����+>ϛSS5|�!C;j�[��<ˤ�5��#߮�zh	ȅ�ˆ���>0[% �وx���]��,E���X�R �c�(��	�X���7d}o�
c�Z+���]/��ʡ�Ź;����x�ܐW⌊��wM/�??�)XefZƓ����`n���r�;KoH�F������`_`e���"��[���<hay��j�~Ձ��6`�j	����̧g�Ĵ�$J�d�ܑ�,�eZ:�7.���Zk�yĒ�Q�γW(_.���[��M���)N(����)����8Jа2�H���˷�|s��D"�]3��s�<;��5��3.,s"�O����7�k?�6����h��hE�BPJZ;15�q���<����S2��G��͆a���;}�����s�=p����"Ŵ�tr��E6�W�Ң��w7��* h}�B��
�{�����5�~�h���z|S���9��y���~����:�~U��ް2V�=R.U�	 /�lZ�pm9�c
!l[�����<?oV���ƨ���0��"^֢\��\�eܱ�3�t�!wGQ�"���C��8B��^���y�XB@z0T��e4�Ù?��x؉'�8m�:]Id$�����5�aC���&��w@����Ps���]e�����iB��,,Pa*�[g6��L�_9=�=si�����^�E���ؗ�֐jܲtf�w8ۜ��t�x8 \.b#
]�|S^/�ѥI��e	�/���x�����>�	{����8��"�6� �H�-�������� �D�[ (��\+Q�O�N?��.���%�\,����hͬm����ҽ��9�n`�z���F�[���W��Qs���N쫒�g�hb��\Oj��n�P�y�᯦��!��� ���f�ڰ"eR3 ���@}��&��gD4���"&�k	.JM��$��7�%	l-h΄�w����Z�ٗ�Y��]���	~ u��w�v�%�h���Ufi`��"�#T���m�M����s�*�~>iBx,8/�v�Ȓl�E)G�b��*u \9;�3���i(�w��.r���/�"O���HT���ۄ�����uK��6������l~Dڭ5�����3f�1���'_ I�#���bX;Q�Sr�߃�W9��\
	~l�}���\ݰձ�8�0²�=܍�Kp��hV�!���;��!���ũ�Z%���;�[�rc�=�[��>Hn{ކx�X���G���?Ka��Z�Ϯ6���T�����>�"=�v�{�ltЪ��<�h��+\]�
�'�]{�[��_8��$mվ+ӫ��:[�P)����8s�MrM��R�B�2xm�.D?���w��[�r�"����b�b�&�*[��-|�f߸�����)?w,��鿒􊩪Cw��mt�3}�X���l~Z߂!Lo�@��Y�����6)����h 9���:��w��_�I��۳u-��)��R�ϗ���U����LS�a�8�����-(�/�@��n��A��ܰ-�e�؊@8��!>��mxU���a����8M0
Rx�5�V�
5�pW�*	DcK0�B��]3D��sǺc����E�yʵv�w5۲��{�����[������l�+$���61���.�F�c�뚆�5`���_�å��茴�|7�8��BFP��u�#����uX�1��T'��a=�!�.�	)��ĎO�F]�8�G8IQ�� uM��&�&�D��v����}�gʹW��{2B\�b[��Y﷝��྇UI ��X7((����I73��������{�y:v�sy��b���Ț1_�&	�C�l�g��K\�I�k�H��K�Ƞ�yWŋ$
`�e�$��Ri�%�K���Qxn����,��M?�x��L��+�Bg�}I^�DD�!k�1�K��񲄷 J)���[�X�?s�V�[}��4��vVY��j�~���.�P�OE"w2�����ӡ������������٤`��w
Ѽ_�"�^	^�PU�����`�Z/Xg�Dn3=�HR�0S�e��m�@�f��5;��	�b�i�(��e=�YF��U�]��*f�P�Ԁ�O�M��!�Nh�P�}ʊ��������ɠ�h��A�����5e���B[�j@Gͼ�F~�V�c�ДBܺ�����5�=�~0;�Hm�Gާ{�ج�}���)6�^ʾ�δ���VZ˽"����[=�׾t��(�PE:�%eHǳ��#܃�NC���WB�'-t���/[�ӧ�{/�K�����&��>F.�SB��z��n���J@�8�x�/�D�G*�Y-<�0T���v��U���)��E��u��4�� +1�HZ�x�\��'�4����g];���q���sK3�[�#	ƫ�,~BG,;�����G��4
t�4��VS�,�9�=�Rۯ�Erp����f��P��5���F�X��F�5uƎk�;��$������\���dK��A(J��A�~�4B����V�6s���V��1�+_�A`E& ���ۥ��M��'�ȡJ����@�n�P��=����lk����$�<q�0Jx�����l P+��G`�ؔ�l�hi��H6��2 S��*@���Y3L,���LUڈ;g�,JU��2=-��I�S���a��Y/$(��0�(e_�u�k}��Q:�?}�z����B��aR��rG��l��
ՅѯA�M$hЯ��2w�����[s�Tp|+V󊙨!�eE~`wk�w�xi�(x.�YSA�$]����z�렪���F��ũ2ŭK�4�'�+u%@C'�:�ʰ�/��;f�+qXP�d���6�2Usx�G�Sޤ�1w?~�r���a�Κ���u}�p�ؽ�~��{��_ň�g~�Ń���
j�0 >�ziJk8�m�{��mT6J3����jex���Id_�b��葧���#�m�ɋĬvϩ��#	���gǢN���D�E��y~I�j9y� ur6���T�E�6�W����%Y�k��z�)���5��U�e��Mޙ�蹠qOS�a-:�K۳�.s�ol�k��Y��:��3�$�N8go��Wj�=�P����v��?\�밿:r��𸗞��]��B�T��.X�:r:�ş5gj\F���Ƒ�~* ��Fn����0�1b��)��o��}�O�?�q/W���#�*�=���֮']/߬(�"����لB�v��t���]�BUd�������qU���z}P�	\ڔ�#	�˕��[Hϙ=X��+��Ar=�����+��iX�y��;"61&�����
��i\L\nJFl���(Ѯ��,��
�Ӊ��k��U����ѝ�p�0`e�`e��`���@2֟�Ь+�������z����q높T��L��B�S/eu �˽��	{�{OwY�߫D+�pw�3i�T�'2�18��\: �=�%l*J�k��*M!��u�y$�>����P\��J7b�I�%q�d�>���D�ݼٴI�!oqz�ަl�dM���w��RL��\RT��L,|Q'�f��@��3�8��aN�r䞕94^!8E ��^F'��GK�=���������z��6a�-���Τ��Z��D+����A���2�\�������[!���w>��`��V\2K�3_�J�#���z��TZ3�F?�m*��msl�V��w�I߀�k&�/`$I\4<|H�K��*{Vt$���:?T��5P�gЭ<��,�2�Wh�@�Rh��օ��F��]Bc�g�9�?�i;��~_~�f9��zH�g�;�e=k?�p93��g?��zi�q77rQ��r�a�(�F�Q��W�!����äM���o���;Ir�/_��F�dA����y��j��D�D'4*��W�lt伥G,F9�YKO /]�*��'H���?���>�J�G��:8��\kS�1Ĝgw���n�ɑ ^1j�M�g�4���xq���\��@�p��X�,���2Z<gd8/g�^[�;��ɬ����̦J��^` f�v|�cG5�!X"��6A\�KAx���TZ8��`$T�%.8�GIż��P�eUӨ[�'�nRP^;)�Qyci���p�ĉ�P0���㨷\3�|I(�ZGވ�{�Q��%d��`�{f�y�Gf�heTK�;^���ޠbs~J"�icO��d79 ������D��M��*�$Rx�(���E�%}a��D�?���u�q�|Ü��2�s�'T$�hw�f/�tz�����՜��;�%PFj�1}҃:ػ��%e�T��i�I�._+l�J9������8Z� ���[z)�c�h�`��;�@h�0P$��J�� 34�,���"�rZ*��J�<�L^T\���,&�d�E��4���#b�F�j����Һ�[��|�N�ՙ�&ȴgKp����X��q��z����P����"�&n9Z���1F-�6�ٯ=/���u�צ��<�p��ohT��n����^�ޚo�����`Fy���>|�k���,�u�� �M98.�G{�'u���£���<��U���x�ʿ Ųk��Ae(�:N��J�\��O����\��?���틔�Rs���>�������k�ăC��8��p�I�P��*� �@#2���C����K	M���_)�2��wU����
�E<5/U;ռ�G�G0f�0����rk�⅐�7Nn�U�\G�,��޲t�i��f]r]���|��e���9���=�X+w=~7�<�Iӓ��j��$��I�[���)6b�*�� �6^���4���0��3M�)�̌��U�eU�\e��������}dmuޡ����êi���H �'�y�" %���?��XO��HAi����jŰ�-c 6H�ӻ� _�6�3�v�l"f������<~�1G��}��t֡(���gPM�{xzE=8��QOX�\4�q L��ޙ�,2��H�3K��e�pf8řI�!�41����l׷��K�F��ǡ�S�]9����Qҝ}Yɗ�3y��������bP(�ҋ��>G'.7�?G�m�\;\;���V�J�j���]g���&s��6	�B�;�����k�]�ZV�����7W�F�dg�����N�9���u?	V���5� �f���k�H��t����	O������v uC�z�����?d��� S}y�8�J��b�i��	,�W1�5ϩ\��Ќ�P$�6�Y����stY��&4�]��33�ЄG��>6{��B�FeT_OeM}������?p��Qs9�]�Y0xݸ"�If�#��-k�F9v��^�3����L�O��
�Fۛ��ߝ��_-�4�%��rx�.�W����bv�Nۅ�r���!�8�k��EQ<D���3� ��hJ^���~��H�FT��+;��HE�4�� ��|��h��Q2�%SR_����N�.�P;L��M�7F�Iut�)��VVl���5�A6�ml'�6��|Ǘ\��QiB'���&m��t��H�����0�/i�����e	�lx��t�ܺ���n����A�v�q��Toi��2oe.Nb/nc[+`x� ��[c��d����q�5N�O
"�*u���gz�?lF��Wy�Aާ�o+��u�\l�Ś �cZcu%����qT��@1�uƐ�ϧ[�=�Og��*,�mLeN4˱�wl�`{'��_~���!��T��M�s���+�<��.��);�.��MPn.DJ�F�,X�)����k:�R���{&38�������*ۺ�Yi["[%����*��"v�4	�%��x��΂���n�)���`&��!7��\9�̹prT������)"�VJW}#;4W�g
��
c�Ń���\i8 6�^����-^kͩ+��ԟ#sBåW��ZA���@<jU�?���"���j{R
��t��~�����g�\;����գB���M\��TTQ1����̡��ƪ
���@�̡�>���Gwu����΄,������6�g|'۹�:�Q*�ρ���1U�(e��r�q������eo��>1�O�B&�H�kF��s�<K-���Lu譗^�����8I�2�����Ӻ���|.��z8�10��e$*�ސ ���1�kߤ�Si��0��\G�<`>u5W�2�۞�X�� ab2 6��dW]��#�!,���J�YqOqh�v&`�{)߽�Q�e��H=⺼������y�X��� (v�PQ���<�������e��A#|�BM�~�5�]�f����K�V.��v'8@�kV�D\S��9zo�{/m�/P�j�V~g���O�.�	�z��c�++
�Lڶ�P����%��j8��.OQ�_y�.�
nL@L�vQN\'��4�C#�n�.T�.�Z�ϱ�5����N9��-ܝ������7�̎͛������;/��<!�N�n�$op|��H�"�T�X����X�O�#�A�#��6.�R�p�f�'�oqC5�b.)8_u3Lmr��Q~lҦ���S���O�Xૺ[�_t�[-c{�MD���������)�k�����~���X�[	�u�+�p��2w$۫v7�R1�M�"Z����Z<������E��X���;��^0u������ m	�z��۬�{+5�2"B˵���z����Hr�qy�O��QU�YJY�Z�f�������{��(���a���8/�`�na~�{�6� ~B?�J���Ό��h�r�y���; ����4*���E�u/�4��h�A���X�ߤp���,�>MeŪC�AU�Ɠ��,.��
e�Y`Dg �=k�c��'A��h��Y� �t�*�*(�aIb�a�m�ނZ��X�<���K=���� 
�jF��Z5!��]�7�����G(� �uTlKa�2l�v���\媯�Po���_K�=��9��Qj�p{����m���h�`UO}Ą
�wj�`&t�_�������b2t��N( =9��Uĭ�S��s��+������b[䚸���/Osi�d�"�oH�l(D���F�㺟�e�L(��"�k�;#b�µ���%��CT6F���Z�$�n%#`U^�o�����mU}^H�v.i#p5���L�N!ac8�u��K�W/� m��Dhj�7��|��c��ȳS���uRj���2xb�Eb�4��b�--����׻���Hc^^+hS�;�ľ��8H�	�1XL�����LL�)��p�D��p@F�YJ�f^��ޥ[F+�&b� e�Fp�7�ED[��Bw�f��P��!2#���I�uh���e�	�C�� �����[)o<�F+��C��m�fS��Ju��C��-e��Go!�1\˃M��$�@��f��E�\A���Ŕ+7�ʍ����l!VY�椺N�[� 3�;����&#ͨOQ>Q��(�f���9_}b�(���P��?�L&�*�ǝ��7��7�!	�l�['�Y���	��׵�p`��ӫf2s���n��p@��<lp��0㨥�Й�I�دb���;���x/�d�jOX���ҝ�����UX��ZS�����]�y��w�����sG�$TM�쫸��/t𸢵ъ�u��ټ�V�c��0��E�90�6}�;_j͟�|��^,$6�	U"Q�E�Ɓ�7�b���Ά�5kP��Ê6Ț�[.��FT_x-�L���.���S2�y�7Y�-"������
� �	jGS�)������m"�� 4�}:S.p@2
JT#���-���yc:tޘV�q�xxxRڦ�Q��]Ʒ_M�A��(=1�P�N���j�ќ���e��`Nc�?�����(�}j���KD�aYY�	7���	�J�m%)Ώ+	�6D�D��!��qX�����,��m}Q�L�� ���݀�����^���m��<1��M
Oʪ�n���7g;�|�j��J	&�e���~��<Fq�wxo!f�KCuc^��}�EK����m�Bൗ�N)n����	�]��6�k�uTt/�G,��������XF�mk���
P1���8�rNʎ �-��9`�� 
d�[P���3a�,סmۜ�i� �̈������X[����{�]�O�����	]������x�u�M�O��m�^����\cE����)�sG�v��!����@��O���+�7$�r{I����� #WtV�	���k�#���5����ځ�uT���T��(���}$A�i��y��>W�:�Uo�&��9�O:z~)��(8^�z_����Q���omF��H�~}�	y�A|�z�;u�����C}�}�C�6׆7,�`��Ͷ�0� gZ	H慷ȥ_5-T4�RԔ7	7y�*�HĴ���Y;#C���SNʙm�����2��^O,m�]�;��g��g�����&<���2>�}�*�Vr:��x���x�`Y ���.�C�L�^U���B+3 �/�rKq1w1
g$�p�è+]��-bf��IBy@�X�\��9���(Ʉ`%%�; �hX ńAqU��"�ڋ�P��q���ڟ�f��݌e�����!I�����$	�3��[Jj��������%?[\�Y�c��$�*�h�]�^�H�����<;J�<��	�����?r�{=��0/w�W>�q	��3N��ݳ�4���
����my��]�9�Q2�Kj˳�`��P�" W��'���e�Y��d�M�Zp7j�^�S�i�F3�G�ISikخ�8��ǌr���~���죸,���gW�D��˺�4W�	n�>ד �+p#&A�2���v��1�w�$OC������M|�6��:9�G*@��'��M��|��v�wa6���{
��w,`\�  o.�9Q/s�zX'����sG�:�� �g�-MC_t��QӤGS�GBvk��'O���:fk�n�P�
ʐ�5�� Ev��}�Q������ l����0�(���AJ&T#R���H,��]`�;�}�0���Rh(�����h�:��S)�Xn5���dvz���J��������	��У^�%7�6)yϲ:���S(�g��'K��4T�^���3-���%ƳPD�����'�ǩj�W5L{�F��U.�DL�G�������:"����M�X��� s�ā�ċs�a&�<)X�� +[��S�g�a0� �$�O�������
{,q���H�P��H/:����.}3�+eA��g�3�J0o����-̊�$;�ڷ}���@y�����K׳��nyeQ�3���7d�RC�r�����wlÝ�oo���ԓa"�ɽ�J(�����Щ~�,Y")�OȂ�Պ%��%[��s�=N"ᾒ��o��&�K�!α�Q�jgA2�=�|g�N���P|�q:�w�r���#K�ؒ�����_���tQ��� f��DY<�'_�����xk*��g���>��W�.�[7���*�_+��q�$�-��/�m�^)0vUV˴�5l^5�]�%wr�Vs���x�X[�Q�w|M��(��&og��{��E��N��U����k 0�zr������|LCSL+���5���Y�>������͜��$� ��TksQ���Et�!Iž�c-����f�=��4(8(����,�j����U>�h�'�)MP0Z��'�iيÏ|U�26,#��p8@N�������ZA6���$��?��״@��x�e�H�/��I~sG�~�8�F_�����g.�^l6*,V��S��L�P�)Ě�Y��1ںCH��eAf%�{I�Iq��	0R(ظT����K����	�cڠ)'�Ƹ��%)��$����lׯ�z6���l.-��P�� �/��4r�(�X�����y�G��%���F���]�l\S�%�	��z��)E��F���j���Y�	&ӪK�]��N���Z�'o9�T$i�fz�%�(=���|�[��g�R��p�H~~��Ac����Uxw\��0�vT��z��=�n��&���1��7M����������ph�n���t-��o,]·+��k;�;I����E��kSU��EoA֗�D@�[���YϬ���І��6�+�	n>.���c��bz�f4=�8��v��41*���]�cXJ�):V)���V�Ʉvw|�)�nb�s��������_5H�K~�>F�)?�(b�����[�� O6{HO��Fb}���^��S4���	����iq�C�!� ��J`�#����" ��d�kRh�P�(��w���tO��.��݉:�hLK�	��6�CՇ8_�nKC��R9p
!-�9�	r���	_x�ωy?ص��|�1m7"o�3�Er��']`.�bڃ>����$��EL0��0tCţ�Ҁ`�O�p��Rh�&�V��c��u���.=t�]�U�v���O�^ ǔ��Nњ��%�@\�pд�4��̌=����]�{m�	���GE�SgHf |���}��˿5'�����N�W�h�C �
V�ks��9B�,�	L���m8�0��mE���~W)�X��i-� ����_:����j�
Y�=B���*]!��`N�A�����<R8%��ڵm@�4u}֘�n�.Z���pO�m�l�]�����(W�F\7��j��]�V^P���sC��h��pR��hЭ
V��~'}�/�y߻/|��g	w�_�POWX��r$8�y���Rs�>�LQu6����p�����+��.T�z�-W���'sb�ݔ�1Z�W�s]B����~'n2I�q���H�X�u@�eH��^���w�0��w�����g��r���ӫ�R���EC۞�6��j��F������F��Er4�x�>�e�3n��k?�Ly9w�~����Q �~��-)1�$e��|�r�e�|�+~�j,�:�!�{�U*o}�k�qyi��=�-�\q�TY1G��Yk��1|J�o]y|���i�Z9�ȉZt��9#w��;z'�ʘ��p# � ����}D"p�\���a��j^sB���q�U�Ӫ�����J�6��.O����%C�Q~�%uD�"�6�7&�$��/��y�&~7b)�V���:˫�s�=�I�e�t��8R���J�3 AQPq���6G��ȼ�͋���~�r���馪0�M��詡�v��I�Ȼ���@���s��Y�����(�U�G(m/���9�P��o��u�'��4' }�~�e(g<J�^�C&�&���a��^.�u���L�a�T��a!�g�}9�9 z�Z[��W+��p|��l~(-i%Io���:����A�=3 �%<֩fu���=�r����_P���1FClv��9��x��|��U� �;;������g�fa�T@�h��1!`)d�f�P~-B�Qj�F��frb�!�gF�wj9a��$z���Cm�E��d�!�'����b��=ˍy����^`0������=�p:�M�G����)��lNѺL`������]����0 �a�N�x�#I��-��ƾhF1Bm�ov�)�=��V���U�����X?���B���Za��rh�	"q��Kn��!�}/a�ֈ�ḥ<PbF�6�j�r��n�ƛ�;XRZ�֯�2����63� u��τ�%jvc �¶��__�S�B�j�w>)��lM#��#pHQ�Py�a ]���;ՈPt���C.�W��T�W' {��;�[$����DA]� ��M�vb�R��b���)�#a0�������(����3-Va��H�4;U'�A`%R���0��%�<�~���y,��<��7	8@W{���l{�i�j3Vܺ�
G����3_78�̳�ڀ���ǈ���VM�
>�J�J�<�`��|�tv��6�>�.�d�����ĥ�
Ѳ��+7Z�H6���m�D]����d���U(m�<xk�SS�`����0A�����x��>K�����\A�_�)3G��t9{=��t�d�H�ǂ�eE/4��E���3�� #Eq^M����gD1��bbG�9�C�6����:z���z��+����1e���(�=w��])�|Gf�AJ�+�W8�R�5��Y�l��GH�wOK}�M��n���Mh��]kל���;��!��Ȕ��3}H�+\=11.ݹ8�M����HX/�K ���)��sN��wD���Y��g�O/� ,}&n0͒��[;}!X��B@6���+�(��A��&x�c��9j��Yj�[.0�{�f�.Q(~�h��)�	�����}�A`�!����KFn�4IM�� ����5zp�B���w�����4�b��!/ �b�Q�J�\j��Tv�D�UwN$�z<���b5t��)f���t��@U ,N4/ѠpzH��x����ʁ8"����tSA(	�l���B�,�ٝ���$�ś �%�!�f�y�V�E2͕^�	Rʲ��&E�Z����~܊]P�A����l��;�������rQ��`h,�pp�\L� U��2��i�m����������Z���P
6�q�A�����1�pG�I���������q9w�3F�!�S��[H��)�R�v^>4��k_�+@�S7����
�XH����.�=��r3�[�\D�N���L�'!����&ݨ����'�\�i��>�Cn������+sP��u�a�Q��2"7���
5������z�	5D@X�Ab��}:ڥFC�Q:��y�g�o$!3;M�o��v�`���)	�����|3h�ÈS"�SӺ
!�eX��
9X��G�u
�}��Gy�N���9Pk�@�T&PvOX�b;�?A�.�[�TK_� V��Lʟ|'(G\h�w#7Τ[%/�>r���+O��|�C��t�A�ݬ�u���Z��� `��I��T���iM����W���P���y�(�n��d�����Q�@(���Ў`7�%(~|h��2!J~����y�����ru���#�b�fq�\)V�$�^����di���N�a'EP�6�e�-*;�TEQ���7|TJX�J��H;upʼS#��~�S�s��(rJ_�g�Q)�؈OB����l�w�^�M�m�N��� �n�↖HlC��|�д��͚_쪙0�&��Dj��.��R���S��B��7\�}+�Q�RL�'�������*W���V,���{(y�>g��#G"?ӵu�gt�K`��rd<��G7Pw؏GT����S�����KI.W�|:.�k��1�k�!��վ&qsS@�x��>ÉEk��P,� ��N��� ��@�U��>~:pʪĘ��}Pӛ/p�{��WV���C|�K��)6W��d�-�*ؑ��4���y�P6�2r�"�0w@Jz&��N]{ԭ�f�/�/�MS��z�q�P�ot�2}ΏF^!��dA�u�������vat?����\k{����4Z�$!{�y�*f��i�����
�f�g������ i���*W���ja;$�0�����^���8�jHY�#a�5�� m�Z-y�RF'	m�m5~�D��z��wg����^��?_R&�/��d훵�-v�%
���#�f7;�g��p���C���T� �w��?ljq�?�W=��H�w�7Jk�>]� w��������gk�6�s�E^���]��s�[����m-�֒���M�1K��Z{>$�f�m/�Ƒ��{���g���Fr����P�5�.5�"�[���3��n�g�j	.!n������E���,TV$ܐ�B�a�~-�H����Kĺ@��L�� 	@a�w��Ki�����u��H��s+��~�D)ӼO"Q��%���oo�y������{�8���
;��9r]$7��N�x��5�5�}l9_c0=3��dz�<�UA�wh�d٪���z�Bse�O�H���Յ��d"�q'���\��r����が�����P�22�m/]P{1���x�������Ė�#��<Nk�5�UuK��m�𣯦 ��,��CqKJ0�> �y)E��a����}�E��+�6n�ay[u������O�ۈH;�e��	n4ӥ��[��?������i��ĵj��Q%^e*��U�������A"��vg)��9�`���e?�JR�[�eB�u�x�S�N��#H|O�sm?��>�<?��V�ɳ����hư�i��U~��uU(���e���\x�I迖ߒ,��9d�늣7��5ل�.y�͎ۥZw�&�VQy�s�m� W �*f4;�)����av��`�X�r�{�$vخ�>�'�mX�..���9�}3FҘ{��,H8 c��K~��>%cK�����R��ܾRN�}��� {�Y)ok�h�aX/ڽ��cϜ�BI}��T�*�V�.�'�➻�F��JmF �Y���o_�\�m&��X5�.DG��Ҽ��u�0�ۀ���A�8]�g��Q�s�覿�SKBմ�����;W������4M�|���l�Bf�%��ǐ��)���R!�m�9Uf�Dn\�:���Q܃~��T��W��^������Ò�	�����a\ӎ�ւj����7V���0nR���c�9�-��F`���x��[�e9����a�/9R{��|պ�l�vA>|������m�Q�d����=rJ����+���;�A��W��&X�4FR���F����_��UtF6
=ggK�\����I�FG�x��gܚ�����a˂|��v��7ɿ��$2\R���)w��j��t'1N�D͌�{|�ўJ����VX�T�áݻ5H�:��^kSn5%���m����@K E�����`�ۮ_�\Z~%;{���B�\�:�	Ȫӥ@�Q}qPӅRLJӴ�K���-�>�-����3��� �E̦�HA��7l9_���cZ�w+3:�2����@"���x��y��>6�"K��!�Q��|y/�p���i�qP{]A���X�F�d�A��a���M ���� ���������LH���	�aT�'o�|��ϧ���a=�`v2$TH�:z�Z���N<��@��E�f���A^%�ʱnG�^ Q�ɊH�Y�"
Y:����PEz#q#32O��̉%�9�!���֠�g�ϳ(b��4K�"�$��ӊ&���s9L�y��{e�|8�#�K<7�:o�Ì��|��r��+x�\l�b�]k���Yս3w���5�D��~�+JT�B./ �D<��U�F�9S�T�)4�����P��eҞ9C�l�ߎ��*�\��7�d6s�kRV�
��Pd�����;]R�#A�Hs�d�C����*��i��.?v#��p���O�a*�����\�/�IM�H��u%T��@�}��h�� ��:�/y�|&;�ie���3?O|w��@|����M�S������=�"�\
��m��)4��Y���Pҟ�ҋ�����XRe���}�°��5�#Y�X���z��iW�v��$7�`�X�.�4��Ξ�~����z̍��n`��9�k^�όޏ�'G�&q��lݛvGRVLa�O��n�ZA`/x�~�;��b����h�4%Q���rٞ�\9�H��ʎqK����?NlB������{Ͳ�S�+3k�)�?G���s�|���,=�^����RZ��'n�܄s6d᾽ȅ�~~|˟������?�M�iK��U)�b���7<��녌\��#_r���O܂ꗱ�[+�K��d�{:�B*���G���q�Te_���������9U�:�izez)E[��y��A��]��p���HU'���D]�����ɎX��N����e���Ḓ���{��S�呠&�5�p��r�NjG���� ��3������l�_����CEGr������$�>B�̙��U'���E�ɏ�&�3�I�qn9A?:>Dmc�)��l=�l��6�+H1d�(g�='JO��pW�nъ�P\�Kk��A-�	B��( E���'p�yo��Rs80r4�=����C����p,>l"s�xJ��ޓ$��=rbO��-f��-O�Z�Jz�;U���,�@�`t"�2[�-�.}6�O� ���+^[�4F�XIm���\?��/w����l8�����L�������4�����7=���W����7��zN�zy@�ݛ,�)V%Ÿb��X���i5����T�drN��h�������<b�*xa�U�9��/\��p_�[ EY�	��v��5�e��CW��%�՜o���O��(���s��g6ȹ�y�/�7��r���>�QshZ�b���l?MXH]+_;m4<���.X�"��n���ڹ�5W�Ƴ��A�5��]B'�z$\�X�e�$�n�<�UeĂ��Z����TZ�.H;J�A�g����l�(�wtf讚_M͆I��	��4V�>�i>�TYC��4�xNH��ڡ/�x3a���_/��8"����$�mF�W��{D��|d����&c^G�x�N
^E�z���^����O_���VQ9>.�9Z�{S5j��*�i�jg�8:Vh^tу��v������ՠ1���ϑ��1��,B?*�f.�uzq�Z��#�P-�fm�/։��o6 j �5 ��E��f�?���L��|����m����}@w'���B�t���d�Hu,�w�:��%����I��2pmQ�P�<�_��b[���a.�/s���}���,f���P�Pc���s��kw��f�͵��[��Ծ�sS"��P�_���m�۬1q��N�1���q��J�,��2ρ�� U����|46�PK�c?KR����|J��}��()�,��&)<��s1m�g1|�Z�F�Iݢt4 �r���?d�#���w��k�<�LDC Ajes�M�l����Y�O�w����ph�	1�U�=P�ݭE(��fnJ$�y��$ 4�Uu!�{�$֭���l/W@��Ҏ��Ff�.7��9�?nm�NK-������-%l���ڭ��K�я��1�B�X���%�W�g��D`$��F	?�;fk���m������&�ۺ�6^��rR!�֤zq��s�� ��(��E.l�F4�T�{I(���n@u�(!�^o��i�q?��E�*3T��Wq
q��,�_�87������X�е@��k>�	����2�T�
MWG�?�E*�Ic��-��(9�Q�}&wy+�/��#����N�u��~x^�9�x�=p\6�(�ς T�'�Z�Xʙ�qhB ���G�<�l��[��G����ڗ�����y�6�Ө���I3�����	�D
f����W�dƱ�j���f=�)7I�*5t>Vlc�6B�F��&��s�7�7sB������S"'29=
֯	�r����{�(o�X��*=�3\m��ȗ�8��w�`�r^��J�7�Xw���y�H�H� ��n�8$�i�����E2�R4�V�e�a��='��B�(=h��ol�)�ZWM��޴6۰(�"yUR|Q���}X#�ϼ�lx���o����?�o�v���Pc����zm�e��X�j-��`�W8��Z=T���X�-ISi�W���,����9��>���~@%�R&��/@��,4��j>;�GlZd9H�3�]}��%�.��J����1$���ܿ�#�E~d�C�cD��Q�UB��9ߩQEk`��e���$*U0HEGtcCHV�,�����O��tO�b���\섉}T�P�ގ��Z�W���ٽ0�B�X��}�D�u�i�n����=�a�����n��Q�ɽ�fJ�:>1��K��?�2o�g����kD�)ˣX����;�����t\��B��m�R���ڏ��{E ��d��5�JCڔ5^%���D�]� �8_������G��OD��'M&^28�m
̟��]S�zZIp������?�*�V!��L�T�AA���:��!e�����?�D�C��ŕ��/��M����j^�T�����{s�J�e8��G�}+t�:�jWx�|�T>�	�P0��D��|~
}B\�q��ɨ(h����S^#[�W�DXZ}��D��Z�S�S$��"�����ei�y���V�sg�w��2�%�h��JY
�f��B����9�Q"��d �|x�hJф�cit�qHS��շui.p��
g!���+}P�����tS�a��*��F3gd��c^<0��� Q�)j&{$�A�X�4M��=]�`hy���Ƈ� yMg�uG|����l��N�w�]cP������bz�q�ޟ-�Q�yx\���(d}��WU�2�}o �bn����ۂ�����N7zO�yP�졅��K�6����y��Wۊ!?�{
۬���|
Ĵ}�/���;ϐ��a�w8{[`��zׄD}�EJ�.u-�ކZ5A��Z�=�ܙD�I�����t�~9����]�:t�c���kW6e���$_3.L��B�%���.�(��k�G=��y6D�����[Ւ����G)g�	�����1x]}�������W<�m|��#�=Y��-~1>ǢK��v��G���m�aZ�\���s!	�k������u��K���mPr���O�J*�п.+����ҡZ�,���n'��(���i��t��27X��o���ĩ�ٵ&����X�c�ԇ�(�=m�ߏXU?a��
�[���
 ��D���ʪ}0�4@��T���]���2��+Ȯ����M��Dx@q�?X���ּ��E9~#� E �㫠1$�OA�~�h�!�Vݚ`�Q.�kbsK1{6�sR��P�⚆�og!��i��c��IBL0�}����ݤ�6��
YW���C޺𸼳��,Ө�(�?�8�����^]P]u���i���L\)Tt�B�;Cp�eJ0�#����:Z�B�:(�?��������@@vmr휴�O;A���x0�]���������+�*�h!&cl� ��=�ũ�C�;[�:y�W[�/� J��Mt�j:kc>2N��O��(�P\�ch�u�ナi�Â[8�v��2��=>zwP%����q�~�$ƾ��v֋��R��xFG� 5^Ĕ!'��{�r��jF:���5�SlA=Z�uɬ<x��P��v��l��==� $�I�3��
��[��z�����_6��� e��_�1�##��L��HsTҩϢ�'c��KgT���������$�b��QTr�H[>�N/�DR���+p�0��:��}�Q�\+����v���u�B������J� ����5ZM�i�)�4��O���r�_�WAXh�BtiH�2뮮���Q� ���s� �!�G�9�i����KԢ�ML�&���������0��uϸUͼ�n�0�:�7�nL��<`ލf8OC�5[d��R%��#�\�А7�K'bfy��g�pâ= ��`e�mk:|����@��g<�N�WILy��t즾#뵌�U��uxZ�s�jv�N�8��\�1k�
%z1�DC��r���#��Q+U�|�TG���p�[Ν����&�q�ID!vʋ�T	�̛����@�ÿr�_aa�Z/��F��g��3%L�j`S���5R����1�\J+�!�H���7�\ DK5-�Cπ3�.��o�:���y$~Sw�����Ȕ��y����6ܠg�s�q����K�Gc}�� �0T{|``�3w2T������C�+M%�\8+A�E��"4�vX����W�kc�z�S��S�&�-���v#�RUv3�R3'ˏ�8e։b	�2+�ӕ��@��RW�0Q,�Uc��!uG�M��ђc��_@ltb(>0�ﲘ ��it���#@�]�'�G�����TQ�*t�"�W=��} ,R-5]�l<�P��SVt�ޓ���4�fGx[�M�|k2�w�i���8� �\:;����D^OI�e�!M�վ�@��k�Ay�Ú|���/�g�Q~li�aɞ�JR̳L�>��t����=ۣ�f��N�Dr�q�7���"G�J[�Nϡ�:�(�O��l��v�a�����Io�/H�	;���
�䆷���(�g�2S~���rF�7 ��Î�q���"ha%h�^$��SY�:ĜU��~���l�\�)���x,���n7�:�6�J�7�6jw��r�5�`�'�uT��U"ꅹ�7]���)7������5����OR�w�7)~|\CPI��j~�e�MS�ɴ��<$���8��E��fg�m��f�x�X��m�gWY�X�a.T����@��N7��1}_H�ť���b�wR�m��R�Ȅ	*M��:�Xq�h�d���LbX��� 0O8R9����.'*nL���z�]9�DB��Ǔ���PR?G���4�Ŝт YV��O{ѧ���:A%���_�C�[�)���U�y����3�x�{1��[{O�Ό3��m�r��X&����)`�I-���\�ц�,��mo���!�@ڵT'��!��=Q}��jD��tT��\���h`��P�I@^e;���	�kKO���Br�F�w�T>T�Wj� p`n�4o[�m%�7y�Ě���4����U H1��ӌH��[S�igA�W�p�2��2�=�#H ����Bq�i�?*�/Q<�<Δ8����~(�Y����`C���V��Z�G� Hń:ڒ��,�Ie��o;��mI9eG��xg4�U=}��!j}W��Ĩ�����+~¬h�;{���v�k��z��ܶ��Aոzh�'֝����!�U�E�^��$n�r2��/Ҕ����]+?�tm�jާ�OUl������0���2�y@C�3Ŵ�Yx��:�7Ӣ(�����J�� ����\;�����P:fh�H:�r��$J����3��H&�(��^Ve�ӷ���Q��zw��m]{}��ݽ��Ll��T��ʝ�:
�@X2c�<%594�2��:��:���M%�I��h�P�g�,k0�3+�j��s�1�v,z�U�(,m�QH�^���r��d�]
Gv�^]	����@���N��Ӗ[�d*�X]��K&!�]"q���Gv<5��k{����-����tP>���� ��(�f�i�~0I_D��z��P��04�2d7��ڑ��;f	�G�m��q�l���ٸ�����>��:�Qaa���3���n2I+Ε����_�Ii�5ct��4��9a;��W2�E@`}� �N����x�!�5!i����Â�L�TA�ԃ1����rb��q�n�RU��.�0�?y(��QU�	ͫ �3lő��s���fr�줹�5�^�5d��'̔zG��p�J�2�`?���s�.?r�V�L��`�.m:�D�]�����٢���G��jfk$�!��:;	�A�H@�|e&�~�D��K��c�UY=�D(-�0����`�+���dv�k����`h^��7��.l<�� NԘX��{��t�H.#���"���b�(E�ߩ�T̂#~+����7��5�����:EbcJ+�s��|@[f?Ox�jilҶ��� F�](��j+�7�x���.n��)���� �bpX��Z�B�,lH�=�; X�H�ZL����������H�aR���Q4RnU�P�u!�3�#���5e���Ь���N��`B���v���C˞;u,�(d	e��T��w�b���4`�_��Β�©���%r÷և�H�O��L^mA����@���zw#S����Ch#�Y�	�*#�Z"L�Tlƅ��f˶���rlY�۪&0�������~�D�TXU5�Eo@��ߔ��׈�M]��Z���w���QG�nի�u*���Vwke5��j;N�>�8��`�J�}�X%��S�.@�@���	�9�-�'"�;G/-����>2L�9\�Ȩ��|?���_G��ɉ��"v�'�`�4��UWӭ��7}�W ����v.v�XJ~���ڊ�L*=��}��i�/�(�́�J��-j�& ����Hr-m#�e?�'ZH��!�GcIDp�!2?�������v���n��
�^��ٗF�s?pN<s:�G,�oY&���rɋkƠ��*��9,7�#����&w�,H`�&p�rg�����1:�ܸ`�M�� O]u��BZ��m�%k<A���,0~.��ј�#>��Ⴁ�X�2_���v1���CG�����'�;H>8m�H��]�������Y_���Us���>����
�Ϫ\�SR�T�� 32)~aJ�%�x}H���R��_8/�%8�?²O��Ԥ��ē���;ϹC�;��)~?)��:��]䓭��њ��ƵX<LS�w���b�������.�=k]�]���v����e�;�?Kb{�z���J98�Kk��.�B<w�ϺJm�2���ϭB����/�6����H=>�\vH
Ӄtx���N e����4́��}��@S�N�^{��}�?���.f�G��"�9�~e+��սܳ����M�e�z"�Ba!�!�h���ݽ��^�M�y튰ڲ�֮*E�W ���X�?�?]3*�c����(Kc��Ur]1�oW��O��݊��5h̓�Jm%(�WQ�2u�d~���|1��пᖿ������VF�"}rR ��/���+���B�:����tb8~��0�p��6nF��g'�MK�Ƞ8���IpY���pm;�aR\��B;�\mT���-��Ž�)8�ul������WQ�L��o�M,]3ȉ/�S��=����'#��_���Y!�H`�/Q,��nCW�9�6$1Ք�V]�a�Nc�<e6)�?\�4�D/�����&�I�_I�Y�g�����T���4/v�U�7��Fy$AMh�)Q�y�d�]��_yX����9��bA�.x����������G_|�I<�
u1٫<@	;5*����֪[2:n�/�%5Ӕa�N���Е�ߵA����>[���Re�m.�!f<����(X!�7&拓0>�
"xf�Yh�89��x���ã�J߾����D��M;�W�
K�8�K�T"�>�����x(��n�n��%������/���ǲWv�H���s��ML�'��/�_0��l:{"lv�M��l��y%�2H(u3���6Mx�a`�:v���b��l�q�2#�<��C�Ƥ��EQ{}�d�mR'�;�7ND�ը3W��+XW�I{�ۛ�Yt���M�w�xF�}E��]f����nq<J�~�uz��jE�3�᫟j��Zl��|�t��ca��ɑ���kW3}��"��B�)��m�l���HI�L%�^�tЍE��@E�v�/�e�("Rs餸�C�P�0���r�c����km�uRX6}��S�Z<Y��XW�@n�<^�[Վ�*��Hb�Z4���B<���J֕
����s�����C�Sup���bϟ����=�i}Se�W&8a�������BX�G)jK͇u^C8�����XX�ma���댐���x���5.��E��&�wxk<��K��2�e瑶*�_���Ab�p�%h� �l
��%�Ӱ$e+����Q��}#�au$��e��C�M����Ƥ!o���N�J �z��Ґ�今��_r���p����R�1d_UG�}ߔ[��[�����'x��Ϊ�񛖥��A�8=M�}1�^����ƅ��r�*, ��rFM�лl#'�zj,��W}$�}�����z*��/&�
��Û��s���)�,�����wHȭ �A��7���6���L���`C��n��cI8��z�hq�$��UC�?�n���Jm<�y��c>�EV�pZ��}�Z��QT7��  Өc5�k�:���rQ��ql���f�␅���gj��Y�G�����dB�����Y�U$��{X��h��V���q+v�p�r�P�[ $s1i�j�;[��	`��j-x�^$�a�ˠ��)Qd4n�4�f��`�"V��u�Ss��og� ҦDZ�RM�P�����Х�X�F�˥h��qhCz����K������'jNw�7� ]��|������lT!1�Q:h�l�
�Y+^�%�%���F��%闍�J��M�/@a�ɘZ-Q^�Z�������4���l��ӭ^ذ� j
Lw�݀�Ƥ-]��k��h�35`�v	�b�p�,SU��PNU9ozxMM~t��pk��v{!(����@㤮��JvhT�7s^��`�W���R��>"`��a��gR��������y0�pt1�l�$(�]�0U��/����:H��O¨�@�;H�sb�x_4�&��7�L7[�;.kIo@Ƀ���H�Ehs�k�b�H�H�[�������+mK硛����gC��d��?�棷���b<�������f/��A�}��S��u�3nA�������r6KpdˤrBvisd�@�:���t����i��.���*̌���㍋�E��^.�2��:���w�F睦7�?<S
�GC�>kɺ{-�J���8%uo���dS�G%����/�f�ȷ>�Q�)�g7�j��m$xoݺS�<��7�\Eu]ɷ��KBes}��5��K��4���#�Z��h�Jk�� ��E����#���O���-q[��{u�B��+��'H�ܞ ���� `~I����x6~�}]M6y^�٠�[�v���3�(�\"�k��;TWh$�����{i��L�1�)�����nɪ�;��,���������)N>��-5�����-a��b�t6u"X�T�_|�l��ߣ�A�ST�Do��ňo�$G�����JV�������0kձ'W=J�|Э$�|��k�C����q �t�PpTW�n+aϺ�ť_���@�	�DJo�Z@���b}Wp=�_��z.x+[B௕^�*�!��S��Ip�
��N�n+���v���H��iA]��*a���G�x�ό^b�Mg�����4��(A��UT3�x���f�����<���k6�B�Q ��e�[֞���G9��
���=���f�*�( (�5I_Z9�����r�xZ�X��)�J���Ѣ�}#���>�v��h�Q7|]&�4T�ٶ��y�����Zq��׎f$�V~�V�2�)���.����A2� S���x�V�xs����zI��vg,��ދ@�N�Q�'ʙ@��]��D>�*�����i�M\J�/��Q��	c�V�UOs{�2���6�*Ns�tN�����[{�Vr�(�g(�i��_����Awۼ9��j�(:��g�-��8�+I_��x� ������N��m!C��K``� p����^��o'.������pğ�@�j��M���.6��ы)P��}�2w%OA+�°�aGZ�v�n��߿ĭG�0���&�?B��'I��d�b�%'����'n�v����*�ޣ��|W?���ZX�
T[�+���aWf<=*V�=1�\ʤ�ǜ��>��
u����3��5v�|�@�Z�u�X~�S�:���΅#��}����V�w�ܦ�	�Z'�k�L׃�|^m�q�X�F�r<a��-�F�TyZ�Qt*�� ?:h��W��D�>��+q�����b=��e��s@W8t�=���nTP�X)J��# z���>��%;ي��Do�~/�o�S���H���̹�\����>O�˶hE����"e��rVz17�ӣ%)�9B�S�i������d}��J�����v�~�Z�w�^��}3���@M B�%�����m�m\έ��x���~���J̘�,mM��J"�ME?t���G�f��S��-C[e��ʢ�cTe D�+��p~�VNkT@��l�л��7h6P��k��=�hP�ų3=�����塏*���Il$,6��Q����C�R�g	�ς/�s$�'�&����E	d_�n���f^���3�<9����E	˰<IDv��/�/ⷓ�;���5����l�l���>�G*��i��gò�:4m��5���-Y��Hpy�;8�f\m�FR9�UjtUFIKA�J��븟���s~�󂖄�����?4q\H�tG2�����)�뷺�<��׳�.���݄�p������陳��@����^�c(�)k_�)�c%ll�E�L���_��,�F�i�K�_AI.�͇G9�|�U�YL��x�o����=w�|�C���� ����>��ta#��*�6�4>Mok�8�#�(�T��/�]Ϲ��'���DX:��#~�I��+,ݍ�)/[}+w �ٵ�(.�nQ�.Ü��xr	%�l�g\�|����n�����L�����{����TKX7����g�w��ʘO���������,�#��i�;MЪ�GZ��P��5B��ʊ�.�U��1��[�3i�x��lvc�M(�������[MH���,�5͹2���-�R���LX>�;�h�q��Ιc�����*�n���Ѱ�o��̓xy&[$�Ǭ��L��N]�_���n��,�Rx������E���7~8*���m�R\ş<}04�!�i/΋9Xy��-l�͔֧p�$L�.d^n7沖G�華����h��]p-�0�_,�"�r�i��2Gb�}�u���-ZJ��j*~�S|�=N�)�pa�d1r�|ӽ�c#�MO��-E8\~ 9NMI �8U�����3����X�B@m_���C�=T!��yq��B�ϐ�FY���!�����D�o?I�(x�4� �C� ���,��|�R���`��ݐ�`ˡY���L+¡��y��8Li���(F�����~�����A�UM��E��*��Z��ߌMvS����\�$�X:6��gv� ����Gc��+t.m�3�����\<��,��ԪU��]��ran�k	���s��tu���*�tD�A�V�u���.G:�$ot^���I������V�)���1	I�DՉ�`����ԯ79.���mܭw<��i4Mc��}]-�k��ڥ���W����KR�R���vI:��6,k�۱�,�>7�v���	�8�m&1�����ig�� ��� �rGt
ݦ;�<6��n[-�)����w��QX(
�c�He��4+пI��sL�
ƞ�Bݾǝ/~�0= �b��&��b��\̽�u1�W{V=��m�6�lz:�	Y�5x��CO���>bD?�z(��^�-�"�>�s����m��."eRB��OjI��I�v�o�5�Hg��_i�
�R^���6���}����
�?.���	���thͨ�=y�ڄ�����zS�6���:�:;���Y���娣���p�>Ɯ2(C�4y�O�0���(=,X� ]N���ٱ�'��ҺQ,�]�u	9�l�����I��l��an���M�/�Q�*��T�^*���Qr�P�K��h��A����my9	�����Wo�s�f0�s��q��*��t<*ै��m�����f�1�}�%Fn_fqh�~dk}0�[\�u=-~|�����Փ�_�*�U�~���{��)u}ύ��(��k^5�j�� B�8�$�F�Q$,�gP=*(&��u��F�qfv͙���5��5C���i�Jk�/*.'�ڦ��ʕ�/S�@�VHK���G1�x� B��9xEO4�!_���PS���4�ک�	9D?��%N�M���4��rO[�5�9�)�J�D�.������@��ih��d�H<���x��]���5�J��,�z&�0��Vr��2:�T�gЂ2��S�Z���k�o�ʲ5Rw�6a�D�A���˸A��2�_�sM}�Z����	z{��H��A,O�� n���~j��n�WT��f�K����\s�b�M\�����V�"<sR>��3϶{36���QE�� E�^���l|�K=��~w{��e�EW!�F�b om�8��y��`����4��ҩS1��K���0?`5O(��:�ir
��bmun�I��D(��,u��k0j~��ӭ!��kފ�3e;��4h�R���9��읮��6�]�Ҍ�m%�r��#�N�X��Z���'P,M����i:�
���+Z��Z�E�r#�txP�'����K��,�P�-W�1���
B$d0U�+ם׽���������p9t�J��ɼ�l�x:N��P>�i�ZL]�\�M����z�bJ�b��2���J���(Ũ,A�^	;��.n�E��N�7p�O�kf0K���U��CM-�IPZ����c��#��I�ru�����kո>�G�N���l�OR_|;m��ۋ �#�f��)$�W�/�S��t��4���P�����*J�<7^%vf��B%O�Is̯�]χ��HU?��}2yuj�����S̒�&�W(J�s�CH?\'�G%���Ƣ>�º�ԿN�!���}�voz��H�y��9�7��[���U�M6Y�4hE
�Ow�V��(�?�jٳ̷��5�@r��Do]���fٱ����*��	�8���K�	�XҔT���¾x/Q�������-\�2�a�����L�]<�O\�����I]��5�r,�?��o[��f�ks��a��v5֟�'� ~-=�S�L35Npg.�i�#O���n�"�YMI�G5�""h�A�v��q��!+Pz#�A�C�n	̓�5y� �į���Dq��ş���{_"�@�DӪ�B����<+���A��By��\���Pp���+��Ka�%`و��w���a�$���Y�n�B�.�Ԥ��-ų.7��Ń�Gʹ�����$��n�O\�j�f�-f�8�na:�$U)B�!t�7V�WL�2��5g��ߛ������}҉�	gM(|b$�BE����@k�3{�4$�l��Y�l/RYB���Vm
5�\�FKA*�έV
�6p�+�.Ũ)�|ʌ���:�ma/grt��1��|�Il�h�������I��	����	}v�3
I�yRMo??���<��6Cm5{Ʀ�� ��0�+wo[�naC�\D�,Q�>�����Ӟ� �Ky����N��z���eg
rߑ�5hn��T�|�k�[Kq ��ucc��"oBqr��
�]�*"�f�Z�q�МsNqU�M{��Y�A�69}��F=<Y��f�c�W�E��T�%,!p��:Y�si	aL\#�i Zr�F���4&v#e�U�L���O�%�j�����xD�k�:�Z�a���'��\s8�%)�#J��K��Ruy!��
�AcL��C���8WTt%������ZeAe�]�61	�
�@�7'��J�Ur��0@5q��A�<M�Uaޜ�ml�;!���k4a����R�O�r Y��/h�z]fY���f��ܒ�GcE��0�0��A�.:�r���|��0^���<0�P����ֹ�"ĄP�+�݌�-���������g,h2�����	�`�a� �w#[�W_�����������xư�l�fʚ�oB$b����	ђ���H~�1y��\��p���7T�o<Q�ww��:��$ޭB��}�rK�����"�KL�~�t?4�wiOc����L/^5雏�R�V�������������f�eB~Ay&z��cF}��lꢍ, O^��M?�^�]��Ir���e�q�n����hS���W�M�/S�$�9�Q^ަ����S+l��#�O3:��#�̓��}�z3����	�%2ĥ��s5u��z�������ƁsR�:�tiAX�ί����g*� �D�nק�A�PV-0,H��ha:s_;<�G~*寑#p��^��� ua���B�*��vt�Q$N�ɽ��Yn-���WĝU$�{P֢>B���V�r�i�&�������GHB�bSt-P�I/��G@�QU�����읇뵜�]c6�5r[�t�[�5�}��޹���3�B�g����A��T,��Os�l��M:9+����F��$Ux+���蹿���s��
�Zy�!�0D�8%/�Y˂|��_$@)L�3W䎶�C�Q�5@���<`�s�s�CR@�t'!74�o�Y��H���`���5� �H�oI�7���?�q�R�|����u��/�=Z��j��}�KO�e6%q�]�2}��O.9�C�}�o�H{=n)��v+�2`�P������.'�?	H��G�5����ڈ���`Ld���N�B����谿�/��U��ra|b�dQb�"�}0����|�YD���ʝ���;���Ղ�<�����w�L��c|�
��0X�Wܨ���������Y�T"�X-n4q��� �£����lƶ�X���;'���� QE�>L)1��Ζt/#�3qI�
IҀk���P�4�-]��>�:��Y�Êi&�z��w�~!�h�m�S��>����oEh�NE�Tj���r%��L�)�����I��9s��k�*Chn?���$�k�M�~9�ovW]�|�ă��G[wmQ͜��R��RX���^E������(ivAf|ǩ�.�N5=7�����t�.�l��X���jw7�z�?�1�����i�et*+3�Bp��NK�E���j�pye�� 0,U�����i�5��ѡJL�X��~P�E��SF)U��6m 4����y^��f�p�-��߽�b�<l��	f-z	pUۓ�i��Z�D��ZC99��L �	���*�lNS����|�y�,{!F�ۭ!W�^���-�1N���4{�`�����s�㢵Q�� q������Ǝt������,���+�` �p��~�R�Ax1mD "�/Ca�G��]l��~3�*�/]���w�bnG�-��j�3k��Z�{�׊ƽ��z����E�S��8&���?�6��i�O��Cbz����TC
�kK�A�M����(�e�O{���P	�B�u,��_0��&k��T���֝lԅF�d�C��zR܊Q��SP6g�B8���fp0w�To��k�c�i�>�L	�K�"2�r���-U��+c���:�k�!������a_��m��8n�ʄ�(�%��ݗr��ܵ�O�;�`$�S3�(D���SA��JP�	B�`����)�ò��%m�����~�+�u�~�?rC��Q�������\�l�B/��w]㇠n�^r�B��q1$�ik��o~.vN��ȍ�Qu_Rڍ���Y�Si�^C ����3����X���S���t�BZ}޼>�E�-���]���1)�^#JD��r3�tH��$��Z�������v�BK�0x\�F�/�w��f�)��5�Λ�%%��v���v0vp4���U���s��I�-7�f
��#�������5�q�+�h�̾ў��D��d�! ���S�'��El.A�̂�WրU�V��P�Is�E금D�{0||�xV�wq��T��X�z(`�|���Z�t�ߊ�t���Q��XAvYs�3j �&���%T ��h��/�:�̶���Ҥ�?�V���������D��Y�;N�Ý�N�7/d¤�P&_%�ʙ��)؎�f��1?B�>��'�e��{@J��X�4̛åPz��ѐ��0xT��F��+����*d��TP�iʜTo��C{�61�bN���DF�L��I�7�����T'�-��ٚ��u�N�m��D�Zk�ǌy�J�(*����C��G��&}f��W�F��Rqu��V�Ӫ ��L��f7��w�+L�Rݤ\�XuU�N� 󷜄��"���i�G �*�g<�_��� ��u��n_��Y3�!�J��e%�5��o�p\E��~u3W��îܾ�N`>jM��3J����TO���A���R��4g��X~Go�5h)].�W�f�m�X�����zc����j��D!��d�G���P:�%gm?C�6��Hr,��T�ؙ_=x���=����[���!z�}=r�Q-n�t�I�ؒpԑ|���բ�a��-�~�4�';�5��ㅹN���e�+��l7y���W���j�4�ңk,	�#';U�Д`3k��f�����Ԝ&cC��ŕ_� .�/�Ѿ����c�\�,�q�C�/nC����h���x�i���G�v�x��nO~�o�����1�)?1�[�`B��w�*=����[36�b1�W-HD¶��ȯ�J�N�u�:�@��>��F���'�T������0�*S�-�5k%=��}��5l��7��o���gd#?K���Sh��� �E���w,��'j�(i���k�����z�&]�w�)��>�ma��Z*-��mc�"��a��;�X�H�����ڜՠjk
MAӯF�<G�W�'@nt�W=�.��2D���	/O��[4�]/��I�
�2�׾-ѣǿV�l�1=�ѭ�9P��ǯv3`\2�O�р�^C�W��b���T[��M���� E�h�_��d�my�׺��@�Qs@ٗ&f����h�����jQ}�"�����g�G�T�6�r`�%��#�ڍ��Ŵ?��N�p���	Ӵ�Q�jB��F#iɦ���lI�9�a-��<|�� '%sU�$�����i>i�3�d������k�����ƫ�1�Bk��P�/��C����x��V�I�V�D�.h��hFA'էV5�q��D�*�x���$Rv�	�7��#�a�|>����2#7�t�g����1����ަ�Ӧ�B���Sy��cA<Z)�$/{�I!s���p�u���ލ��W*��2�MH�q^*�i����g��O�@�w�E�����0`2���Ge�cBw.T@P��w(lp���V���z���4�?���)���NV>ؕW d�r�Ѫf?c�-�RuШ��Cݻ�ef�2Ů�B��E���ڌ��m��S�b�~u��bOAN�b�zE˓?����=S��[x��"��yU�g
ih�J&~9��N��i�c+�73;��	P�*=yʕ6-�	Σ��
��/7��Ge�c���(��@ ��Jgi�Y�b7}Ğ�,))��������4�<�q.K��Q9�$���nq=����yL5���B�81�K�&t�����˙����y*���r��N <���k��ufV	;er��F�c��8��([�2{R���B����G֘Q6JQcݟ9��!���U�d�㬀�rQh�b�W��Â�u�`"�J���[��ޒ0X��I )]�V�f&�A*8Ѱ}f�8d�Nl��Y�k�vL�)�h[�ɔ����A�V+��F@ZQ>���ﬔ�(YkTǁ��}�C�-ſ�(�&���/
��k*�ʍ�,�k.����?�`RN�]k�R��&&Kz<DT�e����`�{��F����Θ��l�9�:A��DP��_��<+\@��"�E҉"a�lh[��s,��d8�F^-�/68�O��O���F�����3)Ϩ���N��FQ��~���%q�>F�}��$	�i����������q�z�e�K�%�_:k�F�����v�6�*��ؕfԑ*Y���QӮV%�"���Z��3r�7����?ϒ0�sׅ��!D��{=��s�ʫK���3�)D�/Џ-�g�Mĺ���Qr�˚���׋�(���Y��䏊�N��A��Z�Ycz��P�B5~-��ԉN�[pA����>Ru�A�uJH�ǽ�Ԉ��+⮺n��{�W�Cu��.?	�l�XJ����N��=��61����W~�C��Ѫl�"츮�>����:;HGc��ʻ��X����gd~�	��_J����@'XJ�L�P�*�/���ٻ��숅�8�;�f�|죻uy��؉�����bh}e0�''�~�O�Wa���j��Y�dd���U�\�|�)	����R��&�fD�얈�}�?���G���)��0=�Zb�pў�coF,�?���˱"`"Bh�S�x'��Y�nw��C"*�ɥB��Q4�rb��z%�_����2�0���o��Z�R�Gu:'��|��<�6@�`KAa�,S�;8���]BO���7�ݭ�7aX|�B�	��Fuŝ��~�]I�]�
(�t�Y�������e��S�mF����j�/�K���R�I���?�t�����1�4���4�}NC���+Q��:G�)�;������HML�4���t>Q�_c����&-�,��16[p�)piGȞn=��eC�		vuT?v�G;r����w;�	����d���f@�bL`�+Gfb`�r��5�\���X�#"R���֟������b'=�~ikdH�Z:h[ђǒ�}�C�][��+��r("��J�޳'��W����|�ƂŔ����@0;����s�H
�ԕ��]V���,�&/�����E�M��g\h�E2`G_����O�����	�.#���V�mW��u����g���HEp7�=�{^�]O���7�� J��s6�D��Y�Egy�W+"�
�@����[���l�.e�-'�Q�	`ڎ�ޓq���M����0 �iG#��l�=.h籗����PCUa�ZWX� F��4�%;��OQg���q�+!��S����Bآm���揟���L/��>�N��(�8�!7�;!��n��ؿ�T�od�TK������j�Q���x�dg�X?��f���'UQ)YI�"���I��֭R]&�d%;��T$�ٙ9`ud��. ڮ�|�'��1���zX������T=���4Aɕn��%�"L�Nd_"�t��![?��zk�(lV���@�@9m6�STY��B,|��et�p����[\�8@` �9���l� 12V`�î�}l%�0��]!���]���m�e�o���"kÿ`��?��)9h��kk��L�4�M>[ׅu#_��nm��R�QB��8�k0�P�\V�ƹL\���F��1L�m9ѪŸ|���I�Bb=�����t�t=G�KdD�k �v�9��E��6�'y�����������- R�?�c�j�5k������kp��Ѐ��O�vf�8q�=k�����1���@��{<kp�}��~kZ}�ؘ���)@�e/�R��2uܷrF�֜FnD�������`�s�L^W.8�T�PO�ZP���U���j�Z�����\��C��qt�d|���ש�T	��\�������ۻ�����u<�8RzW���+����?�&u#�6|�'�򙿑�F�bo��]�C�_�<j�Uk�C���Z��ަ�Jϣ-��5�Ѳ:��YPsoA�%�&RL��
Ч<��Wu������&�AѲq~.����@� rn ��l�ꝓfm�XK�k�k����cKQ�I�^;���	r�q�T��J<3�8nq)
��q�82@�Mwn�I�"|�Z�y �i��9��?�#e��8���Luc_�ʋ�Tݣ���ʑ�v�S-�Y������w�kHd�ߵ��Im_�t"s�\+EX��r�����E�a����V�?�����:0q�,U�l��)_@�BfnpB���Q�3��>�>�\ѧ��X#�L�W��M�`Zԁ��n�iū{�q�����'��vǲ��	�F��c��7����T�}�Fi\2U�%B챬G��W���.��}(-��I��^��|
�\I��ޘ�^Cꠕ�6y����{�~��&��g���_�u��Zlj����)=]��I4��W���r��{�9k����/[�e�r,.����N-����hqW��|��r�sU�#c�*�������dKW�`���){���?7iئ�P�}	��ӫ���p��	�T�caC:�T��򲒪��"Eg��$����){�vh.�[����W�8q4T8�O�X�Q���y?� aM^+y$�Z����D�խ�~�A������)�c'Y������ƪE�Ά�9>��iL�9�;��W�̧<w�a�U@+��.��=�R-���}	OW)�B�x��O��
 H���߼{]k��+1/�L9gLa�ξ{I�& ����M�Ъr@K�[�Cmc���{Ӯ�d�����i����~^R�np%�=W�$���A}Ք��{���پ�칸�"O?��I�s��C�Q)�D���֏Zn�Q���:u�g�$7\�GKWU�f�WE�W�d'�eOD�TyS����%�w]_][����EYYj;f{����G���]L�L���g>�ӳ��cr ���)����}2wN�/H�/F���K^|QG�N!y�M
��-��<'�_Z�St�&��T������v.BP1\�fcRE.���u����X��]��c���}��|%�-Y�c��Ñ5߰Z��	5�rX�������4�_A6�(�<'_��n�d_��~F��X"����*&�锫�C\ik�!��t��uRy-��:E����'�M�łp�"�)�S4���6������M�P��Yg.P]R/�̛��j����xI�����{z��_ �������!i� � �	hd���&Kf2�l���<�eZXw����'������>�hmؾ���ȶG�X&.�6�ї�
�¼�5�NH2Wn�dFAp��l���b��w��Y�����!�:H���]�ݠ���x�"lbS'B��TD)iUώ3P�,�q��.uN�=���3���cR9�)���g�9�&
�7�����X� ��`o�&s*	^�b(�������f��d�����.�Kp�s�f#
uZGN��4	`B}�Km}I�w�aQ*��	�tO���#���0��+�<E׎�d���+H/��ܶ�n\	;��9��($o�,)��@'��xH��ѩiiv>��#U��Ѻ�Z�O�m��*wN����Lᑜ����ʈ*p~�f݄dʍ��c�� �&K���&�6��,�]�a��<맪��=��˧�pۓ�)�z�����$�]߻� ш�c����˱�ǃǎ�S��+��f�$�n�^��(�����<��8�:�?7�c��L�EF[.*�=d=��V����=����I���w���b�Q�D[�n��ɰ,r02&	�77��2g�.�4�����m�Q��UT�+A+qG�;�rt�6g\V����h��ȼ���n���j>(Ȃ̂rƱ�ӑq��[��Y`LQk�����%7�n{���h"f���Zx
�D�o{P�bl͠�<@�g���R- tG]dN���O��W�bf
�?�xs^- �5�^�F�E1�㬽�[X�2���=
���$m�a��Y��K���w�As��\���E����<5�f�'<���fW�+U�3�J�j����:���F���{Y�9qr������v��������)�}�c�qb��ɰ鶷�����N�:��Íp���*��о�[p5H����N�bV��ה�v��t_脚���J�^�R�}�E�UC�e^G�����x�6r��@
t��Y��kɴ��wRvI_��dy��| ���0=��V�9�Cq���H�,J�;0u�ۣ�t�>a�]�ɮ��ֿ��	�׮�kK;���{zNw-�g[(M��iP9���nm����艐�u(�QR���o�YP�"6;�!H}�f��X�l�)YZ�l�R��܇�-Vvs�G��CK3j�AѤ��tʚȼ����9I�)p�&8��b��1�K48k1�E@��&C=Kb��O��ND�Qe�B h�.)�:q��i~Z��������
,˻�X��^�z��Qi$�3a)�@�X�~����P�Dpr"/�q��)�W�|�C�Ź��'P��{��d���Ga%W	XNN�=�%FG�
�h�x[ƞ�w<�(�\�%W	���0�7���k���7l���(m7�R"]�,�`�,fMrr^l��
����y��[q�n�:��};��Ps�L����0���F�5p��E�*�wV�|B!,����S��+��dr��vY��F��db��c�`V 6�^����yGit�?����)|T���W���?P����rz��y��Г���l��T�T��m�y����C�+�Grnܽ�ܤ�7]�f�А�ԭ���;{aX6BO�i����E�P$3?TЌ%�Iq_yVH��+H�"c�
�LH|	�r ����J�JM��2��j%����p�h<U�=U_U|�n��i���79{���#��D/6)��jϘ������Z���o};p���}ɖ�Sv�a
J�ɢ-ғ�|�=�%Ɵ
��pu�$pެC�,'V���##��٪�W��{ie��ZGK��K�S��������m�_d����,�f��E�H�ř������uj��C⮶^FB�΄F�gt�$�5w�a8�x<Si!�Ԧ}���]W��J+ޝ@J�����9z���Oh�ˢ���w/J��O����&R;�G����|S�B|F��]rk?���Wk_/iV�	��Pi$`���hu���47	%l4��f�/'�eVc� �޳Ue��Z�/�ܴy���K�>�����Z����+��O�C��	�;�Ƙ"o�|v�'Z�K���?�3���<D��RVrŲdVp�Z��1�5ؓ�+�aD�h�azĥ���yd���Egڊa�F��N[�Ot0�����	��OI�듹�^1�Y����֟�e;�u���K�C���wa{MY��4;�OT���
�W��<_9�b&��µJ�[$E���ߙ�lt�&���ks�8L�yh���������hO�e���l W�j�����i��G4�7��#�n�����}��'�$4#��h�\;�Ӛ-{�Z�P��.�Ý!G��M�8��%E(-�no�f!{oI�snL�����[���}G������`�Ū,N+��R-t��k����@R����C��6��L��v9my`�viL
UN��_kj��j�����gJ����iבS�89�y$!�,z��N1�h���b��<V�)���1��0?
�O�R��O6�z�]��b���&ن�" ����o��Qz���[��@�	��G���گ�b4Hm+�t���6�o�З&$�nB+��h��+�'0v����~J�}��Sa�N��/;�PҖa��I2��a��$����^����79������z��׷��:d���4btO����׺> U� �a����5Ny��RA�.���'���
m�3{������2�⺪Y���r|Wg>RQW�|��[��.,yl��	������n}M�m @P�9c���p�پR)�ud<�t��9y�jG��'>���+�R��_�8�7��Ym��nX�P
Z|�!e�p�:�U��# ���7dD�	�w$�~f�M�CVNH3�X.Йð�[1�=����O~.�%�4��1��n՝nDf"��8/wy��F���|��ڥ���{��6�RQs�����
�+"��J��)�}��>Y�C��4�O�|^%� .4?�M�d�އ��\��}��]c��I�?�Tn�?r?xBt���5����nݹ�1#��x����������ae$��Dyx�5%r�+x�Z|3Z��eF��ڟ���u�U���TVG1�;\Uz�G�Ԋ�Ns�"��"@��2Q�y����]oI�@I#wI|K�u���zd��u�b��A�}�Y!@�-<�*���
���v�L��ar�ȷ��`��/���Y�(E�y�Y|6稢�2",�߲@򐁎��v@����^_W?y��K���-T↰5�:���F��G`ѭ����;�*h����k%���{(��yQ�x��h�ztX��l#��|��q�Zl�ޘsιMX8�֟�ސH(_���W�cF���T��R�z����qԺ`~GHz3h՘)�컇b�!�����	���Pq��/��ԥ��5���m��ʄ�i.5W�ͲA�E\2�,@����sl�yW8o�w�GH�qc+�sP���������F��Coqh��;�bH�V"C�E�)�(c��R#\����P�\�olvu-{��J��Axpږ�nW;*�9"��y�W���{<�Ϯ�Y�[�(q����B!2��H�jJ���Dgq������4�<�܄Pj�;����Ǘ#�N7
��m�M���ȘDG6x���Ԣ��!��\�g�Bs�	F�ӂ�d"3�#�t�]���r# Y�=}n��u=u��梴ou��0���G��\T����6`;@NF����+Z�~��|$j�LtM�1�B>����E'J0���d�>��,m]��0�<�`���R���m�!�R�yG�ʪY��#����������^�K���̖(F���&��m�[P�=������+�&�W]�n�DyҍSg�nL�[���~I���d%E�d[k�pXA�31#�c�m�#K�">�e���}b�h	S�+�Dѕ*ٶ�\�1p��3D>	9���Q�*�"�_>���#����ڿ�� a���YT����7�lk�+����W�+�ǩ����U~w�1]���+@��c^n������# k��?֔���3*�~rw�vAy��U[o�[����ſ�0�ݰٌ ��^ޞ}'�0)�\�-�L��.�:.5d;���z�U����O��K�!O�i��H��I�?�ÏJ1���{�St�kvi-���� �N��[��E�&��)6�p�y�tљ(�Ì�w��L9��9AW��a,_�� qU�1o��>�
��i�4��T��Lۛ�ڔ�~셻��O�!s�l\�Mpna�s�fͦ��L[Y��D�hj�C���2:�����	Wk���Gi���G�҄����t���	�]g����\.�����@`8�?qd�ﰑ]J4_� �Ӵk�ј���)4촌fi�̼z!+���� ��ؖ�^Gw�.A'�n�e��^�ExN��78�Ԁ�W��WGu���X���F�T�nu�,C{�X%��`�c{{`��L�OK�~y�WY�Y�~y�Ǖ����$hO��%��tBH^��x���]�E��-�$������j���޲4y����������jjP�u�|4��زR�P������w���69�Z}-'�`qJ��W�q�p�\9��r�������4���E���cTF��&*hӬ��J�v��f���;"'V�P˛k ��W�3���J�����Q؈��u���Hy*7`=�֖�t#�lV�0��*_��z������������"h�T��m�
�76�����[
՝����o�n@
8@6�H3m��B�c�n�Υx��s�T�w(�hU!�#ɦ�FQŶI�ʜ�v�<�mT�&D�K��z�:��S����鲀u��2f�����yp#�:ʣ�Ҭ�<2r�|s�?�Оu6�_�	5^��P���IY�K�V`b���b	�;*��i�/��oT�v�Nof0j�QJ�9�������R�V��r�5/ M����jo��/��l���0�w| AzM�:"8�����~��3�Q^�)?�A����^��t�||~�U��B�+����ݿ&T}s*��֮��e���?���Q��xn���I�1�N:�����.(�+)�nU0FOK�(�|�����<�2X+�R�|śݶ9��r��3��	�{��}�f���$���3�>V�&C�}P�ӱlL�+�4�&a.?��M�?y���H~��MϿ� �6�����-<�8�����#�����U�D��a,V�jN�1s����hl;$,���0�v@L����Z�U�n����=e�CՎ��l��T6@v��Z�C����*��{��q2<6���D�����g>$�Z�Ĝߒ6?E�������F���ݍW�l���9O�(�yѥ����b�V����Pp�O��̛G��W,|;ɲiz�k�
[�nN<���?�f�@O��;[�BWOd�߬���.�c��ڧk�V.c�I0tݟ$�@�h?x)��Z����&����Q1�p���k�NuBO��
(=�{�4����R��[RXd��O�G��/�iyw"�Y�J�|���
�5���
,)f^��
��E�If;�G�#,��$��h��al��t%���X��Q#�8G�T`��-��&�n��T,F������ߺ��*����͝��j�1w,p'Dd��a)2�t�%�g՝����pā�R�u
���N�$�W�X�`O���K�A�B�W��g��(Z.�ґ���vE�mȜ���?�)�����~ʀ��t�ڲ%2�׀H�N�����t�|Lй=��B���J����灹�a
��׾Z��%E�ŉ�ś)?� ��?YgqHzG\���v��SșAXa�N����ʮ�v���b�SV伞(^;��W�XH���O*3"bE���O�[�.����s�Z�B����3_� ��B㸭U�s�*��U��`��y��g� P�E�{��i�&�\� a`�a�pl'.s\{��Ѐ;�`8*5�ȶ� ��)�r������R4�/�zN�"O�`b�&�JU��We� �j�����)����lնi�5�G&;!ǏJ��H0K�Є=��	�[�+��҃�U�0,����7��=(�hV�{�Ɓ]n��O����.>S����V�/1��,;�~,R�	 "�v����`� "!p�����^����d{#������Q%�m�Y�`�[􈼩X�f�����~��~)�Ny)  /����%��AH�O;i�%��W��#����W�2Pm�8[��h[��U8��N�d�0�;��5�:wAlK�����F?�el�ڰ�'��Fģ. .ۮ�%����*>Q�iv;s ���'�3��ZR��1�+�Pw��Vi�+|�Y'�ѨYd:�@���2�?]u !(07�I�IL��y[��!2�# 5w�!xB���X����]�p۴/U1�`��J�~���H�Be ?���zT�&~Y���,�@���Śj�Aؙ�ʪ�J�*g֟.�A`�ɾ��R$U\�8�d��L�>�� �GVF��,Y>�t�;~qy��:ڵG�v�"d1��pS�
��c��O�<hr���ȱܴ��f�A� ��X9���\��Vb;�?Ɋ�w^�E6����1Y�4U����u�SВ�<��A@T~\깫���n��kï|~��
9��t����"�x�6"��5�+�y�7e�f�C��``E�۔<U�3�8yC� �2���=�x���1k���3Q��nR#�<-y�O������X"���x���XR��m�qWI�cǲ�g�ۣͫ����V藞����Ӣ�
�V��h���I�X^�-��"�@�!��)��6�@0�H��OҾ�uH��2)��t���Ұv���O������"�_������ߪv?��J�9�M ��9^��*���&�`�G�o���4N�L���I��#�&��jS�����_��4�{cS��%�3v2���2&�A`V"1�<�H�PR4�s����\2�R)����w�yٍ�HU���|��V��015����X6�\�Q���ъ�|�Z�;���@M�!Z�vЋ���D�3U�f�W/�6e��j�V���P��I|9�6�p��lĕA��9)���L�N��E�;���� NЧ���B��B���&��tՐ�L��x�y*����+Ȉf�{���V����P-��'�����.&���	��F��5��Xce1�kH�+[�*�L�� ��,��S\���9U!@@���FI(	p�n]b�IpB38�X�ғ��73�ٹ�i�kd�߫�0��G��A��G`-�|ӷ;�gh^�Kњ�c�ڋ(���:�K�l���gW~�����2�)�.Xky�5����5�Jړn��6�04+[�aY���i�i�s��0�xQę�88%N����h�j�_!��@4���B�`T
{��C���²�)�@���nA'HJ��eGOy�������R��t4 ^G�8 �ׇ#�qn ,�M"?��Đ~w> ����!���߸��4��������W�(��� ����t�����HZ�wK2�"�̳�l��K���b��c#�
�����˨g���C���D�w_
V+��E_U"��1@��Ȭ��fצ1�N�\'���g_yt��O��S'1��QQ$���M�+R��x��P-�jؠ��f��G�����'�����d���]ި\Џ��Ci;�ӫ��D��ގ�;M�e��qwH�1�Vyդ��7%��𔯚m��Gу���W<�Yix=�h�6�~8�+�9�7�Og��'8�Ȉ����I�rKrm�ע�W�N�_��Ƿ�Zө��_���\��^�K5�����>��dG%(�$'o{V����x^�윅R�8i:vr��+$�:�UQz�t|�-��_
�N�z1�~���#�^�4�#ND��{Pa��ɞ�ǐ+/�QJ޻�lv�zb	ڼ�h�nA1=��(��"
�5��,�7B�a�c�]�HD�b��\k�
#+����(=��3'Do%d��)�c�`��=���7�`��W�7	��]r�6���h;{|>����3���<�!ʐb����L�qL�Slvd^���ӈ�_�`[�^�s���8�T�;V��욙��+S�1S��%�p04����Jm��WQh�-�\S.����C�<L�>w!�1$�~O���ʦ4Z!O���m$����&�V���u{����߈;|A�Z�= ���{$c���8W����֯�$�/��F,E3�z �k��'�[�_��5+{�ȴd���S�O�: �	�0��u�41O= ����b����������y\k�F�T�;d�Y �r�H-b��5�Ǚ�����D{��&�7�<dpӢfT�f��`�3�P^B�8t�؈���|ק��h~d�OR?I��Pچ��ssTPi$x/L$퍉%�̕Q|�S��	��{<=t�ݑw�U��Y��@���t7�u��u��8�bL�n%���a��l���`׿y��[&%��Wը��\/����=�\��8*0��<��9YY�.��rN�/X�c'������mlX��bF}I�b�6��eP�z��04�(kPV9�}Q�LC�V[ ,��'O��DSP��E��`������甒�=���l|V�5U� �b/1M��w����	 �K�Y��v�2���r�e�i{/�v�s��C�V��	��aF[K����o<²�!9�CS�>�&���{���'L�'	C^�X�0��r�״�#$b.'�kCϝO��9$��?�E�mʳ'A�S����c����5�(u���^����zw��D|&(��H.A�x����ځӰ1�j��)�ݜ�8i�t�����z7�5<USu�uEGDk��亿�a�4�:s%9��LDRa��rv!p��$_��v~��:I�)���B�B����$�׫�����|c��t�or.9E� �2� ��B�V%#��.=sH���[q��*��1��Ϯ����y����Q� ��b������R�ּ0ܝ�r���Wƈ.v�s��hK��䖍"f:�:%q�;ͮ��}�k�L���L+{��_��q��0ay������������[�S�Ƞ��������5�.w�U�� �ܵ���/#lDk�w'���%��Qja��:|&%/V�Qn@�j���\�q4��W�ϝI�W�Tg����A�t��>����S�m�e���TF���.�����3nҨ���WFeH��sL������)���g�Ճ�,_�F�s���xY6P�T{Xh�����\Z�,�WH�p�H���E���`���'|v
�"Ӿz-l�|=D�{i����=ΣѹDa�9uȾ�+���� F'��di�����Rq3��c1_�?Q~jR��dXDi�8��O��A�H�;�8SUd���Q�|�v���D9�^R�=��vyxX���%J�L�zL
�߳���g���k���`y�nA즚�p��a
T���t�Y���ϯ�4#��p���V�!cX@2j2v`��q~�%�k���o��p$<?Rn\����R��&��\9Vp�����8��]��b�Y�&�`�U\P?ߗCr�ש�\}�0^���^&��\��?���<�"�W��6�}��@-�3aYK�!�Sw��p��˫���u�f|�f���d�',�vQ���O˵�ǧk�>V�L�>�g�)�|ߣ����YdA?�я�ؕ��) �s�� �]�k��Kgg=���1V�ȃ��)I �
�A�q�u��Q��>:�Lx���ro�`L�l/�bA��Qq���֨7"�M� �״�b�pl$^�U$5=����_b#����rˡ�h�gs9�ގ�p��z����ڃ�J�i[gc��.�S����m
�i�EK�"+̚B�88cW��7E�4���\���%	V0	�w�y�1�\���f�[�Aj��<�CQ��r���ϟ�lKERYH����Y�����F�z=�ʣ�:�����D���d}ƶ������=���<�ʍ�F�v��&|��!�81n��j}�҉"��]ȗl����dݬ����"���}����� �8��@�UE�FN4��/���
T�*�a ��F,`�ٙp���҄�� !Am�"�}����{�Ѵ���1���~�m�D1�i��oA�L��.*�L0b����%��0���)��[g
^МZ3p󤞳s*r�&vQ�-4�6
�^S/E�"d�m�� ,����ͽ�����\1���C�DD4�4��	�����oQ@6/�G1�l���H���yN�W��;�n�����e-��nu�q]���pw��b,�2-Q���!��w�ڛn��#���O��׌.�muk�Z��*rNd���m�~d� ���-��(@��&�#�
D�2�!N�&'�
�U4��_�u�=e��y4�Wzބ���Y~��8_=@�ގ��z��ۆ�5�΃
,�:b�v�� ��h2�J�qC�6��̶PZZrE۲��U�H����d�:ȆZ����c�s��2u�z�O�;���u�pC��� f(�A�V_���]��	�MZ��I�c��-��P�,L�ï���H�ޕ2$�.� ��C\O�
�t��R�B���$���^|�f����7��v#%T#�'�lP�ḷ��n�������u��I�7�x�R?�����މ��Ц�Z��l��1H�!l#/|Ƕ>r��k�] H��Q��G������LJ�b�$���]��"@�L�dml�1�����"��Ak�P������m����p}�]�Ä�0o�C�18�?��R��sI9�@���M5}��L��=QX윯&_&~�B`�x�W�Շ���?��u�L�A�	�)f>#����m��oH[�9�A��O��5�[���z������xOގj�����;5%%oXȖ�>B��jDA�Nb�%NJ�sF�z*����I9�=�ߙE�I����\�gr��1'vG�	y[±���w~�J���ڡ��$�R|�:t!�3��>։�b��h/�%���Lᑑ����}�ȖP�]�-�)_D8�%���=�TX����8��S����q2�/�@X�}�GS�SGָ�q�ҹ%�����4��)��T"E������*��$�ؠt^�����&F��l߼��ǥ9��<t|I�?��|�@d��/�Bu�#,��W�_O��M�����\bW�#���&���R��|zW32�x����x��V�Ұ�Ƒ�Th� c5����]�f������ɏw�>������5�h����1G;�Z=}�Om`-�"�C��45�	�WP����Q!:�e߼5};IPGa��0j�A���W�75[���h�ny�vᨈ~{K�6a���$�ʴj�bd7�ŰQ��Q3w�-A ��p�E�#�B�*�ujV��Jc_��������g����y��������4�5(���w^�d�/���att a���N;x�O�礢+���H��J{�j�G7��-���i���-���i�o4��Vk�����Ԣ	�����wJr��k�&��6u�
�@d�A�x������^w��J��;ĝ�ߛ`&T���_��l���k�wUJ|�HAv��ɗp�B���ӯJ�^�CzX`-�DG����d&Z$*�ϑB���Nj�BpΩ�����E\Ѣ�ގɾń}�iCɺ��,���>u����Q�zn
�H�7]��1?K�M��!�(#9(ٖ�<�G*{5���m$Y<�w�x����'.��@s-�%ܠ9eT?Fyy��$�%ܾ������g�Ih���Ә�M�b�ܚ�&�k2�6��BR��_/�ܢ��}�$1E�tԣ	�*{2�.�s��Z��q#�i�Z�$??b�*��ʢ�#�(f��Hb$Jj�'�l�Ι�$ճb&��*�1O�ϱ��`32�IAu��0Bk�u^y2t� rA1!�%��7�d*5m��)uȓ�����"Z�?��%0/Q�Zz��q��7��.M�KT��J��w��2�ꝳ��T��^I��<�C�C�K6�:��7�i�� ��b͗���X�><���{tos�;�a�m��<�F�����l�l��p�
�~��8���L2x~ӴI�w/��|�f��Y-z�%^����ʅ�}�����i�Z��B� � -�n,z����tP����P�J�G�$0��g�N뚔��}��� ��-�|������t#K���7��	�Uj�4� ��aы��̳vB��)�/�c�,'	�i�L���W��^��yE��[�)�l��<G{�~�vD��]#����?���^���G$�zS&	卑� ���f�@�K	�Z4(�SW�W_�sź��E�1,p�x� �x��d& w���`P��4��T��Rg$�h{���Zk����"��s�⼇���eG|��bȕ,����+��=�G ��ı�]J���콾���lU�&�U�K�� T�k�H��Ǧ�A��� �0��t3��#J9����ٻ�dr�K�-ڱs4f��U�PA�UE� 0��_����_��*ݭ4!s�������R��J�xLo��RȞ]��
��Bĥ��ϋN�3�����=���-���&�@���3���!��=�n�1��r��.
��r"3�.��ʀm[�����8���W�QF�o�}�0n�7�Z�6͘�=9B�?���SbX��t�8����}4%�~4)od\~���Ks�WR�Jb��z�Ny����'Ǹ7�1��m@&3xV{��s���e�͵b[�D�4� G�U�����������X�ǀ0��	��G�q�����m\4R-�.�6_xz��z3*/�y��Vgn�)j��K���2{X�$t���TU��:� ����}�.�UG��A�ϑH�8��g���L��R���&�mgl�A'TЙ�\=��uZqV��V�~f���%,����� .h�M1��g��T(��"�ބ�fmf;������?�
1�՝'l��@0Wν��}����!�&�/nFg:�?��WJ�iO�a��ݦQE��)2���0b֙\�VΨ)6�����mvr�O9ĭ��Hv*1�d��E|��XR�Ayx��,�!�`^a0�P��F��d���)�:ܿ���B��~�����J�%�[:�EO�`X;�6�ޡ`7���8��� �F4�1��!�j�����6Z��k��g�}GSW�n )���1^��l����?Ĕ�����V� �s���7�MP��'������!��Nг}c/jA0�0�EYY[1�"v�w�Y������'S�#�%aԘ��� m\ń�7�lB�܍�1�>�P��9ު�9mZ����f���{�����xR٬M���:w)� )��7p�I�)�c�ˏ��p�heg��[R3|Wx}8Q?�6��@q��f����K�P\�Mj������RM�BU�z�Ó���]-e�3B�R�u2����/�-G��l;��7�%_�
���O1'�d��.M��t#e3���d���i�xЅc�D�ٍYE�+�'�F��f�x����I&?�KD���w�� #��w*�A�C�� �<�M,�MkC��@۪`�DD��BA^z �d���
��jw�9��E޶������iE%����r<�#����K��(�_Z�y�<�����]����4�~P*e�p�U��%�p(z--�2�U���h=��U���p8kȩ3
!��0V,���sM-�*9��bSˣ��Gʌ*����O�;�eA��G��˔��������4�n�L�oR ��F�4��z���gk�oӾ�p�^M�M���s�C+�Ќ�J ��Uy�1�Wr�/�&�!���g�1�"u�i��9"yC�|�k�(�A�]'E�%�G���G-��`B*�]@Ů��
�����KE,�ψ]�u����ϲ��?_�(ԭA�6�~Q�T�Jk��c+�^�.���,���df�r7i�8��zj���"�+6��c/`�}����nF��U{0iCĚ�8EX�+=<�)�'[��c���.֖��k����S�Q�f%%^Q�3�H���1��,�YHUv�'{�vX���1��ğqGȄ�+��SxW�ƀ��H�5l,�<d����AI�o1�e�:
U�f�x���gIq:�G�f)�iCB�����82CxlnZ�z��\ã�:ƫ��B�a��ն1�orj�2�+VO+��Ƭ�J��SaCM[���☗R�p�j���Ql��.U�RjB���CvG=\��쑄�k�(�WF�μ�R�c��W��`+hZ��ȣ^�fשД$��O�8h�)�������<~��mЉ����M-Z?��ud3����3���]ZC����Ef��7�L��դ�m����Ȯ�A���TF�D��C��B��$�K3��!��Y+�]��bˢb��֎o���ׅ�Hj��zHg�~�C��|��ʧ`Mw��K)HLZz�����p%+���h.7�e/C d�t*/}{٪O6���-�
!ڦ��vJ���f?x*K�[�/�,�~��ܑ�Q4�=��e������@[2eL����W�ӣd�8|\X��A"�(��s0g�p; Ay%<����r;Y�lDa���b;}U���FesKƂ��WS:���O�&����$�`>�����|�S(�lq�9(��w���&���*w���~������W���J�y�ϱoŤ�
G�}�Y���<��P�B\Y�����~2�1��
�#��#�J���҃ӿ~/Vpݺc�%d���"V�	$��9�շK+�*��ڒ?{ȧӄL���S�G�=&��*"w�a}'(�d�5�XR��$�URΌ%#(%/B�����n?m���:�n ��
tEh�Y�o��(*&��(cKSl�i�"sP�/8�X �c�3�j"5�j��c,}*Z) �ʐ"�ߩ����b�juh�Ρ�,TbL8+=��4}n�<J���<�O���Db˫V@�t�^��y���HF�&�N�Z�� �1�����f���#+��A��NH�7�Zɡ�k5}������{d���&9���f���`dZ�#���9���]��G�����|A�0ͼS���m/��v�̬�U:o��F�����E�IU4��a��v���O��RHy��P��Kw�2��Ӗh$���E��m��M��"�*�5:[���>���\���.OX<�a+��>TJ(]�������	ހ����#���g���]�BZ���|�_V�� )#�rv�m��7�`���7�w�����fG�����A ��S�.��5�����3�1k�|�,��iI.�O��=`m߁&�$�� ٓ�@���3H�B��t����n+�!3��b�姒O���������fg#N�qik�?�u��LnFj�)����7�$ ��B��.��IՄ�G��ܔ�t�O��u0}/a�a+��B,٠]�ciZZ�f�����N_��d\[c��t$V�0�͔m���Yr�
�e6�+.�	���{��Ete6����H��>넲�������J##�Z���;�$�LJ�%�8��n��i��K*$q�*��n�ě4Kc-U;|�Cu�3S�45�	�'�[�����L_��L%,	epo+3�V#3�2��~�x��8m8����\F!�I���gec�������"���tǃ���Na�Z�릤𑡝�6�tꢩ��{My%G"�(�0Z+���Y�$��S��l7�"f�AY��h��{�3�	�t�JX�d)���?�h�&-�#��J������ڬ&�����$9��q���.��I)��p
l���Ebi5����܉��ӭ��o�fV��0z�<����
�gs������F@B�{M4;1�������'c;�ƣe{�|�6�s(A��Ƞ�7�;��Ն`r��H�+���v�%$2������g�d��@G��?Ɛ=�l�o��Sqy,IR��,|U��]�*����W9�Q-��AոQT�ü�Τ�@��?b[ɏa�p.�
�[�����M�i�sg<���(�1Bv�RR�����^d���c����~D�:fZ���bBfP()��m`���,�>U�g�Pb�O�6�"M�R��Z��j�Э��rԊ��"�exv�b-�_z��]�'���A�-�^��_X���B�?N���S$�Yľ:���uy�0���=`΃��y��zkcD��J���z��? %a��d���k]�g�K�Qu���G��.r��0tķ{�!��A�D˹+P	I�*^�?M����S�,��oZx�pp��04����r�Zq�\4mA�᝵F�e��i�hH/r���S4�z�»/�������a��R��ҟg=+�,JR�N���v���VNP���KMUI[ RtD�psb�� o�GOx�VͲ9"b|u������߆���}M"����W�, �����?岬�Xi�n��}��C��_�b&.�!f�r�m�3���+В��/a;Yӄz�����i�������g�#Cϩ�18HH��OOVG�a�7ҿ\����.�y2ԏ��R5���N�R��b5�<f��uz</�F�nGo�P(����䃡3�t�>D�H��7����E<D�h���:[�CjKj�'>�l"��Pk���]�9��}ΌM �"4~��w<�٪3E�4ʖy���?�BIҠ�=�T1+��^thi@>1oiq��)��E���lԢ��Y�����|���=t�s�F��(�/�t�{��q�ى��U;�`5>�����ˆb?�-��	�Z]+ǌN��]KzS��p�96�^�@Y���N�!����R[70���$�+z�,,Կ���>�l�՛r#��5��Tҽ%�N\5��H�U"�K2���E�ǃ�l�������h*V��f,�d�g��b(���PWK�m��\�DrO�?�C�.=Ӱʦ�z���y\�yZ�������%��,��K�<YmH�3�l�����I����%��$ ���-�C��Ћ�R��.��S;:��o���Q:ɝ��h��w&�}��2�xV����s��{�HK�o n�Y�Tӓ�[e"���,�U�1�j�<�)*��a�{[���C���#B��˜��� �ot�Ɲ���S>c�H���Vy4���mz�dP)�Hn�*��v(5 �#�9ܠ�`�lJ6mt�?`�誕҆�J��0�xo��2{�2�̋�ih�l��@T���RA����c�4��5�L��9p��� D��\��}?H?��d�i���1�oj��i����m/Sa\��ޒx�o[�k0P��fU��k���]$a�
�@q�R�*;�%"����鰯���ȗ�>U�������6�C.1�����,�i�">�X po�9[��r_gn��<R���5���*����3�Ԭ"���|�Yy[\�ݡxb0���c���r2t���΂����nZ@E���9 "�/�^�H�i�CÜ��Q��U`����,�(W)�t-J�K�*��m*��$�c����%VW�ؙ@�4��gX*qӇB2�\�%�o�=�<�ی�z΁���I��1U��i���*�Q���l5�Si�0 r���?�S��S�[�C�������2��N���ꯢ��>���#�K�	;7PxuH#9��f{3ug����N!�<�q)�y��c��gXƴ]ߞ��x��������K���M*%.K#�u2�
�"$�������Lވ�/�aq^�!�z$X�ہ��G����Zוɏ��]����W�T��G�\�m�9�E��Lg� _��s�;n��}�`לTҦ�+4���#�C�9���#ƔQ��l�i�Ǉg��`H����?��$��rV-�p��D&�0'
mq���0���2*���$�C����,Ǫ��5<���K�q�ަj-v�EL|1;`�=V,�� כ($��4�I��d�m�$p�f,� i'�fx�HcX%k u���"�����{*�Ų�O�������>u��܎�-�W�k�&�E-��8Ī�{G�ޕB��9/�d8��ü�6U�;Lk��g���!HeMQ���
�lژ �ƍm�& a��S*΄u��4fEc��לݞc�D�zj���!�m~"�y��'��
[E����
���C�M��4j�~S�xֽ�H���G]�Ҡ/Mq��Y���)CW�	�>H��<� ���'�:�Q�c�T�U�)�>i%���U"�������B�;��B�$�����cm�����$���,�OeK1 ���$«5+�7�����4�XI	�<��0X�hM�%?�NR�81fA��hZ��+��u���%
������;I�#;����(H�xFH�QF�jO��S��R��V�cD���SDƃ���0�랭���D�~�~�>�G�pF;ĺݠ��u�[�CT��&4�_!v���K.Q��0���NR��'[�<�%�D�/,$ZȹFRRI�vss�Z�[�@�>�&	|Ȕ3A�6�mr���Hf����jbr���}�%p�qDUZt#�0|��:��6�=���f5�����Z�Q�g�dTWH�K�l��)Y<C	)�Lp���D�&�؆�cu�;�0�����]��Z�pU�?��H����70��U�MR	��ʜ-D/ā�#��B+N�o��pn��%�P��� ����e�-�����m���p��aGE�3�K��P+�(�mo�ӯBV�>�Ap����!��s�yy.H�b�(_�H�?t����z�<N �GLH�F�8uʂQ3H?�*4�!�<O��vF�u����GoUX���;�t����r��Yd
�J�5�o۴�����@��T����v0���D�z�~*���+��e*/d��z:/M�4p��١=��|�%:��d��S-�I�JJ����+F �Ц&:�٤�~%G�毿͜~ُ��Zl�Gώ���X�+�Rǽ�@�/���{�Iʝ%��vd��X�8�F���%0��&/{J��0��p^�yX\U_CV�ϜSc�n�饒ͮ�J�۠�����f�,0�Ϳ�=�3��iYY���4�����#5��(�#Y,�˴�	�㟼���&�
|X������η$���Eo���n����2��3b�=rlKCƆS_b�Y��Ѝ뵝��@~S���A�ӧ��HP���(�^#gR�R�(�����	�s���e�$a��A�1ܮy'Xδ��VK�DE	J����GX��Sᱺ��d�B����Eb��Ж��ls���S5�g qU��:5��߹�K$�I��-.�
[9��	�]?��5V>+ِ'|����d�����E�ڤ8�}�����Swi
�/O*��-ۍ	�32#D��_<�����P�Ռ��Qh{�R$��d���R��wyWqL4\�O�P��XMFШ���c`���*�MC
kf�h��K�_�����n_�7	��[�9��N`�X@沽���'R�}n'u��aj�D{-�Kk�d7R���{��;R�{�z�EX�BĽ��2��d֘]�ږ&@�@P��\�`᢮p���oi���A���;4Z�S'U,��Y�,G޶�ߢf�gC^�^qfIU��\ڬgw&�B�D�K��1��ZFtt7:���#-�FV���E%��݄�ruܧ�'�[
˖�@����d0Rh�[b�߭�� P8�tV��vu��@kPP�w_�����N�&�����9�<���wk-�i�M�d0KL��&��N�&-���}2�q���!�@�D�K�;8�������w�������h�q�p��z��D��m�����|���s�-㘉S���hdQ��,��{L�K�5�ُ��4�s<;�ۇVA����YޣEu��h}y�:ڪ9C��Bh/�O��/�ve�)��J���IaA깷FB��ڇ�D3Д�H��̗v=$���F�AI�u��rՖ�.���(�L!���:�z:=r�?���tL~5vp�a���8����/�IY��i�i�V���+v��>���zI�xi���@��	z�8��ĳ?��yp5nٰ!M ��XcZ��O�Z��1�{��<�r���w�w���5����X��FTnMy��%���֤;�O����r� ��rH+^*r'��x�<���:�(�}c>���p����H!E������8z�ffk�Y@����g�ɨL�3�=�t+D3t�,�J��=��
��ft�:�5�]��Y���R��]�K_$���˧S���V'���Z�����p��J�P�PB5mH���k\d�?	�H'�РR�u�y���<q3R%�"��t6ck6���#��S�퐧8@�4֞�����n�X��U� �KW�;�F��@[��TЏ������QƖ$��������/�&��Ũ��zK¬�jͲ�uGo!00I_}��h^����������L1U\N£��=�C̩W*����0R����5`4��M6���2SC���B�wb{vP�b�KB�GX\�u���4�0�J`��Â�۞�q�����֑��$��c�V=�q.Q�s�) zU-��Veʇ��i5�h���3�N��Aq�2�Qw���\�f-��b'��׈�X�uMʿИcl���U��U6�)�o_�q^ɽ�O�凇Xb�Q�0Z���
���yk ku�<L��x��g����ĳ;zn#O�:-��u�����=V��J�T�Sp��� ���>(l9w]��V�D����j�^��;m����W>*�䂔�3J��c�9GB�$�A;�ɉ獃��H9sċKe���^%:?	��ύ�W���RT��O��!r�����K�6�bU_�����Vd�E��XN1B �"|`BS��Ih����|	�M_��x5H�0��Yo8}P0(���0�����s�u�k���z|���ZV��t�ԭ5آG���#�l��p�~jw�;4�%d��]t� ����u@����Bs���|ȝ���RG�E1��H��Y1��YV͋��	h�̻��C�+���S�e<Q[��[�ЇĘ���<<��� �<���c��-Qh�D�5��ɷg],�9xuD�s:%�7�ɋt��׏�s!� M;4su�IHl?<{�]tP{�r7�X�� rXˑ������:�J���������8H�&���W?n��SQ0���!��n�7�,�	�18��)EB��t�]]�/�ʫ�3�n׉�l��%�E�\B�|�l4[<0��!���Ԙ�r,N�����Msܱ�������~��-I��ŷ�\�j/ٴ�z(�d���0�m؇�H�e��`���D���Ηf���ru��`O�$	�؆��W�]��#PsX6NJ-�=K�I�%�eר_Q�4G�x�"v��[�(��ǲ;�S��B�{:;k��y�>`ڟ�ӛ>�^��N6�Io��� �����*%���k�j�^�;DS\�v2[J,.s�WM�������Q�3x.`�I���M�<H��X� ��l�f)�M�$Ef=k�=r�_�>�v����U� mWQܵ����8$&3d8�ߗ�i�o�0�B�9���_<���CMmM���u찭o��x'D��Wt5;'E��~^C��ƕɶ��X.H�h`}�e�N/U���������N���W��5Wj��E��҇~@�E�Z�m�l�����b�����y^e�:��ޭ��o������7?b)��;7!��~\���S�u�����͢c\��q�ۍ;g߉������惆�������$��w˦|���!u�Dv1'�b
�V��Y���#M�F�Gq�ҹ_����(bq�	���O�OPư��a�B��*�c��(D':>�~�yc@�������[��Q6���VO���x&�st��H�u�O�<��-�_��(
��`�G�З�P�[�©T1/���.f����)�W� �r�ZَH�7�*�U�	�;�<�	'A�N�����J�;�S���i&������i��G`�.�o�L��T���{����њ�_܋�x}x�Q��a��׃�q��¯]dX�{,ґ�[����"͙@w�
��ٸ�!��J¦ԓ�O���T���Ӣc)�[~��A/��Z�Ћ,ܱq����6���G�!�Sϭy���jۭ�KId�e����RI%�(��XIw��pIQ|��F��,�hy��!յ�b]�Sfd+��zL�Ns���4>C7ec��X���3:l�}�3z�)�<�D��&����*�W�J�,Ґ��kv^�w{�Yg����9Eߒ�@��CycWBk}������g8_;��R��?��/D������
N�8.A͔��0�jǟ!���k�e�]�ш�]��K\�,as"�vЖ�@uT6�e��$��R{a�L�J��.�{�bC]f�H�Jsj}`9��.p�������U���R�����*ԥ薴 R�`6�HT=E^�9��8y5���V[m����AɊ�:��p]%�4���\��SCl������g���vN�}��NN�E�/ɦy��9�A�h�]]u���jĹdCR��F:���3����F��Y�thy3�z�'���e�t].��O��i���x�O6�1�9�F�ޘȟX�
�t�ƀ*Z�5�%J�p��J]���m�?��,�\��	��(��`�b��a:��
I⻹���6Cu���?i�8�{i�g�Y9���/-�gZ��80�_7T}�~3�._���f��WN��mu���!S`�G^��%���S>j�dL������0'T"��|a�]P<���Y��,�{�������� ��~��4�����,�#��#�]c��=��%����_�z%x�A��'�f��0��B���1��n�gh㋿j������3&|�C�)�O\�R��F�܎��?7/a^�ܨ�K��j���A3*@�@��%��p��C{$U�-�ؘ�P���@+/7*\E�: �FUw�$�߈����a�RV������ﮩ�\G����5���8����|"ڻ
1�e3�F��9[�8"�(�><�Z���[�]VmN�*���uu�:=�X<U�q/�	���~]G=y��9����m�Ul?�'0ُ!�x1�O�uǪ%_�,��`�E���S%0��*Cj䫪؎ωe]t�v��C�h�		�����"q}�O��@ <�?�4�a=S�A��p1ʂ체\2)�ס؀���F��^_��/���.M/	D��f�ĴRd"���Q2�lE��tz>�7Ŭ�+"zߙQ�fL�����D�ڍ6�܈�Ҩ�Powv�Q���g��=��I
�-�����@�ﺘx�W
R������f鮎#�9N6u�5U��D�D#��xg�� �I�!�VA���4�'����ĦvN�e)S��-	4^WPp�$>�<���1��?�`�V��.!s��Y�<���Zdb���˞�̖"�La�<��������쉀'�����-tl�0ċ��"�$A>�@5b$�g,`Mg�fg�{���O(<�?�Z�H�ӻ���[֊H�&LV�T]�*'��P�_5��+�O�� KFᗚ'�*AD�B�ˤ��2Kp8��*��>!f���	���p4��i$j8�h�J�� �M�1�w�b�*}���
��nLN���6�I}A>�7_�w�E�ś��U�������M��",�0�I�K�)����Z��|L;�#͗"�X����OK� ��@uc��j?{b�R.�7���E*�V2(��h�H�>�1%�I��O����\�l�P���I��ٗ�B�� ʖ��Go�j���<qܼ7ռm��/��5 ��.�U�[���6��{����G48�i��vMN�~L6������r�Җ�]���3�FEnG �b �yE)H�Œ�%�8����ܣ�9�eD��o�"�|hж�|c�M��]kz�bRnu;9�;f�8v �)�;�3y��$<BW�����D&s�2_���Bj`��z6 |��df5��?�����|lŶ�40^����w�<�*Vm����=�`�j��}O�O��ã�P}x1��(q{8�m�L�
c˄'�����0�����oQ �5T�z�\&���7ў� ���蔍���9�4�Q�	�tL<?F؊^�'�OS[�m��W�~/�~��`�pPt�?�,�(6�������5�F�ӒX�+t+��N%��(Ays�g����[�g�#��w}�/��ڥ(<շ3�n­J=���a<ǐ���-�̋v�׳�*T),�2o9��]�[5j���1?��	��ήkU�<�_�bULT|F���h�[�#�Z9�;.3�)犬�zy��s��IH��{���	0�Ӕw;��ܫC�染�/9T�;_�@t���Oҍ�K��H�?<1X���c���{��%��V��8I���B*��-��ֲ���&�1�ԈUֳ�2Y\[(��W2>'�[}��a����7K��i�Mm�\�u|��)�i��,v��7l��ˆS�R	h'f���G�� ���Yۋ��c�z����,���k��1"=Z�ؒ��N3�5e��K�'a�$���b6���]�#m�h�@��P��{Z`f"h�����/�|�-0)~L��^�c��\_o�m>�.Vz�f�	Y��"2S-S�B�c�v#	��/Uk/�I�ش5ӎ��P0�&�F�N%�Z��/��g����%æ�؈��iPm�BE�YL��NB�C0��9����Cf�f�{B�{��oȕ��$�
�����I���OJ9�\Xc���X{�˅�������[���5,�^���tڧ�Mu����^ir^�$eS�I]k��f��x
ZV�.]��Dq��B"������w�k�/8!p7+��LS7���f8�<��D�g� "<)�<�e-�FC>� ��<X�?O
,��4��_e�1�1^BM�J?�T�tA�� :���PR�f���@��=�������>g��Q��Z���;_N�u�hMB3Q�4��?&�P@Qp���J��W.����#�td�1�hI(�'�2oJbm�24O6���9�&<�E�����w��c�� 6	 ~�������26�q���G�)�O��I�=��#�kq2.�����d�&�������|!v3Ŝ�[]���"���/̽�2�I�s���+�n�8�ػO�]/e����dVDۭ����6�9�k&=LW�,�W�����]�X?�ߌ�����7HA!f�:�⍿W��#�$H�D늝�WB--���d��*ħ�����Y�U�[-���nq6��F"��r/Z5�oѯ� 8�E���3r���T�FT
ng@[�����ө@𑠯H��W�H�_~K��]�U8�� �\�^Q��0'g6���%���>���<O>�rݩ}�eti������1���w���W#�t�9LZV��"^����qL�}x�:�&o/9��1�l0ߚս!���M�� k��Š��{4x����(v�9�✒��#�Q�B�Is?s�;4����|�\[Ӓ�־��J)��Br�͐�2�jFT��-d8�W0]؏Z��$Îݵz�U1��n�����&�-�/���6�g4ԏ�� g��.^���y����Մ;N��.Q,�~ E(IW��V�jA�P�9UGƨ�gH̏و���o����{C8X����N��5� ��gzeJ紋b��dyչc�ZO쐺)�m�oώ��h�S_LR5����<�6�R���B=�=��ҽ�&eo ��W�y����k|I+cʢr@:u c�:�סzVu����eO��uBѱ:�q_OO�� �P���<��Ob���	�Y�\?��'�ؐC�k�-�g��0�)�:��Q�EJn���W��s�M ���)����T�� �)�^�ɺw`&�B��g���P�F{[�P\F>�Kx�2"Uu=�S��p0���aZ��Н'*ՙ�Y�5'L�3@�X�sj�����2���F�T~`qǶ��!��7i7 S�����%��lq�� W��0X!���F!	6��k�[�����G'/��d��B�|�E�MuS63�5��H#\��\�}�4�ذ}������� o�v��	�m4/6�������/�z�c��#�.��v�]���=Q��3��Ǧ����	� ���Y�T�V��,2�o]{��+y�������,c�iY�z���h��<o�r�?�8���S�wHZ�x���Rk�%��t^�����]_�U\�蛐�`o�aT�>��
Tel��L��-K���ތ{�p�HV ���q��R�S-�g���d�v���J����IՓs �
�0t��.B'�{�<ezp��j�D���,�����
��)������������?���''��K�c}xg�uR��"��p�m��74�eI�<�5z5�x��"Q���0CS��6�A�$�Q[lt�"�%j���ژ��C�DweB��F]l���9[R�h��T�5S�hܑm�%×���H9N�,����� 8:�4J@m�a���O�����F�f�k XZ�~��L�r�I顩���es>|o�~�~t��h�B��Hl����	����9�E��{����wJ�R��-���=^�̚��1�.���k�{?�5���yϐN��:tא�����}���y��B�kI��]p���VF� s����b�m
5�jL@���;.vX>O"��� a3nD���N�h�vwpA ,;}�3 ���9*�<�V+P������e�f�d��a����W�G�~Gsc�]���-�o��^�6^��rhp���x�`�<���I�Z���Zv�5�P�4r��F0傠����;E[Aמb�Uԙ?H��5�?����3���M���A���oС}��5��b �en��L�2�@�cqit�y���O�]=.� �n?{Y�� �ش��P!�F4�����lǪl $`�Œ���
���	O���,}S��GxX٠>@3���[u�>!�4�BD�0a�0j�.M�슷A4�iF]�x�y��it8���%(5t@��6D��&�|��׺�|HĳA����BƦ#K���� O��3����8�\Y]/C|��*��>��Ϡ}�ܧgP_͌��Z�N�&
'wP�� ��O��e�H�(ܟ����µ� j̋]IL�*<�l�Q���^.���nW�NdOm |��?_�?��3��l�'��?�-��x��7.��>��t�_"�O�~��1_ao�Z��������M��\��T�K��ix��1��\�Ij̆9�Xu��y�[��B�y�]�\��w��DAmkKkP�gw$}�䥾������4�+�ʖR�/Su���� �ֳ���X��4ఫF�}r=��$x7��̮�:����-0��*��1� q��qKO�F1)6�u7��U��zh%^^WYz���(�����+�dr�&�^�G��.��T�m�_ճ| �_���`�,_b���eɓ�SsNzS�:n�#�T'
l��oOT�5�i'	E6�8����_���� �ޑ0Ta�ҞA1�#�e�$�qa5�[lh�����<�?h�ǧ�!�F��1�H7�i?0�mE=j,{�/��ŋs���GP�+��C6Ǿ��8�p:��DE��MM�,0��cӭ�u����%��� %~:�Q���  �H�� ��j�� 4�QSBJKF^cED9�qt��e!�v��3���L�-姚tt�OY^�9����LߞL�7������0��c����'���w���9�1��g��}���8��*�s��;'�7�yA��Y�eu��j,nk�'}�$.�y���-Wol$Ev���lq�kS����QX-vjG�#Dy���/��D�����m������wc���O��O[�"��j�2\��^:HZwk���m�s ܍��M7���+�w���p��kH����@O�c��޷ЕaRZø� <���T��p��{��մ;LX{\�R_ү,�hPy+���L3�	��ZY�]�`P:�;����~C����R�Dg#x��z�U��D6F��z��<�+�&��ԕ�+=e�4Y����b?�rz��q�Re��jd-�9�_�B3�u�����@�a�
���Q���&H���_K��.�&Z��#����I�^�3�ժ�oC�=�8<Ó���>��}g���������.�A}����@x��b���Qj9���/-�2�yH.)���2y\�A�l���AQ�)�-To��:a��Fj?=bt@|D�Ts��?2����6.,��S��h���N�v�kŘ�i�q��Y�y�Y\��%f�l7��2�fd;�)۴M�H�(�_B���<��G��.�,�/�������J�!���@5k�}��� ��˧j% s4�N@�u~ە8������M��ּ�ݠ�M��ѕ��.�~�MH�e�MB	<n�犮2�%�|��O�	]䣜y���S�V������]�o�n����M�m����Z
��-v� �A�?DI%&m-� zI��`�k��h��_�4l��: ��l��,���!�֥�jSCW�f�d��"1BͺmI�Ί����En-3 v}=跔64���Z�� c�)��uW3�/�!�Z����6�|��/�J���g�5�@6^��k�� 	��Ҵ��L,����j�~����ho�TU��E"�����9M��?d�]�� ��HaҌ�$��O�	��>w��q�PL6�V�����Kd�/������n�����C�Ū���U6}ᡶ|Kf�{��]��q|�v-/{mJ"m7�檕� ��k(/���Lٞ�-�CC9{- R����'�*��9��
��a��b�f���	��{ �8CE%�k�ц�;�34u�C˅Y�|>ؾ\9r�pʱv=3JV�\�F�mY	{�� �<5"a|�������Or����� ǳ#�Y��#��	\ �������g��S���)�
F��ϼ�#$H"�H6=h��Gyq~/�����b|����O{�����C/�Bm���Z��k��uW�w[�[˩��Oe ��#kv��Ğh�mӵI���	�[_Dfʪ���Վ�N�3h��l���4H� �>I�R_LP��/g3���H���,h:���Ja��_{��%�Ѐ�W6!ƿ�2�.�X��B�r���92�h�J9����ﴳ�g�aOv��!rU��������f��Jv���O�~��xtr%��!cҿ��-	�T�VwVȩEʥ;��'<;ى}ކ��ގ�-����t|~Z�x���U��z�퟼����4�3a�+~m_�^��H�f��J���7mǿ�>�jX��8|�(Fɱ�y7\+��VFa뮀�z���0V�ra��5�ņ�qd�lA*j�\?��Y3�1�O��6�!�}_vbK����R����B�,1��V��:Ӏ���4"/966�텉o�Wd����P�L��s��M}�P� ��� 'u�Ht� L��������������w�V֤��'A;�� t������?�#�_���0��4�j�zq�Y�@|3�ݬ�X�$��A��U�X���1�O8�5�ү�7��dͦ%q�7"�w�L��g�͔�{��ve��`U1�v�9ě��C=1�^��O��Qf�l.{����ֳ� ?
���6���@�I�l]��n�QU����k��2=��F��@�u&w�w0�Ǧl��c�ls�[s�>��b�M���o~%֣<���p�)#���n�����L�������o7��<(]��B�gr�I$o�
��b�#��u���$I%���g^H1��ԦPZ;�p�^/��yvvC�R���n�q]ZRy�OP�~�&�9gvv���uu��~����	%�wy�fܽD[/�^��])�yCL�R�]���&�	����(�"UiL���˂�w�����\|p�t���~���=jҕ �����)�(�CJf)�cɒ������`P����(����k}��$��+:��^~h3@����ʋ�M����{��z#�X���b[g��ݾ v�;�Vŉn.�z�b�D`AU)�[��$�C�V,��5*_�8V�������Ub� ����Xxe��5�.��z#f����Q	��!�K�?�}�cl��j8[�l��Bُ8f��0��i������{��g!�����\IH�L�]��*�Y����mp]Yז")64`@'yn�ep���DIرq8N��E3��S��`u\���;���/	�<m.�4���r+t� �N�~?���,�4v2 �3������>��$����1}6*�t���8�w��j�!�q��9��q��S�;�� g�5cC�ʻ��&w��;�~��2�g�;I+��~����s.�!8�nޤ�pm��@�:��i�e(�ض-�R��������|�)+a@����xi;�iQ|'�x�+�ͭ�k��η&�c��Ë�Mh��s�/��K�P�IS��i�}7$�V�dfP�-qc)�e���r�e�:�Y��IuPihg���Q�����fXa����}��%���:��"4ʈ 
�ܿ���A*������b������7��q`�2�p.����J 	Ք���=&������ �LR����NA�#���p��$v���C� X~{�T5�u����v�	"
�ﰨ+�P^��\|��rU����8������ډu��u�5��K�EE�V�R�sn��ĻԞ!)l�t)��!n
�C\u/��F�G������!�hR\H5�CkC#��>߸E� �z�˙�c��`F|��M��{dR�H�IQSq�+Y"���&�[�g�&�XjL^�U�h��K}�PG��n��*.�7������5��!��.�;�ޡ�.�l���*�2x�9.��:����~��v $W?�y�ZԸX���)�O�|w(�e���!���Q܃��u��i���̯�3͈=:���GH�4;_6���B7�? ��
���e�I� t{�zn�e8�I����X�0t�KHJ�����=r���W_�?Ux�U%���j6u��^�|>��b�@&�O�P���z������4���.�q�a]��	���'F����Aa]�+����;��;Ҿu`q��٘@1_�CG���^v!9�Z?UĮ�=�~�gnE�-�\�/A��������� �#���)��x�t��A��*Ŕ4��f��rc�0 �Ǒ�S���v�1�Y9�%��y�D�؍�=��w�}��[����
���2�{[/�)6145��X��s��� ���3L��X��C��uX7c5�{0�g��F!6��X�b�u�)N���)$�ߎ�J~
�X� ��{d�Nv�s��C^ &��r�Du�����
�B�M�(VO�.��a |Z͑V1�*��2u�8 1U��O�ю���xڱ����B�#39(�`�a��Snځ��6�ÿA�~�����Cks���	���(��ذ[2(/�S���VU�B���`��o㈨E��Q���9ь^���� ���H�O��L[t�>�a+p1�" )[��+=�����ͷ�����LU\�D�
&���B,�i��u�	V��e����2e�``K(�fE��0�o��/RW?�@������~��s)�ɽ��o�R�?�z55��^N�4Y9z�zw��7��*��\�_o>|N�[�|h}�@�3o�ģ��h�+8>�ɱ�ྴ��P^(4$ɶ&���P*"7*!.�a��
11�M���o�E�9�����8e{���G�r^Q�lX� e�:�Z��׎���ݘ-�'���J�')��`����z�Ǆ�����O�ipm8r�����	�24S��{�#�O0������}�ftS��&$�Z�V��7��x)�'��B/�'����ۈ�� 8~_ ��� ��{M�l�o�='jOK�2v�CeΓ��oI8��R�t"��T���Aq������ɶ�n;\lۍ$���?�Ir�g1)��ո��j2ގC2����3ۭ�T�6_�n�6g���u�g�ZbM�[E
�w����\����tYy��d�#"�m�խm�P�����<"mm�baÓ$���\�%.��*�r�r�z*�G��ľ�Q�XRH�y�4�Nj`��Z��(��Bn��B*�}��~L ���3����O
v-�<���x��=C�&��ON�W�ѻ�:�G���Q��u���]�WC(B�6���Iꕈ��"c6`�p�\@yc�g|��pF�����
ןn٠�oq�8��w�i��,4�_��;Wf;��pU��B��H�W,G!^�(^��{�v�s# �&7(� WG�$�IJ���Yj��+���ER��(=�I������r�g:h2G� 3J�G���3��j��u,�T���5ih�-��2<FP*x=<�&����̨��F)y�J�O���
�x��նG����&lIW`7����¶���|P���-�]6���������l>f�ќ}����	ݷf�yh�w�'���>���mw�ϝ�4���N�lB�x��'�pu��.t��wޒ��K��������}zc6�֧�7B����D�`l.��h�V�1(u��ߋ����xG��ع*�J��L3V�������$ڇ���,�M���'�	W�{�c1p�O�Ҡʸi'��Y��zs�H�����#'�TXB�V�:m
ݙ[���}q��"���jJ}gm|�!���S*�+��{�h��b�L �w��0��o���q`�`��a5L��y�T�A��9�J5ӧ���Q��ڭa����^�����B�jB�Ռ��R.�PS�H�̎�����")w�T3���d�f��Kepu�g@J�b̒�v��Q�t_����#�5�7p�$x�wuK�F��W���0��V��p���Ut!�LWlӆd��L����ٰ}X]��������^;��d̆��+�2�f�,����@QA!�2q䶁 R���.��E�nY�J��9�tN�Y��;�n�����8v�e��������cQ�� D��0�sk�@�F�P8�ʕ~�,U���NR4�����e=��
���ZG�ʝ�:�m/�n�>��nۇ@%vb~A����a�7g�0O�׽`��HZ�9.����f��+�K
�z��z�2:��<֪�>��oчR�7��� �,��SG�)��?�!���o���@��g,4�Sv&�u�T����g=��ś���T*B��2�\��:�/N#�O��EdfA�=E��z��c���%z�Z*�	�Yv�]���Ok���\^Z��r��:+O>rU_y�0��Ӂ�����lTw��.�=�*ϼz�~sV�#l|Y�<�#͌�bY��(��s�-G�u�"��%�~��+��K2a�#�fS��[pm�_�Z�p��l��D�t�k>�JK��`E�J
�I�"����G|Эy�Yg7hW�?�܌�hca�]�Dr�N�]v���ι)f�т[&���aַU���R�\�M�"���6UxEE��z'��X;�ʀG���:�i7j=��=�� >�x!CU��I��'L�G=�tEMԁ�����Z6ւR[^A�1��G������e�ɓ������ᔎ���3�~wt��a����h���Vl�Rl�7R���z6���J9�}�H.��\�mm7,�U��lWU.g�ݴ�����ե�:g��Rb7D�VC±��x)�h;*v0�>�|�����s�;n���'3i�]��3
º��tʅ2/�H��2z�w��g�O3λ���<x��=
�6�E��������8{�h5�5$f63�����l|�G����h��5�Y�cN]X�*_�"�f�~���	�dj�dl�I'H���s�1��A��y�h�kHH�|��cx����j���f3�� �w������6�BI�%�J�g����Պ���Dܤd	��Gk�?�	�����N�y&UU�����2IT߆%kw��
���1W�������ģo��,�r�U���Ae��:�{�f��n����"�9߻~���p����^|�s��FiȶP. ��`�$�#��pqwX1=�k��� äc��
��ʃή�Y-��8���'�a��U�����}���q8�S���1@#��M�yl,'���2g���b*�ic��
�d<3���s
fީ�8���e����+i��H��k��t��A����Ur���'��fA���g�LK{O�G�Ǭ�H!4D���o��d��iE�_�bpnڨ���5���^�+���ĻX�V��m������&R���l������PJ�g�W�7�H�LCy!F���:���*x��$�Щ��S��%/�t�5�-o�yx���i)�^�/�������8�����RB%4g��(t9rsD%nd�����O��3���#�v�� ��4�社aM�fM X��Z��8���z�#/�uo	����Q}c>�3s�L+�%��K�`��*��k���
���oo�����m{fڋ�	M���	��GWWI��
`��#��+<n�����IW�;r��62 �3�@o�}%��%|��m�E����!�rz�M���tOb��+<�S��G;�L[�G�`b|�f���c0�����Z�m\Z����8�HY����[�;a'a�}}�LT�ȭ �i��L$A�;�5�Gi��k����vH��j��KzmB6)����Ҿh��2�5�">KU�M+>�c QX�6���̎���YB�E~�`��+^�%f���FY�~���J����Q@Y�KܕO��lG�"Y�Cl>�%���H���_���]�9h	_�S�OH��	�e`ƣH�^���-j}�_��qN��$2)6.v��^A4�I�]��%��4����~��k	*<�}��:�v�����Ra�I��=3���6h�-�ax����E1�����A+�k?��t/��Ût��&W��g�IG6�M-3
"�I��(!�q��cOb�~h������doG�U�x�hA�}Ɋ��G��� Y!����z���R=�DPh�a$1a�--��H���އ�@���~�!�Ŋ��&���jQ����d� ڱB��v��\�w���A��Ŕ���[��CL9'�qNv����B���K���؄���[��C�B����F�#�i6�)�K)h��ŏ�����p;���ٯ�W���@@aTp��8�t�ź"��m �D���t�e�h!��0=���`�[�.�0����[_FJ��;e���Ɉ�o���!h��݉�V�JO�� �A2�p��s����P��5�b<�������:�K�`�ǟ�O�=��������"gf����A;zm�_����V��&�Ocɬ���,n���8�.}{Ӆ�T��T#/hz]��mI���	�3����E��|r�E3�x��>��>i��WDG4�+`�/3����V���sc�&�Wf��;�Fm�ƅ��I�Qj��;C����'��QHx��2^�s҂I�tf��D�KBsj8B2��àQK(��ae����
D������"��zf^~��V1�aAP�ǒ,�)�n�ea�Bg�kq50�fH��V�6�X�`�/9�v#B�B��q�0�isr�Ǜ,���%��xe������7E��tg+M��,SL�!�6Z%�I ����b�hc�h)��5���reP����k�$|���|��A��pN��1Y�h�iglER�q����V_?�͇�m�M֠=��П_��_Z�!x��Ǫ�n���h�&��g�fa�T@�)���|�5^�M7(�u��E�O��S���]Bq��Mbpj����?�ĥ��mK�zo=G�Y\���}���͔i�r���l9xnb(�h��WA�L7��4\����i7AnNB�௵�Y.�w�W{�\����v~k ��v����Ǝq��A� ����.���U��c_��!�PץX�ؽ\YR�5!&���؋a%(�W7.��3�?P[T����>�>�[�kӷ3d�������<XH!��W-�H�";�n;�? QY�]�ś���Ս�A��K��u
%�i"!��+��&��\��f(�H���7o�kN���K
�Jf~?)����>4��d�mcb�c"4�>����<`���]ъ-���C��QV�nMP�#'KU�K/�r����'�P�"��;���Ȋa\��ŃoP�8�D��"�ül]2x��@�}�i���S��
�Y��H�	�g�I�H��)x[q(O�dW����vժ��8��r��.f>��Y�"���+>g����0v�0�V/��*�9Z$,&浢��.����g2�}]e=#8y�֍�h9��9�wvQ;\~�yŋ��t�V��fH5�"�9�{:��l��]�i���{ӹ���X���>h��I�{�Tb�� �����I`R%/{�jr�� �~�YҦ	<��j~�R	��D:��u������~"��JۡIleཥ�*�Q8\w~5��2�Ԭ({���%<��i�Jm��r�
�ݽe�;��Xy�2�&�f��bڬ����x&fw��҈�����Czsv�3�Y�2��"���a�%4��(�w�7Nc�$�54�q���5�Mae��c"�@?i/ɕ��7�m��Q�lR�1���E5����r*)������I�>�2�F<gj���ǅ�J5y:
�L����C��S�$�Z�A~�?a�i�E�Rxe)�tL���� �p��Q�"%U�T*S�dxv�/n1PIB�9o^�u���$�)�˿���q,���x �����.����A8-P��$�����~q��S���0�-W�F�d��[��TL�^<L������eUv�Ǖs���27Z#
��3.�	o[���#�s���G�94�T�'.�@���||��tK�"Hub�v���a-f�����^@t'{W0�I �b�N}Z�(�S0���q��ɸj��s�we��7'K6���` <��(��T��f'��Az�A����� i5��y��~�9L_�`'�o��	RF:�g����P0p��n �wL7��V�*�K��������a[z��� ���5X���������a�@/�I�ҩ\�L|!^ ��>�}�3O�����a�������;w��f���}�G�K���t�ې*��tf��:��Q,�y���AB��O_
�m���Hi`R�M����������xb�a!�Y�U�@��pYx�,���.�]{�EӰ9�z��	 ;���K"n܉���HxW�����E�{mC�����?�]{)���	m_ł�砤)��ٹ� �_���X6nsdSR2=��fO?�O�ǯ�� fG@^#Y����.����>�1u��
���E�q[*�,�/̋���8��Rov�n0��+��Al'�P��f�Egl���92��(n�OK�lq����d,˪�ӓhf\���.umd�
��U�q�:t�w�^�� �S�ieKݜ�
S�ӬOܹ��
���Q��z�*Ck̑��
?��0:)�8klS���MH3u+�(F茉��q����FL�қ��tg[xU�Z�&	�J۔K��? �dT>.����-�[��@�OZ�B��6 ���� �F-�W��F��ێ:�A�?��=B���-������[�v@U�k�!~#{Fa��95��a�n�id�@<�*q^�݁���e �$�+^j�h�x	V#_'��7,�z ��fLm����T��kC.q�Y!�R�I�U?��睢 � &�&3&��{"�hS;��_s�>o!V�=�Ei|�N$P�l�dG��Oɵ�Z,q��"���3���\��?���Ϻ��o����QΣ��y�lN�,5j%P�މ 
�>�����1+��Ƀ�^�����]��x��d ����ڧd���lU#A�ɕ��%�E�f�����������FΈZ�|�]��gO"�4` b������J�v5Q�>��&q&�ΏgIA�R/�s�VXOt4����+	X�5F�d]�5�Ùi�k�������KW��
)u��H�or�8_���gR��$#?&fKy֙	Ne�Rh�c`I�'c{q~�tWT)@!�$Q�Q�(�ײi4��W^M)Q*�'�[8�\X���Ix��l�h���N��.���ʳg�(���dO
g�iI���*��S1id��\ƪu�Ꮢ�Ű�N��}�X�P��T����<��j���߉}�e�B�$ͼgf����`rC���]���ɋd��D��i�����]��:I��2�|��H�jm���n�5�I+ǁ8Q��1V�e��B�̐m�I
K�}ϮpS0P�0�r}AJr�-�L_�p�Ε���}�~mm7s�#r�]�
�@�?���n.����Ծ4Ӳ1��Ι6�mqC��؃y��=]$�Rw�4�׆�H�קL�kUƿ�������Z�n��^��� MmL@|��F*�/́�~�hh�y�����݊@a&��!�� ,s���Ӟ)�el�u����	�2�;*��ܑ�-i��� ��͆ܩ��;e�gn,��*Y]4G,��]�ۚ��n��o�EJ�as�$b�B�'m�Hf�0��|�P2�y�y3��kL��� � <y��4�
�w�1��R��r+s���D-\{�z \�$?�-t��&s�.d����K'�=����'���%N�Y��|�礗�ʆ������z!+���0�督�c�&��O�|!>}�H�uO�p"I�B�)MG$��LE�<�6M�\\��f�����T���׀BV+�x"���q�a?���uX(��J�߅�Z�B�UeH�4`fhr�#M�SXQ�����"��Yֺ����YA�rdZ����R*L#�E��t��tӽY=�FB|c2V��uR�]b��Ư\��,�Ӳp��`�ٝUy4�	˛P��(e �E���Ez٭B��%H�4����uNxo~���(�^�:%��푧<@h��]����T�e�;��߫ ��mD������u
^�:��ٝ㛷��3GI<����M��,_N�><��$�=�;��x���kb���ZqD��S�O��'�´Z�L���#+�o�V�ւ�t�9��q5��Z�˲�U�d��*�0����F$��/tR�5W&�1������biE�c"�*���Ɛ=��=�����|��� �d#�b��r�����������0�Sj���]��T$B�Y���4L��
t(���UG%�٨.៵�E�j�8܏�X��R� G]AM��1���kNI���i�^kA&���?�Э����ϼ�5�N�p�,#p�7k��]�0�$�u��i�RkwId�K
&�a��һ�*���o3�[��1�q�+�Q�o�ߤ��j�ƿ�`���B	��Ǆ}���S#d�6?X�sGtD�7��6�
0���3�|�X�g��@���D��\�w#���oI�Ǽn�����l��V��P�l�����Nr+V+rHD��"�����ۯ�_��z��IFe��5rY/"Ԃ��'뀠;�_�#�E�C6�~�N�&�� �l�!D�ߚ��V�[��[�L��t�$rYqf�18�r�|V���ʡ�$��Aĳ���pV�*�d��5�{�~����b��G�1gg�usv�9	{��l��R��C �Yeb�`#7��<[���v���a�l�ʸr��"e����d��!�
s�;���F98��t�+	mv������s�J{��Fd$-��Z��[�8� ��Xǀ��3����u�û�8Ԗ�G���<"A+�<�էA#˭�>�2�2���P8<��&���Á��H�\#_����u���z�:��算cvd�8�V'm �h�����^����Az���|�2�<��M���s4�4�Z����0ф!����R@���N{qJ%'R���**e�ũ<x��A��Հ��!0�ȗV���N���*,����=�E��UV*����eD,�������`anĵ��>�[�_mW�s�������]I4IG-(M!dPGkv�t�>�\�AN��X�e��>��l�c�K�,���A��иg�ٯ��/<;��f6%w��:z�'r(��a1x�B�0��nq�\R�\�c6���0�ufC�_��VvL�q�Α폑�7;~����MO=I�|�8��v�=�k�C7Z}$ɸ	8�*!){(��-�����?.rl;?�T5B����������}NV��Z�n	$fz���hg������K\pv�wGr��hjMY���<� ��w���6�I�o�Y�.e�w�ԇ��gQ��c� o��Wx�q�3U���v<����gR���B�ʷ�Z�N|��
� R��G1��o����jYFħ�7r6��O������1�|�9S�*�������d*]�u�s!X���ўx%�ui�<���+�|t7.G�r��:�qG=���9������4>���7��~N��'��Xm���{����_�n���GKh�-UI��d�����<t�X^�N>N|,,6v�H,����?��H_r1w�����;�\h�%m
�9��8g|��� ]���W� ����+����;6,�j�+H�Q#n=$D\��1�N���2�$�%�=~��z~�k�qш�N�	�]���f�`��������r��JcϨsZ��Q��4e�FÎd�0>��f	� Ֆ^���f�ʱ-,}��ZTf"պ.q�;`+`�T��?;���hl�%.�m���ӈ�q�����j�b`��J?n������ʹV[DA��g�ү�I��3h���\79;�T��y��%D(�}oO����#V��e����+5i>�����ѕ�<D���B�i�qn���^���v�joӿ�@A�34�I��1��5��JNG�k���$I���u���xe�K�ӁI~W�-�,S#|��?���A�z$ca����
�e\����$Ea	�<�;�^�䕪��cl����i�)�����p*�1� 5����&Cym�� ,,�c��W� �t�XL8�I���*��؁*�u�<K���ԩkD��d�p�	�9��c�%���%)>�����Ķ�'�b�w#�aӌ?ˋ��  ����sRz��c�!սQC,�H���g��v�IkK���u[�А*}��c�5�ڔ)������sb�݁t�/���ЗQ� �y�b�������s��\ ��X�K��4]�&#��Lӣ.����WCNc��޴����B�0���M��	�Y�bD��vY)n��Z`=M��Z�� x��8�?=�j&&�1h��_����9����ה�,�m����!TG�R�6��$<�'Nk@w2i�9Q��u�C�	����?$�2�y�0ބ��gY�N%e[i Z8༅��a[k������.�Ά�[s����(�)���H��Qm�D��˝���2��:WKXx�Ϭ"���pt��i�$J�s��c�Y�~�5�$�7a$�.6ٚ�Ӓ�]�?L��܁$������G�,��>/}�z��5 g�v���MZ�7� 5ب��
�>���5��0D �-�Dg�3���a%p8����$�Hב�Ki'�jV���"^쑀9�WP�㼏����Y���f͸��+��@�Y��c'<�o[	�������j�������dI@Y�v(k��eX�Np.Xiz�5!�A���:u�u[-h24l�#�3dZj�f����e�	�o����	JA�:ܭJ�����KX�Vԁ�����;�̾>�|4��u�sNJ�/RwDa�8z���HV1x\.��!Hf��Ob�5Ϟ_&�
���m3�WJ��L&��sD-Y�?8�LP1Z��vC����F�x��m-�	.w*�2Oކo���U�O��y�T���(�@�\�T��������W{���o��L XE�£Bn�.7HA���qk8��I�y`��2�[OC���r��͎�Gի	�Tg����\TO6�w77H����!@D(h{�b�dZЙ%b����f91%��6xC�qזEQ��9�k�a���fə����7j�(�M��/�9NY�/��r��C(d&n��x]�L-#7�����΋��&�O/�ho�*�t�rf�lWC(�=���p����@U沖��=��(�F��+��e��N3�#o�FvEL�1¼��|���㯭��KꛫW��{#''	��r=�Kkz��s�c�+�TL��ך��D�!t�����*�gI�ǢFӘ_�����/~����;_4�ZOBkh�v�X��1e#I�7U�fq�8e}��k���X,�%ٙFK��3��f(O�� �OJ�p~w��Mد
y�b����J},(�U��)ST6h���N���Qz��\����Bz���5��rs5�?����0��� ����:��"]Z$b�Qy��fC���*Q��w�02���y ��;�yI������ˆ��y?b�{)&CLv<b���_e��Om|K��M�o��i�����d�N�:����Ⱦ������WH*��K�I�Ɂ7�;�9/�2���X����Z^ h�ܩ.M���E�{��-�䄛b�U�]5�
ix��P]P^�|��͜6@�����:0��I������X��:^Gk���.=�Pn�(Y��j";������gv:ܥOB�/���\�1�
_u�B�i@-����Ў%�?�, ��>�'��Փ[��C#�J�n6�ԡ��x{c��V�y�7�,��?p�t�Ÿ��l]�]����);e�&dnk�ee��-l�(�~��/�*�c�ʄ��7#��Qh����0�*�"���|PUм������}�%?Z<[���CB��I�L��s��\�DSL7���~LI�y ���p��y0�ż�ea�:.��b��C_G 	S��K@�t��9�O:9�q�׆���D���,�������,�V��H��&�>3�EK�4��Uk���/�1H��0=������b�1�m���M��|7��1�v2�l�HoՊ
>IO<x�e�Vw=P�$�Ar'㝓M^�P�%�f���Y���W����$x�;�{u�f�B�.���Y�1J���4�~={a��X�Qj��Ş�х%�)��b��` �-�"όT��zSq ~���q��r����WUrn��.�ȼ��h��W_�cx�${��
Pd��@�6W��mR7,�s�"�o�5��1g�]� �I��+��A��-;ܕU�%#��⨘��k�~�-����(ݔ��q3Y�ĝ�㋝ֈ<�eC9��x�dMOĎ�ԘJ��y����V�H�~Dԧ(w��?>����C峴Q]"V�Hv�E�(�@�O$�[��h�'�"�8_�3-���{������Hc�tU��T6�?#�<BtB�ܽ��x��Q�SkLT���!�W���uX��1@�͕�rJ�K��Z��Sr�f��`��Gy��e>yv2��6�ֱ���	�EN�����:ʚ��@O)�"�<�
1Ѝ��:��=�+��x���7S��(��w�,	�eB������&[��τ�ߏ�$�����@H���b��OS
�t�;�=y��L��nU�����؅�IJx��(�Wvxe1��pb���_�o�tw���p�"�v���7�eL_�(�j�(��c�`4(���l� ���&T�G�ϵ�N�na䑔���s[��5)�Ny
 & ��?G q�C3[�_�E[�@b�����VN:�a8;?J�t����<UVA�٣��ZJ�y����~��P"w������8��G7�77�u8��G��7���>FWI*Q���qT�`���Ru��w�.�%����L9��-��sQ���e_v��g\Q��[��8[d�6H��E(�/��b*P�h��_�k�r�T#�t�@3���A�I�~	��F��{�UG'p���㒗j�j|��DX�W��,,rG+*���=a�,g*��^%0k0u��ݼ\�KD	"�4�R<�(G�����{��
���wdTFQ�ަ�/á�2�k�ie��D��~b��پ��	�Hˮ�H���^a,�ok��QZe�;r���HM�,r(���"����Wu��~�F���񬰦I��=ز�	�N��=�3Ɏ�� �,��*g+*��� �X������Z^���?!D���N�g�x���LF��6d8���dÿ��m�>?`b@�hX�f�o��q���f�,�;G�����ǉ>�Q�jɺ�1����V�p�4��^�Qۡ�EUK&]��u=� �O4A ��7ꚫ4���P��N�T܃n჏�]�E$�G��ΐY�h���2��P�Q&!a7DPb0����n����FqO���GC�[c��${�Y?y��b�d³�3�?9���.��*r�X�(9�k�u����%5�8��C�}|�iе�5�7�y���{6G�c3ީ��!��'����Q{s hv��^�s�������t/#K.Ř�~��Q�=�ϙXz�OKe>Ѧ���q'`��(��q��P3O����H��)�8=��9�쟐�����&���9h �}�b���'��ɓZ��c0��7���5&����a�^�L��8C�q�\��-o���¢;�%�6���H'��޷hE������u5� �5U��X�q}YXR�+�:LpG����|�L}����*���5[�E@�Y�ޱ9_�\ ������`�ٜ�'�)�����,�C���p��M�#'�����)~"��b�»"@��>`��Lk��w��Q\2����^_�IP��0k�V0����Z7N��ܘީ� 	0�햺�=�V3а��z>���+�q
 .�:~;��^�hI?I��R���L�]�Z��	�L���?B�>ҾF�
��3��:�LgEto�J�^N�Q�w�(2��ڼ�Gi��S���m�&���:��y�@���f}���x>&���ishl >Q�p?�}oL���_d��Ò�����έ��ؐn����R�N:˃��%cx��ܓxt�c��3�g�$O�[E{���b�g�W�|�`1�=^�����s��M ��d��f�����-W��1��> ��W@���ۏ��OkK٣�9�����í��Du�l)���%�SU���Q��
u "�sU�x�}3CH7t��7��I~�-��_��.u�Mo~{�.�$0" S��3Ϋ-�d�A"���ĳ�K����^c�vz�'�����<�{۟_���LЖ�Jsf9�4�t�}�E��֕���{(�BS����#x0���{���r��a4�֤tv�&~9��G��(A@�SBt��xBi:��d$-��*DΌV�i��u���Dɓ*a���ەR������IBd)��d�����Rk��������*ƕh��<�@y�a�8�88�G� �o�g��?�o(s
t۔0��7�5��L}1�D���f(�H������{
w�L������TS�Q�9k9�	֮
��C��\s��١�
����H�G�ca'�W�7X�Ŗ�3���������ZH0�w�n0ZU[�(�
���$T?�hV���Y򶹋��O�{�P��+ΰ�'D��S�� w�Cj�Xv�/��3�����<�ܖ�}M��cl������8���j#�`��j�Ց�W���K>d�U����wi���F-��%�����+���r���*Ag�h�_��6�Y8�	M�_���M!�l
�0�A����YuP�����)?1 �ρJ�6�����E`�{k0v:k�K��mQ3ohK9?�AT��-7g��ҏ	y���vo����VЁK;n��$����E{|h�{���Y\YJ#�c�{�T� ����"���C'��c)�C:��K^�q�0��7[���>=���g����6���l�����90�����4�yW{A��+yV�ў���O��')GȢD��W��(���>n����N^&υ�.Dj?ߥˆd�&�(�`漅2��X�DƑ��y=zٟ�п���|2v�Y�D���ˍ� $�?����׋yEJ׺���b�����n{߉D#O7�%����)6�'t)�,�h(�O���}�ߎ���.%�;D�|�P��0z؛aa��őhw��w��)^��H�Q�NC˘(�%�������x�BL	���h۩"�#��;�:?�Ys��\=��S�����&�S#�YH�T>�|��K�L�e��C{7�=f�E�x�B�[�6M?t��_�1r�ʰ[ou��8���/ѝe�3�}&ka�Nq��+&P~s�BD�[&l�~�oHO���(�C�+��-�ss1-�q%�6o�g�㳭`�l���/�}�
�u�:}��v�}D��k�v��H�i�p�^���~=��PWjW��{�|W<��`Eq�;y��2����r����ٍ�ƾ�q��t�S�S�d4y�v�@�oC PpF���?��.8sw�a��=Qb]�$ƪ;�ȏTf��kc���^D��#�ם/.�t�Ϡ�<��w{>o�n�%���rr��d���N��}�3���̝;謮l.X��T	P��i,�l9~�xب8���Ƭ)�'�4����p*��1ZFt���G��l&4k)I���F�%T��A.�����WkVe?������gwv��4���Vx���1a��lW,KkS	;�j~�)��r��=��\�b	�.
U����.��B��^FO]��C^:�ʍ�+NH#<�K�{[0������qV6�-��c��%�Օ^��^�3�쮋���f�]��d����liU��N#%��6O�@ۛ;G%��O�$�(���-��l�k�#n|c|�s�̕��A�f���Dc���/vRr|�CUV��}�
�hI���J��p\������zV�8,�(��b0�QTr�[Cj�,�vA]�ȯFN�<�ʀNڮ�W�s��X�3W�}VI���:��va�wȍJn|��ܰ��.]�P�����������Ck��6�:��_�1D�����}���OlE�ŕ�6����d��-P����ܐ��P'���fi��jȦ<��O�,)i�ީ��Ζ����#�Gp�b�E���j��a��ۓ�U���Iy��]y�~Q8Ֆ��9��V]�!!�/�`i�>�ȉ���f~�Ή���jݒ��%��{�8Eoyߠ���Q��V_t4�e2%`k�������i>�(Z�ܸ�p(>�?�T�KC1[| d���[��0�C~�����E�cPu�2l��cH>?�/aJ�v�.��"%T\\��Y�P����ӄ6�~�k:߻B��c�M,��u�ՈՏǲV��ua��ʻ�{i'+ځ1��N����.px��:h�y���ao�<ؤ�U �D���ڗ$�<��b��?��Ls\���/Έ���?+5�IyޗQR�
�0L7�V���s�s�"��$�*;�&�J�6gKn���j|։��w먱ar��[ҍl����Z��!�\��@V���ܻ��{ϝ�"����/B���s����cl��dn.xn{��<��#]U�jr�������#�T�pҬ���u��E�F�,f�l��k����@U�oFM�X�żX�}��.��`d�6m?�i��є_��vOt����44���s;�J+��<��.��b�����/���T2_�:�D.X)�9�%1����q�lW;��EtݪNf��V�hp��V��>A�Q�/B7==^��@�<�ǲʳ���/���Z��/���k󕂵݇��{J*ѱm�q2ȟD�(�J���������la����&f7���۷i�Q)��44����	��4���4�O5Cз�����q�[6T���u�#�1��9���'j��-N��o;u��B�AP�?ק�^��_�l��9��O )Ʋ��ҽX�Pi��~�h����ӆu��lj�B��L�d8�� P���=ϋ����GIE	1Zg9_���ͤ�}�s�W�_fh� e��B+�Xఒj=|@"O�Y�~�����,ZV�2l�=a)�?�9���-D�R��EYF��_
L|!����{J� �]x�&.�ktj0,�������o-�mR ��ueĦ���
y<Njg�"s�Z�N�\�l�s�%�1�QB�ja��;5�?͑~���P�'�$��ƨ:;(�T���D�Eы��L�=+	B�����@-�Š�*��A[}l���o��֒['�#��M!�s���{��ӵ	�&��5�I1"��y��3E��'�_��$9�g�A���)�L	]A�iY�2����"���
22����� '���\~���YwT��0搣��(4;�Z�.���uvd��z��{�ML������έ���L(RB��X'l�����!U��� q�@����GZ��`��P%�[@��(X�;={W��K���F��!��H��/O`��;�e�E����	�TL����B%��)�F�t��� 
�f��_�*_	ߊO$I�@�"��꣩��hgJVb4�X�>_DW��B{.�r����-���뽗G������SW~Ři�"�\���u�Ρ2O[Tr@�����U�aPBh/
t|3x���k��26 �c+3�UȖa� �0W�噇z:ݾVOU|Bf�չ�Nz���
s8������;�N9Af|�!N� $b���hqju !��-Xl���5������N���,FA�;��O�1�ͷ�3B}d�\Y�M呢��Y�s}E�^�X!���L�Tm��������֝���j�_jP�a4��T@��Yq��������i��n��y�h��j��U;�i<����jჶ+�ID}v����)�H�.C�1#��*�[�
��G4���"}�e#J7�+�:x�^�PG�P�(��o�%}Ǭy?"_�����[\QN�u��h�̡���G#���e-?����iZ�����U�l"��+�.ɶyzB@�(��V(g�ʤ���rW�|:Oc�ߞ7�H�q�
�o�$빾]4��r*�H�w��DVwc59ff����60kĞ�K^���E�)o?A#��Z��XT��? �,��7��8RK>|�=᪁g�fk�s^T�7"T��OB�.�4Z�cwʚ\7���<��H��+i�W�bd2P�޸����Uw��/4�b���ߨ�@����d�Gm*c�e�;�@��=�vE/�U�;A�kT�˗ߚc:�ĵ����p��1�L���W:�X���EE1�.��c��n?��.��9���
#iX��8� �/�";�n0~Qx*��ٮ7+��`��4C����a�/�O�b; �;!��,�H�[��!3�`��7�M�)`s�3l��<^���x���8��&�x�H���$�g-_"�J�����%}��@�� I��a�	f�ZW������F�k���v^�9��J�P[21��Wu���GZf0,��y9٤������o��w��<�7z1bd�n�d�F7��s���})nL��su��lRL�����qu�ﶀ��z�+8f>����Z�.��j�2�D����8����6��*6���{8�T �~�uQ	_)~�8V��lG-���3�_�(��D����n<��I�f�%dRa�[7�	ӈ��ju^� vf��/�Y�@4I���w��F,��&�:��R/��ڑ���z�P�z3���QDA��12��1id^0���D�C�{�Θ�J�K���N��Va8G�5�<� $u�]M�����`�?0�$X/ ��h���L\��l!;̞�}��ʧ�Po;�9��US�Zgz�EO�1�r x]B���n��A�֟i�*���G(W�x��<�y�n~vFrw���wY�*Z��!�$�C��̖�������d?j
������yH�EH	�ޓ(Ķ��A�ʵ����1���7#r�꿎����=��Y��r�Z�㵦�8��%n�/�Ϩ��+�E� ����چmm��>��B&c�zW���{�����֐��Q��4�R}Z� �C�ݨ�|���+)G��1�O^�pQ���neBH��~��K��,��+Tj['z�<^��R"��˧f��O�ݏQ�i�ћ=r2֞Iф�z���tŎ�ʣ,fw8��̵��B׻����Ⱥ����ę�aN[��@jl<��r��:��P�0��eҙA�$����m4��ǡg���Z����tI͒ ���N�E�<kSwP�	f�HoL��Rd#S��(_=!!�f"�@�� �����Cd�TV���VE�U5��������"LM�>D!��r�	!ޯ[�+��
�L�rw�(}���Ι�Z�b9�|0�mR[�ǪI��.�����V��[��p8��swa �^V�����qkJӨհ�A���	k#���3`)AV�����!"EK�EpP؍k��h�5���6z�w�x�3�8;)���߬�Tb�
�j��D	{{�ծ pu42hʰ��h��7���F�T�s�⦹���݋�;����tZ�D�y$�E����^������8a��ɾ�ez�_��w�NS
DZ-�B�J#e�a¬*:��a렣�?
��{c�_�'����jrzA
���8u�庴M�G+B� WXO�_�i]n+/A���dA����K?�H����ҽ)���z�K��x�ԐOES]�V��b�й�1_�.hth`"U�`�$�fFyc�+;��*��������XW.��Wb���ק�;+vG���	��j����=ʧ�]�@jpq9�I`0��Q B�9�у�d���4#(8��޺�z�:A��w��f6��r�x��%y~{:&Qw���j kq�H�����EF�#w����0�9�^�X��P�
���c������`X�-���7������](�o�w�Y��nKN�A8K􁡒�ů!ĺ�E��V�v�J$M��4��Q�m�y�R��!B�	��M�x8� ^~>-&�<K���I���tֈX?�����F%A���v��9��������TH���BN�u�#R�TK�	N���!� ���S�{��_���KD�iX_�>:Jw(J��(��2��I��b�
�)���!ԔP[d��5a3?WV:�˰����Ӂ��i�?b6Dw�S��M�򼻡8����վ���g6�~��;R�6Y�����Ȅ�T��݊YP`j��@�W�w�l��'�I<5���)+�yK5#ز����&( ݚ�DȨ��Ǯ3u���Y�YL��?ɥe�8º���# @��u���G�����}?��"�����K~Q����?�
WpBlZ�ߊ|K�� �q�PZ"�^�����6��-G�GAP��p��ڍ.���O��z> ���;�����(s:6#�P�onJ�Z���9��#��_�*�޼J�|0(+��Iċ�_\�'zgG=��V�<q�G�!�Ž^ Dr�F���Je��uߩ�V.����θ:�Ͱ�t�����/8��S�]N�޾l�ٞ>�<�un���Mg�X��k~pJQ��\��~T��f��(@��`}�590�b9� ��/QPz���4�;�����k�b�p��L��_�EBy<�X�(��,li�W�������;���0WU��O@b㳃Z|ud�j�ZȽ1�k5�д����U�6$>�T��c�4�&cf�����
��A^^��\�'$Y4�G�Lی�	)#MW��Q������� �>��w��aB�z�l3)ZE�h���ب�2��[>O���;}n�%"V��dM���G�]DD���5���kkj{w�A)ڰKS�F��X�S&'��!v<.������WW���T��]x�LT�l rċ�A_�����&�DKc�I"��:�����Xd��	|)e\!U]�����:o���aVC!\�^��K ׺��g�X!R?�p���Tظ���,m�� �|D� �\���1��W���B�Bo�h�=~6��-���;8�f_n��E�;X���i	%��{��Tif���zN��tg,6k:�OIϮ���>�"I� I�0�xF���_�]�+�WB;b��Q4Y�T9��Vh�D�BS�0$��?I)i����[/�Wn'�%�/��r�Ξx���g*tg��{�48ga�k�[j�<����B}짤����b,��=bb�:�D;���G�G�7���p�}�̪,�<�
����� {1�b��9k	����I$O�sg<a)v��"1~ ���(�p�/q�Y�d��>{� ��D#'�F���}L������UK#�i�PZ��S�D�N7哷�Z���G���Gt��+�I���V���gC�.|m��}�Ly!��==�q�����Wed�L*/z��V����c[RE��U�"�=�L�i�T?A�˟��Ǘ��l%��ms�m��Bg��V�~��C�� �!�y��R]�KF�/`1�N�ȕ�!�TtY�_����Z�sY�c��l���ոl=\�x/�Ud�+t?T�P2Ѩp�Ms��5���6L�	_� lR��j�F>�9��Oe#?˾j%9b���.�9dnJ!����PF�?t�P�u���E��Pn8��ͼ���呵�B��xe�ّ�z�1[I�1ۼ�[��lOH7�"����	ksx��j5�O,"n�_��X�D���ظ�$b=6�G%bթf��]�w�7����ͱ��ʩ�ݠD��u,�Hi"����!s��t?s��������l�M��#���V�2�K�v�ЭA�m�t�c�6������)���C��ff�O2�R��y��e�awa%K&Z��7$����]��	J�	��z3H�0V&q����*uf�͂����T� r܂&�u$ѷ X]���� ��(��-�Y��#ZheM��H���(��c�V<�L`Zf�$���ȴ����B��~�$����;hoY�`{��$wz��2,,�K_z����B���cۼ,�b�	�ٟY�gN�&G,�o�|��1K�ևeTg����95���/���=�J�����T���M�e81i��{Y�����uN׉����N�9g!����q}�0��;<Ej@:�����`�Y�v�}��A�f_��6�~T,R�spF�t(+�0�([���(�-�S�I|���a+��l��;r�2,�_�������O�� �c|XM�ps�sVS��&f����2KGȆ��Z���֬��ҿ�K��g�:tB�0ZW�9�tѓ��h���ƥ���7eY� ?��>��7��K�1��廗e��]��@�P��Ŝ��Z�>�At*��[b�;��?��W�%��"���n.Q�B|G��h޿/�7Sz��|&��h��~`��U/��yr]-|H꣹[�����eWA`\CM��4�����h�L�f�:�'%��An�'ܫ��`O��Ĺ���Gq�D�-0��i+�o
*�����a���~B⑵=6Ռ�Gb��ĦrE?B$��?���*�rO(�&��<7���x��;,�H�ա$��Wy�E}�k!���� ���9Sc ���<�E�D �y�l7�E�Qm W_���J}S�*�K0V���݅�Q�F	�If�r	�C	�С"�j��B@�LY�b�����>I 	P�qe �.�>���7z���D���م�R���d��*s�c�76�FH�$��U��z��1���X��Μ��v���TW/��PЃ�=;���4�����Ϲ.�O'oq��;^�3._�B�"�H�m����p[b�4��xMwd-\������\?A�3@�u����R�c�+�ۻ�!��=��7����>��3�R�Uˊ�tWTa�@\�
�m-��g�uF!�l��Q�YH����+���%���O]㹇[r}��U���w��]:�&�^-���ֲF��NU�q��X�ޖ0�����c��*��k�Kk���ְq��^��E����C��%�1�6j|�t���n���#{چu�%@<�L�,7z�r����2�i2-�O��o�s��3�m.� wX�R0b߆HǬ��	���[�F4�K�6d�����M:^
B2&�=;u �*խ�������P�d��H}n��!.AlM9�����4��2��V��3��������!l�3������bmI�<�쫢�M��ʞ�]%B������X�i�#��I&Y��XR�Y='d��r�Bj��C�H��(�i;��*�d3�d2�ڼ=T�d��l�rL@fj�u����m�ۢ��� B�'d:�Adr�N��]�OW�T�ckC�+�9�K���u�����,�����!���٨i��<Z���Ė���FTk�A��~n�a-��d����C��e��-�0��z�4\�E�FVL֋�F�龨v�c��'�Rj�L�"]�Zm+�c�MB�Dl3���ȩ.��u�|v�)����e)�x��o�&.m���3�z =ͰSn�e��-�_8���×�2R��no㙦Ǌ�f�}��F����1��<����\���b�ձ:� b�Z`"7
�[�����ޚ�̾R߼�ڰv,gr,`-���ɠ��Є�Wњ\Z�7Q�MĊ���!��&&�	q^��_�j�ļ����ue[ݴ"�kSB�<���'X���U�5�?���L5�`J�̴�U5+7��hȂi�䵃��5ǃ�}�q��(-��pWL�s�a���H��ӛ�P�����J����b��B����;-�U�3�+JU1�]ۘ���ڢ��'藁���H,�Z�gFҤ'd��\V|�u�g+��:ў��+gx9D�� ы�l���� 8�V��E�D���K��O�uڧb�Έ��������O$�}�ߗ�ļu�G/J<�j��Ģ��Z��賊Aґ�vG������q\륦LX3)`���Y�pJ��+�n(WN�<�H*���O���{G8��6Q^9U�jy�9x��7�N]ܒ��Ƅ�[�uT���<O���T�G��eٟ}���( �{@���N ����i��ђS��}���`�����O"�Ip��Œh��j�,ʆ#4�9�nȋ�쮡�O?j4��A��7����Ўj�����9�h3)�d�,�j�Q�H́4�u���[��{��,��=��Ғ�?������)N���/��:�M��.ድ%l5S�Q�̭{2Ҋ���Bs���<)1��UV�Gyû���CN5>����D���|�x�>�l6�l�b�Oe�����0�2(��4���YM���v��O"L�}>���x�B"�XUN6}�G�J�n;� �8���CFB���DP+�;�� �mñGm�Wc�c�ZWT�D��֩U@@�W� �����m_E;�D�`�1���Ƭ릲Jt���Y�o�YBdE ��h���N3a�ĀJD����@���&΢m2!}]����;�2�9
*@^�C�� ��ˤ7+��ލ	f"0�_ㄗ�Puiv��RY��h|�J� �X�`�v�·Q���m��g��%�y��Y���O'(t�MFB�N�qY�h1������wc��w���K��u�B�ƃ���XN�l.��CS��4�5=��pV�mA=�\$��:�̔B~a']�ͨ&Q�B5�&��8z����"�/b�YZ��
�0�m��lZ�OY�a&���F�A	�`�mu��d��|nc޳W��,�|�̝�

�䍗�Y�S���|| 0B��-���k_�-��kNB�ɽ�-�=A�����6���5^����YѪ뱑�k�����,�f^S���q�SWP�Ũ�
!��ٱ*��W+����W�^�H��c����to���&�N���1秤�|���jۨj�l�Ӣ�c��fəQu�;}E�'cjP��r'�&���(O��W��g��nAI����)6@M���K��P�ξ������E�wYΪ�&��M�#u�*40<҃��e�ip���*�����Ô:e�����,� $�o7�$���^y�$V��y�@�*�����9��D�Q}��mG |��*��T|�UJ{(�{��ӄْ;=FTh����W. ��J���Ե#|�.r�a��#�x�}qxqҦ�IA�Ď��ඓ+��[5��,�����d��Z���jR=Fh���YlK��X��n��r|�=�aŞV:	�t��U{[7˵p��;^,�q|�DHvny�A������0��o0+��v�.'��'I�׌�]L*�_��Y�0��X�dߖ���H6y�?vAO�4}�P��)��U��ˡp(�w�s|��P1�%f�CL�c1�7��P$�%�P������C:^�C�`)��f�|k�<�S�aK�����5�6k���/*rX�M�D���C�3��
�(��;��V�[�p�S���i�Ǥ�T�2�q7�m�y�"�լ�uf���	�g���8
:.��Uӗ�i��SlG�m	�H�Ռ�87�Cla��m�a��P�ʣbz����o�g=��g͈^h���kk��$ƾ�]I���5[��
.?�� �p~H�.��bl�4vi�&9וێa�
'�ގ��^��+�c��Y��W���9g;�L܌P���Ȯb
yO5���8��i�U��NC(2A*(�;g��B6�-��|�ޣ���"0�Y�C��~V~� ~�'ng�gd�gmԯ�%㮖��1M�u�y��n硐���ޚ��r"_ͳ��.��u��<��PG���d.�ί�P��J�uy Ҙ!��L��xH����]kA"ޓ��9��<��2���so��El�T��1��=�5����t�S�
�;��M�ӵw�7���3�iy���/o��E�#����yHN�C輠?��!{��'<i������o�N]�'Rm㭥��Lu[�!{�o�̴���CD�x}X���i��V���eIg�d}=v��Q,�P@�ݫ���^�d<��6h���
�
�[P�SO�c�F��d�0��Ev-�����,x�BF=�Ng&vdB��FY0:T�.a��,�h��)��w���C�Z3;�Kx���J j���B�1���ֻKk�Z������Y
��v{v�3���l����$�wu�y�A���|�"�2ش�� �5�p�����ϧf9F9�nyɌ��^%d�d�γ]W;���Ӥ�a�c�tUT*<2u7 �\�h�*�p�~������"�ua�����ҥ�,��cF��Z��=m,^_��Q��3�+�y�c&�]�J0[� C���cG!t��%�|�#s8�v��^۸�	.�_�_bٳa?�N$�=���j�}Zs9%���h$��tWK�^�lH{�*��m
K��?�����ꨉS^9�����F�*4v�ݦ�-�tr�Z8;r�jl�.����G��h��q��λ�W�S���jZ�wnx������xB���<
,ygҴ�w>�6:���bL�?Rl�,;�M"����\:s�F���Kb^���F^�.�y������ �l?O��7ӌ���ۧv��V���B+j8&��_��Pb��x$Z��=��v���M%޴dg����/':R4q�j��[=��X�@̏1��&js�o��"ޕ�T��m�����b�We��ȶ���&�<���dh�
�����n����l�����7�E���3@�u���nD^f��;���E��R�ٜ�e����I�X���7��2`��g��dݨ͖�z�ɷ밄��m�`�]Ȋ�̃;#����vF#�R����r�IwGHNt�!���@8@�#-����:I�k�gS�a�OԛrF�d�H�8.�
�Y�bq��'���O��1�
g�Jm��� �SQ�<�$�3��#^&���ޑ/����^����k�I�'�7b $�4�@�%��'	R�Ra�(��޵�8�֞c߽l�yO���KmuNƫ�%@˳��\3�����Oe	u2Ԓ�������XH�B�
��+⁞��y���҄uT���x����Hq�)1�@��0��	�}w��w���m`g�6Ӣ~�m3c�"k^�C(�^FO��<ǫ��Sg�9k>]�d+������E��ê辑�M�K��2���/�!<W���	����+����ږA]q)W5�~i��Y�C�N�U��)�rʆH�%kG�\a��*�Kj�%"��µWM$�~�C3�L�ڴ��>�z'Y�nZE���@�g�D���q��/^oƲ�x���N{�&��
=՛��q�����ؖC�<��l��W�U��18m�y�ޫ�f�ե�˿�e��H��ږ��sY\�ؔ�'��u$%`��xK:b<�G�"EM��㹒��O3i7�8k�Kq��Jɏ6�0V��.p8"ܪ��ߋ,�Ft�V&B�_1����� ��ꥮ�k��*d��ؤ?f�2*fț��5��	��0�E��ygk�`��ch�#�n⓮���2a=3üg��U��?:VE@�Ъ�T�?7�b��Dԏc�%���,sL�1�3���sI���V�'��=5�>�!Kw�6��C=�DLN��q0�zs���#f���|��ҵ�(�l瑬֠�I[�xK$�8)�L���;�jI�ƨmz�m ��������S����t����K��=�Y�KY�3�E�Х!
k_!u$_�q�	#(�f�P;2+�K�������o��æ���^i��$Ns�q) Nw���hQ�6���a0n�*L9W��^��(w߽.~+���\5`>�)2�޴�5=�L��l��ADǖ���Q�c�D�jw������+5������]�=�93j�?�/�]M'�`��dy�<Մ4��E��c0�C8`~�W�{�����X��bn�{=Ԫ��{�/���i�Q��	i�����	]�	p��J�.����wf�5�`���E�!�:��@����W�Pa���ф�<^�r������71bv�����k$N���P�-�Y�P��`@�]�a<̼�՞�և�U5���q����~ue�$k����£x�i�	
pW�l��J|��)�&�3�jYO�c�͸]����.l$��B�\��JZ�����آn�_�WB�\ϲ�����l�Q�%9}�;��Wa^$�:�|�#�n��DB�?^�r�|���Z��vٟ�GB���/:���Q)����\�ôz����%�d�?l���N��ٹH��=��r��I�vc?
��f�ْ���O)U�)}�XfJ�S��٩笄v�k��(�y�B�>q��qg�-��>N?W�u��=���4S�&--�����_4̾��Ľn[RP�P.6��)�������������MN��n��	GNg�dm��2h5�?��RC~<F|qN(f��J )�}-�:!�A+M"�b
q���H:'�B�a,^�.�D�Ā�)7f�s�+�)��XI2�5��I\J��T!�k���� ߈<C�$�|�Eb�[ � m���$H���N�4t�]'�GK�N��!0cls�?���A�r�+`��*�;��a��"x��y����d4,�
	s׌l�A#�m}Li6�F-D���{��m���]R�Wp����g�q��ˢ�4*��ϒi���J6�C���w�f$	h-3a�:�0�)�S-ň,�ڦ��z<�:�d��>�OkM<�$�^c/ٙj�n~6�HF�S�x�iZ��>X����p�=��Ґ�5�R���j��	��6�F,2B6�O�% O�>�
��:�5T� �p���Z�{��}G����A�����H�1�?4�/[V@���NR?'�I9UY���_j��,g��1X�v�7��(V�U��k�P�$۬���l��&ݑ���Ͽ)����א���~��9Ms�a\�GO�7��ذHU��@�B)���o�M�,cK77ܥk��:�[s yި���[q�F~N��)��ϡa��_7FeJ�*"vD�Z�_��"���گՙ�&7ӭ6K˳L�.�R5�Z��"T��v����*O*v��t���T��Ǜ��X@����u�_�
�F����l�\�$�c�ȋ
�_�>�*��X�d�g�^t1#{�2 G8 	��VVwbɶ���$q�8� �Z����0�����a͙M�1 �y�q	���wZ�V����C� �21�ӵ�3�C���ԕTJ����2FuOҋ&�p�3��o��̄ٲ�-b��t쭵�f��l���yƉ
 W�v8v����^�D��K@J.�Tǀ�^XJ}z�7u��F]-�1��f�2e
�$sRa�{��/�]"��#�T���T	�p��# ���koT'B�#V�Fi��c4�����-G�2m�-�޿+��Z�yVM�ea����2��r4��>҅������Ɇ��L�f�P}P �I������Ѣ�G��`Ф��� þ-p�vw��8�)�cb�S%Y�"@|i�_.q���z�?��~�Pz�W`L3�-��%9 ����}Hʕ�Luo�A����E
dm&^ww�>K��������D���:�?z�btw�~���`��$=^�����?o8BfU�T6��8���;��g�S��r��K����g��l_'��d�����C�8ք��;}ĳ��It�f�N��d�';=�g@�����#�~��s��[��fImξ!B�U���٫���2��^×�"7U����Wu~����ײݾc��9�n[>��}��^�%�-��vH����1�ǔT�(�j��)wzv����>�r��$��G6��m~�D	�v'4�5�BC͆��&�80����v,w�x��GoG��H���&���bi|=�c���O~�E��Q�C�]�CB�**m�X,ժ��!�PYq&S1^�]�k!/�i���1X�N���>��[VV:#)����)���Ž�rhl�<t�p��\&�����Z�]���KV��|�w�10������Ǣ�C�V����U��>y&z�k3��r���64ޡ�����v�{}̐^'�������/�jLH�^�)���W�db�m�E/�v��z�π639&��� 	T�Y]�5ޑ�m���I���B����H�i���o�0D�_�����8�A��6���Q���0o�y��P�����s�Bn=t�3"�hq��2[|�j��������-1���l�T�Zd'�B�s�����O�u����/��<�e��G��e�aW���k���=&t�X9U��Z�`P�U���x�j�K����C�Ȧc�Cl7��ș����H�Jm>`x�m���]e6w��{�W�2����5Q@�#�ؠ7?���R՗���,§7�r�e�nq�4�"(���f��D�Ƿ^�#x0L!�t7�\"�Cm��P�p��ŋ�''z���(?qSK�B�%���mG���$B��;
h;7�'&���qT#�J4e%3H�����������T���4��@6#�R?� *�/�VU��a����KD��uѸ&#q���X9x4v &���z� *��qӲe��p���R��0���v��fk�W�.�QX	xq�K�X%EϺ�m	�@��7>J����~�M35m*j�B,�Y�j��k	��<z�����ד��|W�,�ݲ�i�Dh�>D\���t�XҤ�����{Bia��nit�;�hk���l�V+\N&4�mcS��PE�;��e�ؐ�"#�Г�<b��t��;��M�e�3�-��S����TG�^���q�:˧�����b8��|��^TT��?�>����A�9�����K;&f5L-|�yI7���.@"�6�6U�x�B*MA"�3\�*���|��1i��o��$�_�/5����th��<M�p@IW�ٚK�{&bACs.��܅A_]��٘��䲄;���N�������1Ry$>�Ew�Te�F����.ue�̺qN�a�x،Vk�v����m�Uҡ�?
�{�6�D�kez����㮜\��-����~�4�ϓ+3Ѓ���|7��W�*��H�G��Q
�4a���گ�M���{(fc6_f%U�R�h�!��c��.� ��a_��?(��G�]�un������W�}����7p�"������$F�b�>�j��Um"e�ĝ�8����� ��Nvf|��Tǔ@�.z\��#y����d�'�I�K
o�[�r5����uGiےGݝ9��\F �"��A�����´ß?r�L�)$���S�]��ª
І:`�g:��:1�M��3�!=�l�ч��!5=f��-��%���bQ�h�S�-�فF�7��x��>���jE4\%$�Ӏe�ҸdUzìS�˔$~~��%7��i���P{W��gϰoI���K;G;�Cڭ��ʵ+�x٥aQ�&7�[��z���df.֢E�i|�\<U\��I�l����	�=;�e�*�0 �F�2&�-Q��9���oV?
�٥,�<�8$|%�1�� �'��ެ�͕�T<C�Yq�/�h�U�H��U�n��Dy}�2�cĩ]&�M_Q�]*�n锚r�}��d�(��O�tY-��@=:����*jR�tWݤ8��{:�ɫ��2��F�c%���&X##�R|u}{NT�Q�V�p"�܊��d�If�-dA#�>���8YzGeG����R��UL8��6i�MT�2	��O�6/1t�
�ą}s����.����]�#.�)�I���4��H\1��[ �[ *�=���ָ�@i��nI3܎\4�,ހ1d�9�e�E!d���cü6���~�y�Q�f����O��7T,�ׂϔ�7�M�qr�g�������L�����0��1�Ԍ��i�N���_K����S8^��2��4(�g~��sptT|���Z��V��#OZ$4�>],��_Ʀ(���~T��B�9,��a�SUI@6|Q>	�@��)�]'�,��:�ڪ��B9���Z����g���wD����@�.���o����k�k�F/���RB�h�.unĶ���G��c_��q��zP��ܕ+b�� :�D�����K�+��)�TWR��
<�(,d􈿤>�ﵩ,_��w���a��Eu��ű
���tۛn�m���SW�T-J-�
0c��:y!W{Q3�\w:>��g�~7������C��3,4�����R��BKp��v�x�-/=ê���#�L�sZJ����+�3�µJ��Mm�DC]�*зK��o��鱘�ѧ�+{�E��l����d.��@\:���#�n���4*�}2V����Y��,m�4|�R%��/�.�)n�-(�Xx��G8�a��h���wK�<�@q)��v��}���6�qQK�<�&���̳*��t�8�q��mR�<�<��6{��`<��E� ����ͺYB�//B#%�cm;�^��VHʷ*w/Yj\"4��>S@=�N�����u;��gԇY����'�z[��{ Q%�C!����f�wz'��L��ȩd2��I�`���T�E���2 ϟ:���J���O+����	$�{��p�jB �j�-��������nx�"Q:4o���3v���x�R����jlq�>��'��wS�_ 8_&
-ji0�Ic��$t����rO�>�?vP�����|�( �@ МYI����c�� �P�5�E�G'�4�wU���\��͔�xq�u�U4��J�g�ft�Sw���h&�z���6��=� e�5��梽����s��z�AQ���ȉ�CNR���<q�4�����'�1RBf�N���tPl�E���v<��~�n_ft�)h�-|��g�A�\��3�ǃE

|Ep(�����2n��*0����O�27��%�5�g������ih��#�[x']�x��