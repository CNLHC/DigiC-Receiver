��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���5p������H�4�z胖U��'��$-!��M�
�yx7Do��K�;�-����u�4�m܃�Ϙy"5De�#��
�k��@��ϔ�kr� ��c�m�L���/�dRJ*Kh��v8����@js�����ǈ�5I����C�.�@*�ת������:`��"���`�4�Q�����2���&B��bY�=<)�;�ӄY,b�BY��9��e��V'W�.�L��M�)c q:�F��L�J3b�}(\-(��&~?o<�� el6��y�l�6f�(3|��6Ӭ�6K9m���+���BH�L���-�NF�l٧4������鎷���Å���g���ey����⨈{Y�����,,�@��r�]?�:jM��o*�A:��%e�v����ò�
Y������r�7��(����pڭC0\W������ؽ8�{��f�(�5�AV)al�e��{��+���L�gi�$HӏY�ܧښ��a>�H��)��{Ee�=Æ��·���!����R
>T��,�����=�������E�:qA�4� R�^	��!)�1X0r	��<%o�yWjs�i=^����ߛ�T3�Y�0�B��!β��T
D\��Z�{����H�"'�/��w����l���;&1t?1�����:s�ގ{)�
� ��x��,���������N��M�����U�,6�^�����0��jSD�X�3�9~W��qFF�J�=/���ҷ%Dc8�ߤ$YT=��{���2]�E6�u��L	�pU�s���Ǉ�	�k#�U=h�l8�Dn���{@��^Rt�n�gBb(rJ��m��q���+h��<W���c�j_^��4�OrЂ3h|�?���s��oH��o�cT��G��}�M�=�S=?��oF�/O^o�Q��E�`zk�v�>&�P��m��*�N(1��v
$���B(@���W!yw�%�dWK�}���>��A�j�( �"���X�����$�E��G8Zn�ܱ���uD�u��8�I�&}���B��a*���_��pVJO�RW�<_�g�x	Ů��-��F����3)8�I�^e:�����>�� Q;�g��1_��ݷ���T� �ݿ�e%���A����+`I�����3E��i{����zb&���10f�����,Y�Ԅ����{�i�l;�3j}Z=܌����)�.��-����4�!����NM ���j��T�q� j��6Cf����&��
�?+\��s&v����Ax"~"���Y���p�I3\�����͒bl��,'�0!;..)˼sp���
Sx��8�� $tQt�0����-^������w@����#����$����	Ģ��[�_,BR�u�J�w�����]i��(M�/���T� �R�޶%�$"�]�ЗԀC�b]���B4�5-gJ�b�2��|w��k�8�2���N�k�T��@�Ϭ;���h|��u���h���c.ʍ�NxǸ�7�NMj�FX����T��%�Ng"��C��~�V�I�!K���9f��C��O~u����]��yG�~�����ֈtWODZέ3Eɴ����C�4ۯȹ�~�?�
՝���Hb��Da�M����J /�n�����,�}e�*�x��#��cd	�Q�ă��~�J3�����bV�[r�i���.����� ��n75�Ѵ� 4,�i<ߤL�K�fCc��/��Oq��˳ԌEک%/"I���G5�+�ϻ�%t�*�� E���^>7+]��9�"��5�s0U 0F�p8�j`���x׵��]�?%��`����@$oO`�pP0���!b��6{*'�Q�2��4�A'\-N��"޲h�����j�AZWT�J�C����ǀE���ӄ�������S:]�:Q5]��īg㾇��D:�J�S�A���+�ǖW"����;�.����!��TΧL�|(���y��m��\�-��=<X��c	=
��|V{]���f����zt8L �!e
E�����5np���"��I�˔\�Hۅ}�[YX���x���
ߥq���u>�1�Ir�ф�9Fʮ��,����@��O�O}d��1@�2�Ģ��������؎��k5�)8��N��^����u!�&��f�n���K�JA�uDja�����E�dԠo���W	!��	I��M ���rŪ&�N�Ҋ@�H,H�.Q@���.'������	T1��}�.ٸN����H��U���)�@]��͕ח����,;Jt-�@D�a�+7��m�(��y��q澯 �W�,�Uv��YD�N��wW�F������6]3	"�p��ڹv�߇�_p"�7��i���F�c���m�^C��,�=+�p���R� 9	����'@��Q����
��,� V+3&�C�^�k�lȘ�-�ӻ�'��s�O}�)�:��_{x���@t�|��E��=�MB��}ߛ�㾟-�<�:u�HY���d��3�TJ�.D*��/��X4K@ϧ��L�C�~�snٿ�C�GG(���8���eas�U۞~B)i%�n�z�� P��8&�ۈƋ���Ny��*l�wN�Y�N_V#J��R��NQ锑�PW~��e>���~<tuf6��`��=�ǵ�� �U�����Ҧ�C�Ij{�`���uRp�["��P3_�$�0&�mWL4�}M�>��?���`��sw50v�����(���;�ʒվF9�c~\+����j��b�����πZ�b��Ϟ?�K��e�@fj���J��~V<�--�U��=.�g��e��⿔���ٰ`�2�� V�B��	��>��`��Q�R�F�����G�����#iי_���ƅ���*���c�^5h���q��7���.��|4*�'��`)���mbVa�U!K��:�oh�=����jZ���ݶc��@�Q��%�[����_r��
Oz���|�&W=\�,�j����C?t6��u��LWÈ���m1�O2��G�����׀X������ȚGg���U�~~:��Fr� *q���<xb� �l���0dky��F��^�a���q��R*J����<�q����:����Q| f �]��"C����@��8���̑i5��x��]f"C���Bo:�I���,o���bh����Y��REc���
��MyWjg���.t;����\lB|"��B؂�X�T!��o!Bʦ^&�L���@�jz���\�^^���=���Y;网�����: ��+v-^%�":���³OI��[�|��`QI�����e��3S��%�$�Ց���-�����N����,�H�Q��ݎ��B	wch���/	U�{
��=��wLR��P�ސ��
�5U�!��(���S�,�ԇ�C���4uuUOAg�쨧�����2�17��.�nV!��1���v@�X��A�L�]l�-�y
�Zb�����V.A����������h�
�ą��~�j	.ϐ��C���v������9�lE�V��ɠ)ݪI=����{*a�,d��IB ��EVp�&�wSHD c�I���������~PDrX���`.�˟�f>/�-f‽~�.��|���@P}��v[3\s�a`Sw��x��QN�<C�b��E���I��w�����> ���C��/���x�	���$�&څ��P�ߐ硾��=Mhj ����z^w���ߥ��1��Ȥ�m����{6��%��{�;x����<,l_��z{��l?�	�"��t D�-A�-����
������e�m��$�G��>|<}���]�6��ךt�/�������ߴ\~3�#R�"�Rn�h�R�ٌTT�Q��ty��0�9�!\������ ���`3m<��8���(�~6��"����Y`�V�#����==|�H�+�Ѣw�Д��D���1��h�7��c���	w�hD��A�a��%���2�D�	�̐f3x�������q��2RZٸ?s�fq�ǰY��v�ٖ����
��I�TҔ��5�{���{Z(�K�V�K_u���HBO���N��T���ei�	��m��
!�<��� �n�pD�����E�ϋy�VdX��;��^�3=���'d��b�:��]S����H�U~�b�# 1��Ԧ�����t�T]�� �@�E��\��vꨳ��K�{�g��6y�fpF��/�2�i@�5W����d�Zbb��i60Pr�2�Nv��1 ��L����S2t��r	-x�%?��{�ΐ|�=�Ʊ�s��k��˅�no�G�0��Nv{>`��"9���[�y���aN��3#t�1?�馮��7\_4[7���5�q�ϐ�V��6m�1�X�;�5��q)�9 �;�7�+އ����C_aC����W=�!k�HW�fz���C��R����k���v��,`��<n@Љr4~�ƻ�`�'r���ۣ�	j��3�غD���BY"���4r7O�� ��o�c�KΡh�.�CY0p��Y�ca�25��?n����t�/n�����%ܳ�fS�G8hkb5C����g��.� ���`ܞ�
J���)6��OXS�5� n��0�i>r�D�ʴZ��=ϓ����ۄ�qD@�{������C��<F���cّ̻ҫ(�Y�MY�6ܬ(��� �m��x�����|��L&�-�b�#+.��I���EXɨ`w1\�;���P �QN�}ol�g>��n���2"g��,MF쳮r�p��눇<\7���̿�l �T�kz@pS2ڷ� �!>���0�ճŮ/Y��,I�d�6N����];h�Gh�0q���nqU���7�/���o����.�k�{B��L��fӰ�x��\~��d��cu�v6C�M��d����/{A���_3��\]((�V�M�h��^�.c���a^P��`V��7MAk/8�0~�Cd3�\�r������!7��)�GW��O}#ܓ���3pP��iX�	��`.���pD;�A�/�-��\�$��S��菉f�U8��*�3�T�S/?��bbh�h�tCL	�οť����hR�o;Z����D�:�"/�} ���dcp)�h�Ğ)�us�3��(��n@6L�-�3t-��4��"8,t8��6ܖki'*>C�"M�<?�MKlc�d���U���U)�˵�޻�j��__q�t��iW�@�ճ];m�TZ!��g=�=Ir҃��t���c"��b�W�~��.Z�6���������8:�ȶU]O��9�!	"�U��d�k1�d��j�%�A-�_Jb�u�b��������F�#��=�s��?̧N(�h����
��l��@�|�qm�I���f{p�؈�4bm��ԩ�c׺WP�t���8P���h  sZ>����KbjJ�Jsi�R��m�����W=}��,���]���-.������l����$�M�����S'w#ȗ;�h"�����$J>�)%Ce~!`�C~���Ƹ�Q2��Ub�9@�6�λ��ɿH���� �_CX��tsY�{(�,����������eu�(������,�Ek<�r���ff���Z�X%����Do���-u�1ڰ�T��|,�q�r��#���f����4&��2�������X�3��ѓ��Q��6��ƪ���M��:X}�n�>Ȑ0vv$�{�E��.@,���r�:"��0�u���L#����3�vZړ�$,��HD�o�t��T5F*gZ�jI����˅W�l�6�C&%:������K�NS�}sz�ѥ��
�b�x� we�
r�'\��*������ G#�/{�9&t��EumV �-����<,��a+�Be�r�����&5�ѝ����2�����N�U��*.ZP㑥_)A��I^ʺbX���D�v���|M�F�݈���$��%�w|q]y&���n�+��1lw�y�+ǡ_Kn�q�f�e��ڏ7ĸ\,~��'�~'#�c�Y���z�a�a��!��Y3:��/��&u�ߤ��#�`J��V O\,�py]��f�V�"��Yq����Ҕ��&�>�f]��Ӟ��� ���#�c�;���u�6��J��L�b�"�!q[9���"�]8�×�o�M}���0�����1����x
�p�����-#88��	<j���v�-��ɽ\v��OH\��a����QHv�d�E���Ԇ�hD?���ޣpVom�u�����~��ghw�H�����ϻF��Nҳ��/,zhıeDɺ��N�q���o6�]Zx�aER����� �.��,�"P�ڍsjM~fq8�����jhh��߀��0}�vB�~����J�������c����uc[4Ze�}�NM�X�8�)�9qԀ�IZ� �]t�cy-�m?���D�<B G�x�%=m�e���܍!TG�Yx����8|q��k�����g7��� PTҠ��.���XleЙ�V<S֧�R#�@Mˉ ��� �B��A��`����/A&��:zX��!yo��]�c6B����$����Eur����?.��ކ/��eC��Gߔ640��[�i�����O`��+j�^�W�]���� ְH�90B����XL�7g���������/���t1yYC9WJ!�}�L��&�?J�?����6HiC;��+�1g6�v��*⎉�����Υ� 6R�p~;y�����kH
��$�_��
�K�j*���x�
_@Xn5�f��E� ��<2��U��Ͻ�v�������3��C�6�c����K�;8��6����^���fu鄨[����Н�J:�
N�w`�P?�4��C6����9��5��D�PG4Ρx�k+\�����ܰ���Q�56�ɏ�6E�2t�D$~
�1%�ր�kS @F,�l���g����~�4_�l)
[���ŉm����	�}�10�3����q� j�����L�[m/鸜��Xyb;���sð���8`���PO3-�O1ID��u��U�z��䐟�q��x?T�P�+�,a�E��wl����5>g�$>�\m|N��!����˾�#����Co��<�7%`-ʄ�많a�O^��Ȃ��3�X��X��<��%��e
�g,���i(�Kv�C�ec���AM3`I����}a?���b@	�}�e���`K6b�m�i@s�� ��9����3Đ�˒�������씷N=�SwB~s�]�_�<)�7﭂/ �Qrz� x��L8�ͤ�;X���u`51���px+��S�70�+�Ț��:��\�h�AY����=�b~3��k+�\ک��|�O��M?13�0L�$K�×`��(+�b��B�����:J���JM�����f-�Ft�P����?�LO���%��L%��2>,l���k��.*����Y���8w��$�8?e^>�^ a1�X�3�pP����Ò�c���׺�hs���P��yQ�x�����Y��[Ex����� ��u�o��{�9+BE~u��~p�Pj׶а�<�a!o�Pc�Xb٫&LH�8�$o#��θ�)��ƜM��}7�ż/N��rin��OlOu�6���j~�:�'�'Ma�L9���cAB+�ą���`� ���oUZ�%�u���k�B/�S�剢a�$����L�9MgQEG'���Io����<@�^�5����_��~�ێ �d��� u[B�ӳ�O)~�,���Ѕ�<��[����r�g�?����X�q�����CIG*8Q2X-.<�-ゥ�i�ɲGP�`G���R�� ��G+,��_{gM*��G���gf_��_:o��>Q\#��g���|ԕ�I/�Bo"Cܨ�BVI�����c���8�B�'����X�+-��9wU9�^6`���	�^~�l�t��D�e;�b������o{����#�0�����i�e��&W�N�%��;��T��ֶq����Z� &p��[�<�9�/U'x/;樤����Ĺ�3%�rLZ)��v��y�ˤ��&�����!:�P
.�Y���R�T݈H%�B�700z����}���ܷ��W�0�s��`���R�r'ǂK�S�\L�}�/�IEEc��]�%o\�U=��X�T�I�+L��_�jc��t�Fׯ*�4
T�a����*�tk�51��� `!_P��
SKF��*蛊�R�	�:���4�p��ŇQ�K.�!	g���lĿ5�y�72�B^�;P�]���"OZ��h$��$dz�])-��3����؂Muh}�jijq{�`+���y`���6�����������b�V���X�>5�E��u��
+�4%%��Ad��ͯ�tw�����+z�Qf0y��]U�8]fJ @6�#�QwiXD��bᔢ�,�c
���;4��B�?��u�_>�:,qr�z�A[a�oZNut3Z7#�!R��W�̒F�~>T&4�����NeM�O�gV��י�a/��i�v�rw��J�i���CZ[Q0;G8�́{�1�$~䵺���m����HJ�ԃ�W�)t4{�~짎C�/���7C��:�Wo%�i>�E4������	d�c��O��f�z�TW%l	���~��ݦG����@�y�#ܝ�d�X�X��$�$��������(�JL��ֱ/���zĹ 
�ŜW�ƚ����-�F�c^]i��p�
iz���'��H|�o1�jo��� DFOʟuU�I_[�\��,~���G�_����g�Ž� �e�sdtS�|��%@��^	a���M��؍��n-�5�y��s�ț�q��LM��O=��*ma ��2���D��~ŊVx�յ&�ۡ�_��@�?ʨ��������h��
W`���%霳�ju�9���h}}2��J%�20�|hɿ�,�_~UQ�Rz�`�)_�X�
��@�)�7���4BC^�U�����R�n���� ��[�ˠ@�F�n(`�����щ)�p"��i�4�GyE���EP,��)r��Ί���O7�DJ3����Bk��Ǘ�����Uh`a�{&���ެ�o�^W,X��bM[՞?k����[����s�.����*.�9�?2���,��@�e 	|����Nǥr��i��K� OB�_́@���9�^y��[���j��:������N��)���--ɸ���\��$��a�C^��ï%g�5,���24�3���\M�OQ��6�Vh�v+#|�\�d��f��*��K���ʢ�l�1��;���,����\\�)���,����VNs����t�:yC�aTH?�xmz�x�w;��AQ?Lώ�(z4�f�^�V�p]�=���A)�+�^5�9aQsx�E�q�b�xD~8�&�[B=�E,���V��� �� ut~$�0�L�c[�@J[���)֦�`ו��`��gL.�I���|��x�@j�e�"��T��cB�W�����W�se������o��$o��
L +q�_l�B1�9���,S�6�� ��PÜ��Vp��=j��=�S�t���i.��U���F<�#��o�X)�mZ��K�������?��xb=ӭ����t�P�LS1N֒���ƚM�=@;\�Ԍc�k��ӟj"��>J����gc����#j����lߕ�s�G�c���ϘϻhN�눙)�\5�����f�o�[0ʦX�U��W�1�?7[�:�|�x��R�	'�㫎��l�yލe�x�fO����V��1B�k�U0�������'d
�4���B�GK"��Cj��!��|.jy����z�W�h�P��2!Qv�d���7�����遬�P���r�HB�x[�#�2�\�G=iy$��ֵ��+R�hb6�Μ��� ��2nlH�|�-�?0?O �>�ȝ"�����pt�R$��9s�QH�p�
�ua��P��n�″��+' ̀畤rSN� Ǝ�
R/��N^��N�M"��5鋠��9��㮎%fG���x�eךm�yg:����R��{��ۗ�E73ppr��\�����~����j��̽������C�=C1t�~�F�VD0��@1�-�0&y3q�D��
e�u�Ž�:����2��;6�~�y�3m{V6�Z&�uݞd�z�6���E}�l�Y:V0����6��Ϝ��A��}JU]g�>�T<�0�����Ѕ4�|�P�8/�������Pv�s�4����B�l��6������	������f�&�ZfM��:k�����c�be���Ra���k��H�:���!��D���Gh��A��TNi��w���((��O�A�O��v�9k"w�e
0l�N�~��ě#�C��G�o�"��(�/�X�m�$s�ݶ��Q'Zo�vO�ş{+޳�������|���+��(�2��΢	YQ�a9�Z]�!�`�� :�F���p'-�5ƀ��?ĵ�U6yPP'9�IiW�	Ng�@B��M����s���R�è�U�
�#�k��3��U�������_%�p����@��3�j;�^��ڷ,����O�A%*�����c���$��=��F"WkF���?H,�M)y��<�,�j���۬ԿDC~'�u[h�_�/�Kڿ��eWws=�)YO��d�=D�2�B�������fz���\��_��~
��������h�S7����5���ƺ;�����G�J�~Ϻ����;��æ�|���{��$�+ìj��:�!:�@�U��F���Ƣ-/q�6�Qޮ	'm����e��Y-�S�a+RG����_�U�oa�UZ8S^߃#O�[y� A7��W+~��r��WIN�Ɏ�Ȥ���]ؚ�����R�Up����w��J�g�2ō�&ǭg?;�խ&��{�-�Ⱦ=�Q�?�B6l��DE4׶i�0R$��Q�щc� I�L��	�?r��mt
)Y8�U�MeZ����9".F�ϭ���o�y���u�7UW����ڮ8[����|fa���q�s"���r#�ܔ�b,k�8��<��^�p�+v�u��]$Ŧ���%��2#t�+	�8�ıE�v��e��P�(=d�)%-ŞVI�/͘�+���`JMY>�F3�U���交К��O|�Qq����<ܜ[��*�:��T�.�W��S(���� oB�7K`L-U��0m�����h����e�P`���9� Te�iZ���;
1燵��q�[�hO_�iu��� �*���$.��P�c4d��409�k�CϽP4�ɐ6r�ju�a#j�Y_F���!K���]�k����㞑����ޒM��L�"~l�/�����O3�f���yܼ㓩(��gμ��t"H�%��h�~G@�9U՚�=�G͘>SSV2�ω��)+�B�Z^�U���̚���zD~�������[��H��%���b�F�E����Q��v��Gn,Y3�A4r���]�]��y-}�O`J��B!j:?E��`�
���In� �Pt�ɜ�J���	�Ob ]�#��t�eqC�㰻.�FÌ��¹5Cd�[*F�MF.	�Em�<J?t@�u4׼卤/�e���Z:���;���x�q1>>U�ũ� �:7�<󲷡&c�NB(*8�_�gTTwn'uc��U�<�&���:B�u�rl�����z��f����ɬ����ƶ�T�o2Ce�
��~���x���ɐ�B��YM�^Ll�}�C�B[� �M��|��X��9W��{]JCB�)��$h	:u��{6�>^�F��<�"p�����w��I���^�BL��=UQKQ����$��MpE�ۇ�<�ٮ�	��S�z�0�^[`�-q�<��Q&q7�\�-�=}�|��Q���ur�K^B1�M'ܖ,��'��+�*���81�L$�J�HO��>K]O:�ؠ�F�۝�"����z��d')	Ԡ��u|��g�p�+*w��۶���@,~��r�pD�E��׭��L�w���63�2jM3���~������ʇ9�h���5��8��:z��X3�O�� F�r�����T��2|{@���ؘcm�G<�{֪���:�~��4:�d��@iL�y����J�$�ъ���J:�s�#�k�z~"��Z�p�n��H	�{��֝����"w9�<���PR��H��cK�A�y1�M~�d�RhA�Z�h�߀���ieÚu��ɭ���gPI�W�MA��"�?=��b�("�jј]K'�A(���r_���Q�'_�fmB\�I��Pg5�-	 .
Y�⊎��
j9���?�迁��CEj��'H�_��"N¨�u]ַ�u�K��9C�F����jH����6c������p�����گi=]���D1�(��A�3�H����8S�~f�dO�N9��f�u�fX9�%c3ln�^5��O�� ��"���߂���Xg���o,O$�xd_k-A�yJ!TE�GpN��0��@�v�M��z��~�
ΪajϹO�2Lk�b�?JچM�f��z~a�f�,ET1_��q���S�������;�B,�i����BL�����:ۊK�����d�4eIE��Q�����L����V��a�2�3Ȯ�0���E��<ʹoA�Y')9��j����