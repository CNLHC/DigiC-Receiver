��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ����u�SM{��D^4��E�`^�����A�6�������v�@���;�6�*��Jf,����1�$���	�-��I����L�`*~,'V��`�l$A�q#M*��G��Н>���b�jik�F�EU��ýϿJF��=�@��N�ʓ)"i�P��`N歏���ﴏ��i/f��̐�]b~�����|��%Ɯ�e2�d���=N���x,ޘ���LK�S:�؞xN��T�_�S�ɵ*�/9
����Q���X��^7�5v�-$Qv�	�
�4.x��Fa�a��:؆�>�e;r��	�Bh]A��!�UL��k���G(U�}e��G�wވ:ּ�MB�?�	�F����GE~�ED��,VsF���y;�.6����R~��5���2�]��[��[�Ɖ@iR�]���Zp!��Dc�r����K��7md��W���,������H��'0������O��	��AM���)��B]�ހ�E��_hS���)ZV{�(�S�\�#���G"g#�4?��M�%�垜1A������D	�ֻˑ'dYM�铿'�����咓�}�m���@�Z_�[;
'^�a /���(p��7�'Y��ȫ��J��2t��u�U��H�2�b[w��߰������|n��Q����֩�?��<�Rm�FE�A��5F��P�c� �L�����-|2�����QY0(�틛�&�=�_�<ˉ1�f�����/o���Z�'S��2�Z��@��N�'��u�r4��{��������� ��7��g3��+���`�\��t��ل(t�]����i�_߇{��+a����l)�\�d� �!>�&����E���F��6�0vX���:z���uC�/��%��Dr�PrB��vt��H~�O��@l����I?��,��H.�����9Xr�=gV�%�h�F�"y#����>�P�)��j,ڞ��%a��mA*AT�"^[,@4D`B�P����Y�Ӓa�H�~a�վ�����Qܹ(����4bT��X��0*�(���\[�$��bg�CNn���9,��[��n��bU�,���2�L�_<��Iva���]]sFp@�	{��޾������B��P�����3q?� ��f�k�};`l4��t/;�#o�Z�X(س�|��x����^ŷ���H©Dl����וx�Ύ� �9��&q!̰r�Y��z[e�{CC,:h�pЊ�\��HZ��_�4'Z�T��)��4��R�)Y��ò��OvO�|e'P *���s��
O��ش�s3*�6}�ޮ+R`N��a�{�'��C��;� f�Go��uľ��B�@Gm�� ���p@>�jTAj�C��szSp�&	��ֆ��E�9�lY�*��s�y�]�o�(h���H�]��'��N��:]{�P��3�א��00��'�j�[}m&�Z!w�,���D>M�V�=��,ܛ��SC��-'��tY���FK2�|3�8�Yd��1?�mB�A��D=`T��p�{�,�i0r�aOk�y5$oz������
���J/Ϊu�tKdX�)R+Q�P�	Q��T��:��	�/�O8H�9�˘��.�̜$G�b�v���a�nX�a�Z�D��Apz?�yk�$N���.�n<�`�|(ڐμ�Ɍ��92b���+��sN�#z���Hfï½k���l��9O����d�P�q�x�m	����D��	ѻ�8�
h���e1�_�W�ڭ¶�z���!���N�*vx;�E;$%q�և|��c�~ur����h�,��o}�+�,�� 4ꤹ�`�?�B��*ut����67;��1Ɛ����tt.�JVo���w��W�
L�4�����e���S�^[E��Qd5�>�&�1�reL/�Q����?�F�,�n^���)�_ts��x�w2t�d��? ���ɇZ��j��<y$dlx��A�-2�Zbپ�d�xE������ek��|
J���L��b=�:�?Ƌ�;���FMP�3y&-|f�BYr�+"@;���pXJ=~]��+�ZB8��3Z, �����A:mlKF����N����q�,jh��]�8B�@	��eӛ�R ���`?FF���!q�w<�R-�9���]-��~�D�C�׻�/~��c	��@��Ҙ��j�C�g�N1����O�U"J�	RW)�}[��H����A�`�*��C~�jd,Jc�|�^�&��>*{f2��̮�z�HVu��G�<���a�ݕ摂/���4(	�R�j��(=�GUe�<��=oA���>�A�F��3s�p�����<�
@C>_��T���v��s����(Tq����ka��{�pi|� �eps?A�4��s��re�6������@���h;��t�D~@{�����R�*/蹂a1�[=^�$�AS�����(}����2=�*�:�J��N{��5�O�Co����K�{�x ""-˩�u��Mx���������s�{`!�����4B�F�n2�U{m�ǂ}A|�7c3�i�zv�K%�]T-���2������,>˅
{�����nm.P�����=�Wɕ㊗{붱Ŗ`G'�����^ܼ�=Gƽ���ۛ���$gP��iS���d����U(��p��������n�@P{A(!����@βYb��W^>���C���������&
���Z��h{ �6�Yx�;h�Z�>���� 2Z�?ͪ��V�h[0B��0�$-:�|hk���e"H+(�5��h����)����X	������7�!���qe#nǱH}'Lج��l���g>I�T�m
@"�g,\���C�i�zrܰ�-���:��cq6ޑR<���Z�`�z|��f�Y�r���m�J��A݇PߘSr	e��gӀ�����YoX[On繦�)�-��VԋY�C�r�֊$��m8�s̡���dS�q��	\��J#u��.�w�#�jr�m#�e�5Ա-�C�5��Z6�q�=[3*�;�[:L�GK�G<��D�Q.�V�J0�h0�VIڒ��u��j���P�QlgB_+���rM�W��ჰ,;y�rf)�B����y��Z���]^2ۮoS߮-����^`��5A�N�Ԡ׍#KK.'M�,8�C�oS`����08Ŕ�+�䭙ṕH�,�a%g"�.̈�3b�}�#`iİ��1�VT���A�C<SF�ۼƎ�"��|s��&���O���`�YQٞ�:��?.�����l�E���	�;�{r��'����U��sĘ��a%U,��&6� ���1���{��A"p�� H-?U�tHo/O�
I/�^�R�LD����|E� �q�Z�]�z;��K����v{7(7��9�7bʷ(�X4	@���]u}Z^
� �0ѳ�f�^�����2�@l��v�!ÎTs�yT�`c»b��J{@,�C�`����>�piӺ�2)£`J�,7��{�+�|�����k�4W9X_����U��sqC�tdA��\���k&xo;��&���&�#A�Gy1��ui�d~ �]b8��@�9���qT��є�:�BL\��1���4��#j�2�����`���`)_IÖ2!~��3�޷�����&�1(5�ȭa|���'�c +�Pj!�D���>ļ���+ջ`���1�]�g�d�H��Y߫$k[�hU������e��*:k���Ư�%�c��p�{�@��Q�8,[T�n<�����Ԃ�9@l�}`�n��&���7����32B,��/�����@��(ӑ0ż��\]}�M�:��Ti�>��w,�Wg����h����~�ݒ{W'`U�!����Ags����ֽ�%�Bн, ��,7r�`x�p����*!X���ÐZ+�+�kΆe�s�?$:�v�DN��ϭ��)@G�ˉY?�O�߿5#����qx��Q���2(9$GX�a_�X���0&j�<ܳ?@�G��,3���)+4�rGo�'IB,��[�{k4���a��4��GO����$`�ȳ�����H۷�����#�1�7'���]S�]���^i��T}��T�y��#�t�KP���� �faf/[��^�%�$[�L$�o{����T�S~K���r���즥Mv�>gV �IϹ� ML^�Yԃ�{�A�o����z�pp���僐 >DQ��0�3����͊P������1S_I�D6�_���׎T�"��7���L3�I#D�r��a�����[-����4���4�LG�P�C	z�j5͋M���N��� 4�_�	vD:�.����I��l�𫭳�% ��ϰ�ƭ�X�5,�z,��s�$��]h�Ty����t"�\�N��7?q#�w bX��^L�v4@c`f�ȳ����t���>FɑA�H����s����� F��"�~�:I{�"��swն���=-_O��a a�A�W�mn+�0�Z|�U .�C�B�[�#�b�4�!b�3ϵphB���I�z8��rB6~5�GE�۪4=�簪(�g{�U�K���	^�]���ZwR��#���C7���[��(s�2YC�_��]��b(�][1���<�`S���u�P�J/*9Zs-��F@Q!z�le�Qz�:ߚ���W%c��֐r*ب������?yħW�>~o�{˸�i�i�
6P�2�hԹ�K=�l��Ɔ�Mr�|�R�4���f�}�v]5��x<̞�9�r�����A^$Pn�:H,m�A8���!+���k��������N4��c%�ix��k��$���y�7��"²��#P�r��~!ra�q�$���iQ�!�[�7>J����Q��J�{V��$���B�vFt����C�NbD�;��A�I0��2
��d����k�_l4t�j�J�<��T�"�
���98�t4�Q?�=�c>)ShP'.�������y�8׿�& �\��w��&5�^��Â������Vbi
-���N˶7ql��8�A*���9��o�� �1��C∼O�2��_G�����:�5��D1��t�5Ruȉ�kX���VtF���l�t�v���ɦ�u�zc-�"�Q�_<���k�i�@$m�����k�h�Bs'wOۛ��<O>E�1/դ�؝̫�ޗ��C���c�Z�5"�?sj%�Tt�)�M@b̩�[Կ�ݑ�?c=��hmL<���c�������҅p>�DTy�)1��{�J:7Z�o)�T?����\7��4���mݬ�Y�hLGq��y�r7�̍�_�t���<)���xہ]7�m)J��L�To!4"�u���R��*^뾶kN/���<lf��Cb���C�/q�ŃzvYūl;�r��n�	k`�{��������:�������@E�FWw¥-A�s����St�u2���:@9�}DmB���-AL��"�� �8,���b�)E��?G4�ĵ�CƢ�l��0UƆ�p3��,*���;�-	�Y5XL1�ǡ㟾E�ܝm����E���;�P��*э_Mk"�U��qb��D}%�;�-y�F���$������E��egT���Lj�:��5K�s�<�M��)�b�}'�i��"X��C(���%-L�⢏���\R@䎤�Cl��7��g�XM8��9Aj��P�ׄZh�����n�����n'z� n.��S���A�<��,�Ia����	"�ވy�1_K%��M�{>�0��B�܋-"W����n����j�i�>���a������5hݸ4[;I�M_3�h��`t	��z������<#Ru9,��e��'E� ��Ӂy$j�BZ��W,�5�%'�d�i����q̾���s�- &�L��s����q�����k�$k%e�BV�i��>k��T��G�`��{ˎ��P|�A3�%�t̖d��4+�N�XN*�瞬'y��d���U� �� 	E��ֳ���(1̮>�o����Ԃ����f|�+	�z�L%�m�Z1K�HJ`�%Fs�`aGx1^�^�D�r��B�p+��+g�a�`��7�.����'���Ɯ�+	Y[�ġH���^�v�x
&4=|�Q�7������ ��HVE��z�` �H�&#gr�'W.+�eỡ�j�ߣ� ��Rm6�#�a�`��G�e�⍯��@?�AZ�֣(Jt����S����(�1K>yb�`TuPq�G�U!z��8��F��g�$9f���n����CiyA��ջ��I�D����6h�@��A5��=gb�9��C@m�!H� tc8,N�ʤ��F�r���x_�6}9-i�j��B�c����n�&��cs��}z�[�#���Ge>l��5-�?��\9�4�_�oo����',Y3r��I��!#��Q�$1�SWOۗ�~���ŲRģw�چ���3�#����sy�^G%�2���:�3s�WGQkqLP�7>�s�����G��y���'��y��)�*Hﯙ�g�z��|r�7NT��Z�_m��Y҇h����4��Q0 �%�(.|�_�mw�R�U�9�����Dr���b��>��
H٤Tj�j&w��&�>q�Sr�zwu��S�ǈG����+H9{3��k�4qS�I�Y�u��
�Y(�{q@g�#z>���+�dS/����| "e&�%�;^��Nvh��PDA�c�!~g��("�	�A�M*�C���r;ހ�@����+v#H�f�IP�擡*��$Wʴ9� ��A���$�t�j���4`7��|���=��0�?vP�vC�	��s֗��hE�N�(l.��G��:{`�S�1��y��z� �8��b@�ه�X �M������,��`�Qsm� {�&\�C���R�}���ή1�	%|z�H�E|�)m�\���K���Ye�z#w��u�)y��n�0�q��<䋺g4.'�l;U
"5����s�%-�}Q��5'��ၟ����R�{�����i��f5�x~����q��<�������y:m��$�
/���'�b������"�QGw��p�'�!�6h���2�o˅�F/��,6�!8�����!��N]�f�y��Q��W5�i�d�R��%0��<�≧x�]*�
��S�=������٪��L�r}��r�^�����~���K��wM{�m��s�[D�+�#�8}'[�k�=���9��T/�����c(��5Cr�	�����4����6��q'|�2�ɇ����tg�b�j�ВL��ʙ�T�P�ĥx=c~-汘&9�Ki�g.�mԟ;&Ҭ�h�O��*��0-#��u��B�b]p.9�IL���ս4M7�čX����.������|/<�"�#:[5�R;,�W���������ڏ��j�^t^��kI`d"��K+	D�+���3�:]ࠑ�9CQ~�aҀ�L������2�-�y�[oG� �+�ʹ������O߇w�ֈ��d��.i}��_g8�/rq�޼��X�������s�����򖰡ܬu� �7B��1f��� 1��z7�gv�.F^����?@O-�<^�&FL��	P���=!��J�ޒQ{��OJ��R=v8�v&F�v��Kqz�ڑ�4��*����G��"o������������6y�;�mby�ݚ�����g�� M���.���3ʟ�냍�"�1_c��1U����}���U���b�`��bލ\ "�L �V�ZU��V�"⹿+��.�� ��w(lV������$Ӈ|r�W^ׁe�$���J�����&[o���19\�f����̯��QU�����4ks�
;����I0_�r�>��q�o%dj���6Ry\��Fe��K� z���T�L��E�5��|����Bb֫.ݷr�Gg�`iQ�I���Gy<��P-��--o�K�v���aHG��^�%�� Z���6MMI�-��ok�V}�Y�bg^�K4�4d�d�/��� ���U���|j��U���
P��f���ÿ ��(���]�Z�:���{	ݢ+vQۮk�D���;z�Y~şa*���S�o���.��	(���R��WG��H�jW��;lFy�i~֚�MZ��;8�&��d>ʘ�\d�e�d�P�H�9�nк� 3�!{�ɬ(��r��v#'���T<&�#��:du�p���l�R���+�ғ_�<:ßH"X�gH�6�^p�Ǫ��:6c���o257+'����
z+a�.�Z�	���"�1n�A�B�5g��s�d��N�:�0��Q9��9��ʌ�� ��6܄��A+��ڸ@�.�h.����Ώڃ$��?�yF5#�����<���]{,�-�#����ч�/���T�����t։��]�ٍJ'��OU�"��	�W�G���`׎Z�Z�9`=g!ɽ�`;s��r_��E��2���e~+
���[�-�-L ��>����$�s�/�.'��=J71�N]g�߫�=^$���3>�"T ��,��
�!��:$���,���0mԲ/��Xp�{�C�|Æ8 c]�O��Ԟ]>b�V�  �؆)�<M���.ՙv�)}r�&AR^�gy,���i�)�1(��m-��a�Hs={��Yz��.�t�/��Lh}*���ChS��ԗ��m�d<4��<�� @P��2n*T��,��2y
9m�~tTJ�0
v/B:ܛ�R.�j��e�����c�xI�[��f�U[j�zP̮[+4�u���J��i��{�^�6�(;1��Vy���D5'lLK�ٽ,9�����`�@p��X/���UW6|��w���<�t����x���=I���5�"�2�`