��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���P<�%���>j��0�Rco%Չ'�ߗz)�.	ql�I�x��N����1
���L�)C�I��Xz�ad���c�����5}h}��p�&>l��.�L+�I�a�/
�e��h46�Q�8�i�u�� �0�OIrL���_^�5g��K�n�\���V���Jb���Rv����0����˥��b�";ţ/�V�9d}���0N���~��X��/�������1s�J^�lq���Ѐ�jeN�P5�!�Ų���h3 o��/�x*R�z``��MHl��Uh�1�O��OP���n�,��EQ�C���Y�(X�����r+cv�gk/�V��BK�-�.����f��|��9�ڈQ�.�8�Q'}�0��8J}T^D�'+1.��r���]<��ۡ:Q�#�Q��+�-�vZW��b�y�� 7�;%[34;�IF`^3���_�d����Qobd`.!��v8&��š2f(��Wn�mG1	�����6eE?=3.Lۉ����T-;�� =�&u/�g�n�"��I3�j�����W��f��c�9s��ˊBGGp��n=6rئ���bdg �U�^�}=�6�U����k���D�!3H�p�8���=tp�gY����Aq�F#�����/��!���(t�%�x1�%�(L�˺�z�'���㈥\�SK%d>�;
����������&��UW�#�������(~P���G���`��"Gi} �(���V+���e:�p���Cy2� `�7��a�����W��_�)q�>��	��&�Ď�1��J�TM��Y�q�tj&�d��~��Pa������W�����Bp
���s�j��&�!�� '���Im��H+8�_f�����i���H�@m�ЧH1@����@Lgg���p�ͭ�h�$N�&��)-�S��QG=�����`hW��AZ�V��W����	��J{��:�+ޮ@��~
ć�}��Y+�5���-���N4yYM-u`l?���h-3|mB��Y4��<q�W�pL�~@�T�<-!�������9"��3���[Z��ЩƼ4:����٬����Uk3u�e�&�*�ۄl�L#=��e_���w�ٹ�a����T#�=�4���Pq$~Hn���� ��gK�u���l�5(׶��k�__g�����y�1W�E��n�6˝A�ƿI�����GMP|����x�@9=/�a�G�j4�Y{pT�3迫<����˷���)�i�n#�qE��q���� ��/�3p;6
l,����4��4^A���^D7���w��A.s9f/6Ɠװ�<�ߩP��O�h�.[�#}m*�� ���/<I�c$�������]pkӁ�*����\�ڞ�U	h0}�V��X{J��d�&N���;���A*[�X�T�Gd��h(�s���Rل�
�P8`x��A��QB��8���ך�_o+u}���X�963Ur�_߾�����F:3��uɼ�g�<���n���u���{�5��<'Et��+��N�y	%w��oɠI4��dV7
�4OT���Q6/ـ��ž����A֯�L��h�vt{�"��um�u G޸������cg��A�(�����J���ċ�*ME��Ғ"�bg�M���DEޗR�Np���c��>��ݶ�`�W��VÌ$�w�[�{���];���7�ͻ��1�+A4���D�w�����h~����L�l vݮr�䣍7�}O���||��c '�a{�n�Æ�s��Ӈ��$.����������߁�{r| w�����\�p2U�&���e`���e��aU�(����yNZ�;c,��/�iZ[�yA��r����^�ߕS�g��l����9#���Ċ��U���0�yޠ����b��J��	��I-�ٍ�����Ր�����d��U���۬�v��h��4���V/H��.�G$��FS>T�ֱ�A��Zj����ē����(UmS��_��6q�$����?���y�8x�4\�!Pp
�#��I��޸V����8tݕ��()���^̮�
Pj+�>)��?{�"��Ȗ`�~�����!Ssu<�O��Ϳ<��H�޽߆��c�1���3x��M;$��We�;G諦y��#d�j8����2C�ݯ��K���Y����h?j��6��#�k�.�Lqaѽ��4*,�'|&:�����=i���^_@=	zv�!��V�1�0@G�E��A�u=�u`i�d�����u�;���2�=#dd
B�I%5���pux�qͬ�O��G���6 �;%�ۧ��@���;s��N����j��@�Z��0v:zueO:!d д4-�h'����D7�駭�^(��PDK�[á¢��{Щ�IW#�収G��[�Ѭ虄4�g;/�K�v�t����=�.y�S��e�G�|	`�lݮ#Hf/YAv���-a�:���0!��r�&�1�Q�����o:/1tm������9
�T�q1%` ���E� �	��'�65��)�]�f׉�wI*���z�R�wka�k�4ld<��,2��QA�=��q����8�^Mu��$��������Ø�J�6,���	��a* b�s�����WD�[�(erBה*��XʄY�2��z�n�e���']@B���T;p�������΍��[dC��u>�-I�9a���u�$���d��feG�s�m=	$r�� �Weȉ��|n�+T`ߌ�ά��������&�A4��#�LA�;�3P��,�W|���*�aJۢ��щ��/蟒7�:7�n��=�+�AZŬ`����Ϗ��K��k^���X�f�T)��?"���ۯ	e_:����3��w��1�-���e��{.~�xT����Q��A�w��[QŔqv��6gl��q�}|$.c�?���2�v��c� �>�����vF"1ҕ]�u��8/:3D,28'5�<�Okp��8�c��u�jXK).�j������D�b�9
�)AYtt~,	j>�ƈi��`P�7�o�+l���a���FP"ƥP�4�C��_[N�����ɤ̍�O�������,�9��渎c�`S���^>�[�&�����c}�CĚ�h�8��1x���y�����1��������>��S�+I��Jq��Cl;�Y���F��[M�����LL5_����r(���~�9�!��[��o�'�غ�V�f�;��;t�L85���+��D��~::\}�����;�Y�Q��7����%{<��j�̬�<�8�}*,�J����	�p@vCF�x!V�!���j��ul��}�G���.9�+g�b�s���sT��a6XToU:��M�H�H;?'f*��Az�����`.��RgP��I���[�Bp����pr|0�ڟ$h["��E0�Yر�%^(���:'�Z���V�S� N�E�z2¨SP� D~'��~d�X�﷖B�G��_�ܨ��;��-���A�Ղ�1�y�RSm��3��P5=&��j\����6�q.�̙KR?8(��w�iv}�<*k#���Af?�����}�T��mj�f:3 ��R	�y?��5�N@�Єzߖ>#TS��n#����L�2%�X�%I�,��SRK�*�X�=�#�S$�f��X���36����E(�.T��~D!��������1G�J�n��>r�;efP��ݮ�"���R�:�K��X˾���Mv���6�*���#��U�h�>��{?�y#�x(Yu��ZK�F%��r��@���un���9\�z~٬]�?��P����>K�p 34X�iy�`�i�3������/�!��Ð:6V@�-�����W���UD���t��<���lH��?�'in�d#U?-f��~�y+�w��C~��ff|�7��ڀ��w͝C/��ŗ��52���f��B�**��[>~��t���iX_�E8�یz�f;yo�Rj�wG���,B�%�)}:6��T�Ĳ�Sʯ���x[��	g�zxo�
�j�Ytu�B��܇=(��dCө�YF/�g���r���`Ɣ�Es蔠���Ju�3e _灼k� x��H��Z"���� >�O�<��Fl�^�d|�`7�Ih-�=��Z�(L|�k#��{;/��L;��97���(���G=?">}����"�4oO�����l"N�3������32|�@�I�	������~}�u��X,�J�	,$c�{�Iip`2��M��+g��'����ǔ
 ��G���oN14Q�����~:�4~��m4�<�����{����p�5I\>?I[�C��9s>�)B��%TRET�;�YC&z����c��.���t<��)'j�@���ސ�0�zZ$�Shi>����{���s�O�Բ�RQ"j�OHP�MЖ ���Jዏ���ǘF���/���2�aw­�[f�*<x鎕��&s�B�@���]ϻ:�P�����(*���8(q��\���q�d������H&���_�9���b��X�����Ȯ�}J�v%d����Q5:bK��!����ٝ��{~�	�)�N�*+�j�LP������D*ym[x��<��KA�(�!d����ؽ����ԕ�_�D�b�A����k�1��lO}2������7�/MKD�ob��e�P��a��f�&'�G���t�Ɇb�-O�OL�`U�c
�.M�E�M�����NG�
^�1�@�_�����kS�^�^߃��)�����	��u��Wby.Ӓ_���� ���_L���t�v�7��&b���oaQx�/j�dד�J��'�^[I��=�!�B)<m��j���w�E-�C�i�{9��Ye��+�T�+"�+�g=}���m/Oʤ-E�qt�n��t[��h�@�/�4�1�Ѯ�T_x�5Vi�8q���Z��n����3����7�\��������}�@�g�֜c's~�յg�/�z�ꍾ�[�͍�_���#.��'8ZC���=X
�C�����g�R�Gӏ6�>{���r�����0���ׇ���٠�RXѡ�$wV�����(X�]��.3��%���e�E�,��hYzN�;J?���&L�jW��>��Ǡ���*�.#ۧ���9���}Np�ƍ��I��s��� `_0[�c�qnM	�R��çOh�.`���f����$%�"�y�����[�u�.��a� �X�l�J��t����o�l)���r��a��xoL��*ͼ��C�bM�RS!J�������ɨ?ʚ1c���t~�v��M�.#�w�o崗�����|LZ�q�����ư6m�xN{d���*R�1��ޤ�2nї,���m韙�W���?��#�� �����\��b!�<Ga1��6c�ps/r���P%t��pQ�[G��ǕB��ƚi��qW0G���)X��7�a(���w��U��+DI�kB��)p�,�Fo�g�%c[��ws�/Wٯ^ܽ���?Z�gi��k� }�X�?�ϯW>�U��=g�YX���ʙ�S�
*��(m���G�T��}�[ ��I=5�n�e4���y�3	���fu(8H�+���h�#	�-ݼ�9��'d��n��7�UI�.
���5�Xk��xD���F���/f���Ʀ�$,�"!��?�:���Z\_V��<��|6��Nԅ���J��Y�I�����i����N�]�����¾ŀ�3�^Yհa��1����a�:���s#J�=%Y+�k���e��n.ge�p b�: ��g^;a��5� ��c �ܔ�]L^u��7(������[�{,�<z K�c����G�M�:����������T����+u��	�-��N��~�R������Æ�ވW^�(<�d���uK�������q;7�s��Ĉ�d����Sޫ�I��՜B�]*���]�\DQn��#��P���5��K�W�z�n.�A~�%U����"�L�e�B��_Y��Dգ�����Y�Q>�P�2�}�5ف1�VqB�L>��O"H�E���<1k�j����K̥EL�0>+^p�qSkp��],ܫ>�ܭ��#��E���¢Tw$�!5���|F�+�n��d�;�V����8� h#Zi��(>N�)��k���c����� u��)���Յ�3��r���	�t��3�2;CO�{��Kd-(b�ˈEd6${�q��R�,��H  s���"���·Q�#�Q��M'�
�hA�^����>�O��,�Y.{HF�d4m,� ��VO�ܲ��N�W@fA��lW�G`~�� ��S������L�P��+N��|W�*�#�
���� A��%���*���<�P��7�&Tyy7��>g'cG��B�I�۩`�t�χ�3]�n��R۵��'tHH��	�f��14�͚vXnïj������jc$W�xUǁ3̊��]����������l�`��c?��}m�ׅ�3�u�{Q���Q����.7Q0�=Z��JNY�JN� ��)|gi�ݺ�\(���w;��<#���YkYǐ�/���$�|¾��:$�E�%� A��Af���Dؗ����+��Q�F����Z�[�j�(�u1�6iа��% ��y���#<`���:��aP�0-�������χVBZ��������2e��\�S�0HP6)�k�=�����V1[�ͺ���aF�Օ��20��y\[d-?\ip�k[�|�L��g�>�_I�������'�L��T�2�0ҙ��kE� ���<�����ӕT�=��>��T�6?D�oCn�E��e�'4
�d�G%�a�lj� Σ�a�;a���'�����s��|S$�p��vl7�6*B�͘>:����ߋ���0y�(�&�m��S-������3X����AvYN�Ocêphga���x�&��d��8�JɎ������.�����`�~�l4��XY�H�ډ=\�;,�;��W��r�:a���<x��ؒL������]s�L����$��jw� ��`P�����iΌP޶��Z_�.�!r�^�Q��\?k?������u`�����@ix�z,/#��^���Й�*���o�����$��.�� #>8H]͊P�3�clL#J���)��%3d�+��u�cb �+��e4B���+̚���ܟ~�n����j5������J�h+V���~LY(53Q!
�y�Z��G����vH���� g�7����Gs	
Uh+ia��<�GYQPq�����H<���s>
rtѮ�P!$���KvzYEk�8ů2���>'l���{�d%�j�7ݍ/uܸN�<W�K��1���Xd;���惢F{��"�?g��BB��5��"���F�&Sr���Lz��i?C��m&S�I�P��T~��^v��Q�B28���:��+!��@HONڍ?�+v�*x���%؍�.�)�Du�~i/�<����f��_�Y9��v\AK�0j�Qr%/���0��;�l�|�aS��E�zQ�X�G/3]3�1ʸB����\:N�wy�?ѮNy~'8	̐��]�۷~'D���1h©L}��3�ъK���T�mp��~�>;}m�"�3��a� �塰RzO�-�S�˪�w�l7��RŤ�=�UTq��,��T{�	�J��P�4�%T>o7ňe��&%�z��3���KFa	o��FP�����Q�/к�i<�@C%�i/rC�2����,��׼x�o��#OHd2;x���pDjY-4�e5�3X.�	�㚚��r�&9�1��*s�����I�|
�����4?��-I��͆f$�^��BÌ�!=�Q��w>��0�,ZyG��*�l?R������`�����:��f�ùw�V�g3VWϵ�FHr�I���z[�F;!������2l5#���]�"�0��m�.r5��� �TZ4�Ux`E=��r�b�sS{����G�>u��d1�	��e�'�ձ��\�
_��p�8x�k�,����ΌL���t��J0�)�d} ����6 3u��Ue��X_S��%n�tn6�2U��n%*S�_G��E~��)?��!���˜�h�|�+����>�<��!�ᤵ��h\8j���S�n+#*2IE�e���h���A�g��CTT1k�ZK\�V1�R�-QZ�S�^0=CĞX[�V@CoU��RA&l����Es��m|=i3�E����<z���z�9C�3;��|+�Z��$����}�k�	�<CZb�_%7��d]���|�Jd��,�9<§��SҐͯC�TM|M���*�zq���� ����d��̜g�3���)�|�/bd������ml�l�b�X�y �n�:q�cW��& b�GT����m�sO�����(��KVW�r;Nks�C5G�!����I�\p��m�/�����4��Y̞{�2���9UNB� +�r����Ѷ�v��ڼg"v�5�m'����Ɓ�Nf�!��瑀����X�b���%�H.;���VK�3� )��՚R,�?����HJ��]�ׄ�\��0'��xbC��ɫ�r:F��K�����6�a=�d�5� ����=<�\n�ZV��.G������i�o�Ј;����x�~���'�1��{ ����p�?Sq�wcP��k����䓝	�,�'�x6�$��?m�Xc��,f�F�XoP�F/`D�a�n9 GO���N��E��i%���AM1����K�۞Y���Wɂ.N��)ZX�D{s%����d�����e������'ɀ��3�S�Q��&(c�̰[�B?x�c
+ʚ��q��`��sAO�A�w=dF�KObw���v�������qS˘͌d�n�2F�$jG,����S��L<��D�SPbC�\�����p��Tx�CG�5��(@�5���/�K�Q�
h��h5)Sޤã�`����/�.<8�e��X,Π*uӥ��%�$�)4~a+K�S4� �3��6�m�",f�!wd�M��r~�rX��C�b{s�q��뮫�C3=�F�<`]�^W�o�z��Mr.(Ć��\O�+�اm��.��G�T��Q`��}�G�>8�i������'9�A�����V�#9���"�cDμ1	�b���uvovZp����?���TOb&��sf*kE�lWWhg<od�����UJ�8��sB��P���'� �E�!9ѕP�\��6#S:~�q�ؔ��p��n�|QM5^,E�´�R- o|1�j2[�ֱ�cF������0q̑?)���6\z�yyZP�gEܪ�����!�� 5��'�������wr��^�1iw 2���6�f-q�[�HK�0�p�ll�#�2����/�:�	RV��N�)yI�B˳���*I���ә��Y���rr�/�u�=)$\�
��W�WJ7�6l�M��� @�-3��pW�z����X>�(<e]`����{ݩZ�m�xH,U"T�Jf��/?�/�"���pu^)�*����͇��l�P�&�b�:=S���W��5�CUֺ��R���1�:�n�_΍��3#>�gVr�EM[Pq ��P�^�S�i2*�Д���X�O��^q� �#�dX}0zU?6U����Ϻ�Յ��T�2�Iaq�;!6|a���&Xo��$� RM������2�ҳ��,��N'/�m����;$���K߇Vl��:u�%�����*٤���������\'���|Ě4#=�ƙm��;��C~9��k��cp�HhN���Ƈ��{i���p��m�CY��`Y[}�m�#�%#3�� m o8��|�~���x�^�1~b�U޾�R���ir�ʺx\���_f��X������@�� h�QL�T����Ɵ�Vc�N��~�;<����d�Ic1Lτ�LC�t���8���]�o����z�at@&,d9>N)NQ����(s�[e�1 SΪ�)1aV�T��n���0O��~�8�6A]�n�U��on��h��r�6ݢ�>��J\f��),MD���n�D�c��(9�M���	����L/�iRUL@��A�t�[�!̒��>��Td��>_���\r�O�z�������ئD�Ô�~��V{h�}�*�a.cu��4K�����LM��+�mX�J~Zd�sz��?Rg��EE�:l��ML²RM?#PUS5$30ډ���㋨�*+�a����1t����Ph[��\�l䆆}�E��2`�#�J�Ά���	_Y����i��7F��ѯ����U�{�ˎ;h�j-�����2?K����SR�c��"+����w��Ww��B�.u���@�Ҩ.~d]�ˋ�f��O{8"��L�k����x�A�w3����jO3���k�9� 6�S����mB��]�����dp��7?�!�ň�4~_���Ƿg݅̌�U�l��T���˨,�|,��n�|b�sQ���aa��7Ŧ�޲j�{�����}3�m�R�4uq�9�W�[�ԉx7����P{��υ2�e���G�)9m�����x�N�Y��͌��5���{�KbfV����.. �}|+��.�T�入{ 3:1<�W�.���QjQAr��B̊ņ�f���/��7X�������m�6%�`D��l�����^���f�)��(������a�_t��$��N��@T��Ύ��,Y¿ w+�nr4X�C@}f��b{�"� N�v�uX��=�"QK9	'����������U[�e�S�Gc�G9ބ�Twl�8�ƱO��ːItĕ��:�㪍Й�0�:v�����.�L#� =z�o��-~��-i<�f[��(]�� V�jx������<�j� �ZF¾��hk�_�yk�H]!�V��{n�`�8\�G9@���z�Y��I8�q�/�K<r���v��V�'�B�V�:,�[����Ş�{�� �R��� ����w72�q�1�	ܶI{���9`��\����/ԀNx��2"�i	�����T-A魁hyJ���w���N7�������vq���=	Fq����骨�7kG�����:3Fժ:�k�Z����p�ON5;���1{���޿�Q:%��w�����2o�I'�v���>�(EP��K[Hq	�H�$���$��`sj>ർ����G8�'!� W$�|��ob5l���h2�9�B5ĕ�>PS�4L��P�Kyǧ�� �D�4���һ�|f�7F������:1X[��[�1aӃ��@�a���i�]��F+Tc���\-�Z�!YM�}�����xz4����S��{!#N�숟Q|۱	��g+K�X�ğ;;L���
2+�YA����S|����)cŔׂ-��(���I�����BoWŘ�c59��Pc��<a��s���3�r���5�s���ʞ��W��K1<�y��ߌ��նI�����%.�=�����ݫ�$�SjU���&$8���Z��A�j}���4���5W ��^����,)V�v�op�����>⮫`>��i|9by=�E�Հѓи��t�����P� O��u�j��/J��d.5Dh�D�1�u�E���o�1��u�
����#ᐕRD�4�D{����=0�WFEU��|�q�����c'������S��ؑ��U-㴏��s�'\2�c~<��}���R�J2�Z����cc7R�8���?��0u�[�5��o�WY%�MZV&�Z�ˑ����� ��=/3�ʂ�ۧߵ�����G���5�"-i�C�l�6��'/;:JAǕF�Ҝ�k�p;���9ZZ�]��Wo��L�M�C��_�Sg/� ��Ŕ��Y|oJ��_��3�r�Dh����� � '��}�p���G݃��|\��gec�X��5�ѝ`=)I;! ��Fw�}�n2�Cpq��B�g����NA*��a��hF%�5��C�b83�W��ZF�\8����"��٘� ��ŸG���	ޔ����5�c��h�H��z��ڰ��{g�P��$ZK�&/��]5�I���z�M��#�-�Zg�I?�ɐ؈�y�ӟ*\",����T0���>L<�UtGyv�ٺu4���h�<��	�7�8z�z��K�rm��o,� FWpĆHo��2��3�+�e�.a�xY��G5��y����X��,�ٜ��mĒ�$�C}�4Y�\�8��<�=��ODT��;`�-��݉I�f����(�NcN7���
���M��G��q=;�hRkigxI	��	cZG��}�]�hj�����wdl�+�>���-�����=�N�/5�sd��L9��v��Jw���!|lВ�F1������jخ�A�8����Gz0�x�yfg���R0۲0����O�o�����w���a��DE~�O���v�n#m�������TW�3���>��/:T��A��-�O�:XisxQw�z�Ng�R����5���ə���#ՃO<����DNk7�uo�@��~�LJ��ƽY�۳�[�VE�������g�.�3���lϳ'x����ȟ��H�@�Ū��q�=�|����_�K��D]k�T�*�Ht}�ڍ��㖩_��O�������ć�o��Mk}V�fR���V��I��h��e/��.�'��?3�Tf��$ۉ��P,�1;��ח�:�Ji@t��ѓ"�k|�[�=2�L��z*�Y��{e\w0&-�J(y��-͏wt��[��b�/6����_H�](#�Q�]^���K��=�5�Y���C�Rnt6G���=���P3�<�5��� ��~w�0���%�elg�sk���3���Į�T}Nza��)��å�������K�.5�{�ʎ�&��� ��楴�9����=��I#��}V�` +�&J41t:`v��B�$��#"��t�[)��P�5�z����fw��e�j�陼�p���q�k�z�����2���x����q�N#�Ļ;+W!Q �w���m�O�j�o*ì�UIϔ6�[	�'˼��?%]�������-��Rȣ�qpD|7B�te
s��"�/==��,�� .sPo��q���O�LB�����rɏ��c4�]��1��=gc�Ik�Uȩ?���:�5���00^ j���{�����jwYUU�h/uf�� �����i!�0_
���҉7�����Y�Z����˜qʕǻ�̣�x@q�n�q{^T�S��Y�l��?���[���j�(�m�����+X��į�xj�1�ql��l�(A@�R�#�kxL���@���z����.�~{�5�σ׺>�~�k�"�O���Ģ�Ww���Z�e�(�����]��˗�����{�-X���w!���lg`��8��a�Q���k��4�p�)����<�<iz���8z����h�C!;dJ���I`Z���<�?��l�ffK����`z�-'�6�?���Z�����d�"��͟�C�ªA����Ɓ>+����E���eft�=�.m9�ټg��f#H���\tZ�)��R7n&�k���`����-���^�� greg�.�;��1�a�K����e��~ή<�tƼ��0�����؀<�~��ϼ�k�x.�9ے�!��qW���D�8Ğ^�T���*}b)���,�Otc���fy�SH�g��:A����#V<����/��H�n��P�Ǵ���4�6}ZU3nF~�?D�U$c�M/���K"�0�g��P*�1���*@�*2�Īx�J�ΩD��,bJ.fx�E�Aǣ�Lτ��ә�X�'>��.��r�ǈ�O��_��wx�W�`G����Y�Hz����BI��%�8�L�8r�Pk��=G�X���8#mǖm���t#�<��B�D����A�E8�+��s
�Z�ڛ���`K��U����bT��\�y�EG���0��SR3�o7���gN�0�����q��\E.����l�՗�%P{Z`��f@:��9us�q`@V�t�ǭ�%2��X���WH&5*������Bޗ`�
�Q���,�^�ʪ���20/Y��`"T�ny���vi.<V���@�;�]㮦HɞXqk�U���9�����V�^��y]$ѿ��U*]�ʌ]n.�<�4U<>��l�H&�����b���[�FL뽥U
�.��4�F�u�Ђ���l�a��	�M�t�"��s��_K�:��ո���H��}Z��}F"��V��`W��ұ��i]r��9�%�t 6�4��C��B�9�ї����,��Z�+�9tOcvަ�
N��x(�L��.T��7��]6l�Y�e�iU%�O);��<�p�6�P*e�ɑbmti�8��+��+��Jٶ衔�X�'ÂJ�j��]�T��`�*[*R�J}N�����|���>a�?�nm��	@)�:�����F��R��Q^0�����#��^H3X'm⿖��2���+|�F1c����
�\?���źGܓh��0��3`^ �&������M�5�k��m���Xp|e��c�;�r���uqB�����)d�T���h]t
�D3�_�t��zqPu�x�u�{��~���7�)�y�O�Ծ���|z&z��ed���z(�/u��=�I���q��:,�LBՄQ���h��2 �k�3��t�8X�������'&]2�s�dLb�5rV��d.�b�EDU(�S��X��,��:0�Ӕ"-��V��r�H>�Ԭ.�}�A`>LC�n�'灌 y7��tYuI�z4]>F�?k׈8�t٣4.\m�ĥe&0[��Ө��H"���s֩��,��M��M8��<`	S�ߝ��,'9���8� �55����!��P%R�wVO������ӽy��}o3rKy�R�d���9
j��&��/��!��b��3n�/ɢ�j��(�}-���4�������v =X�HMa����?�x򭿴mu���xv����[�1Y�/%�~���o?��9N��a[�`�IA&��p�]@b0)Cۨ�%��'}���� �ۃa�w����>��=�����fS��.x3T�c��� b��u�ZC�ܰ!*m��H8� ��]J�6n�
E�,�ϛqk��yǺ�dՒ��=�s�<�#(11�Nr���	K�;���u3���~X��y��ƍ�\�H��� ��:Ò�э
��i(�3��$
���-�I�G�_ܒ�ϗ�TWh��ƽ�����v��\舄3<�C�fT���-2ޫ��*'��6��U;�V&u���Vx���Fd}�L��Oټ���f��}��3�����!�6�v����K$Zdx"t�L]+[��VJ�wa���W�����q�^7�d�0O�J:��hT��9��n��o��any����$��e +�s�>7�30���¼��� `p����~X=�%m5�ǿ8x�U��h����V+�8l�1lC�<G�&S6�R�f��C�B{|#�l�+�.qų��RHy�y%���:�� �jR��6x'-���"<�`8�+7��הppew�s���o����9�M��|��B�Pc<�\'N�]춂�
2^�Y�%��fL����.rǗ���x?��n��E<k�օy#*1�y�SS�V�[�2:�	P�J�ZP�Ah�l�d��g�`ߊ�� �!T����mWT>�KP=���'��X�췩��YY}��J���zoZ\��N� go_����J�!�LN��9&�;]�t+� i6˹�8��n�����a,LJ*D;�h1��n�9/��jz�N�������������=���V)3�_�D�
�s��A��;�
�HL1���_ԓ�Z�0���+�q;�cܱP����8T��;�j��&�.3�Q��9ܻ	EGa�`�P�4G���Э�g�by�U����q�ÿ��N�Y��g����F���YRP�A��K�ѭ� �3��v��@�b�[NY������)'$��[r	����.�?���R~��?��6�K�����k6y�
��I8����)�	~9���T��7nA� g����2s��̄ùL"��Xm�K�T��\��>���M��!J��ӽP��s�rI��ݍ�R�7P�?�Z#���X��!_��RM�-:��d�R��\�;�]��z�`�D��Q{y�"0;P��Hv�歐�g;�e=!�dƩp��(91)��~R�`�${y�]&����=��X�[gZS�d���+�c���J�[�wG
�?�J�ѩ��%�}�qKg�e��1��-�?�
����9�-�� �'a/́Ɍ���w�:��c��a�J!x�؃�7vf�º�޻Kr�D��h L�Q�����Iv�!�.Y��M�+���1);>8^Fђ�K�ó�8���;�:Sz����R�q-��Fk摇\c8�S��ԗ����j���*	��X�e(\���;SP��f�<�b�j�g��'8�z�BᓙMa��/�U���0 ��Q�b����E}ϣF�.�m��^"�I��U'~���W��0焲�N���MhD���������D`В8�f�� ����!�!�p�l�<�X٨�?|v�0�{vAhW' 9�KgV�n������С�o��3�b���B����ID��iQ��0�T�\L��(w�����'����{�htgؓ�4�Ge=_��N ^ڪ�
��S#L�L^V]i<S���)�,^+�l�iz�f*D��8�(�[	@\KH����7�rPv��C��d���Ō��������7V�'�'^�@~������qOe��1�*a�<tyn��s��VN�����=�	�q��p9�� /�''�.�rcot4��A��F�@:��'>���%89��qOS��FȆ�=��ƻ#BF�+��yq�?�^����S�h���b���(��W�4�7{]G�R̤��gv����*��@^��b�D�f5���s���%O�&\��x���O|73UT��.�� �?W�'���yG��I1���!Dz� ��#�pwL�"��U���E���w��y#�x��Z�ـ/�߾m��X���{��Jbb�6/�Y��ejȀ�S����x��l�k
k-����@��DX��^⤶�lg�JId�`
�Rv�<"4/���X������j��>���-z������L����N^�Ah>��s�%~�*,WL�&F�5.%�Y0�_\����E��mw7Q�o�?6Z�	L��F��I��J��\�_�E*/гy�6&�0��:�'%�>@�Z���}���<�_%�G��>�p>�#Q�G(D��������[q��0	��P[[t)3崣v#��]�h>��3o�%�*~L��Y^e͔v��v,������m��b	I8������BE�N��!`l�3�eZ�뱩^�@c24�GY�&�2�`B+�	����w�FQVg\v 	^�7�U0��m>���^�t�� ��?#�,�5;��L��QI-�7}Ԋ�da��)���X][��*�?Z�΁��+�X%�u�܍�O�^pp�C��=E�f��I�(�cd�\��[�����6�/�݄��2�)����J*��(ݐ�Z��a\����'^VEe��?\~��Y�|�V1�N�u��g-Z0.F��Ѩ�D���w����q���Cs��p����=�|����92����ɡ�6�`T(5��wj#%��������e�%���"���7R˒���.�+A>!����>�u1W=� 'kt*qO5#�A�u�c�e���¸URK�A�r���\��A�"kl#��􏮗�zLR�[���k���qJφS�2���u�uL�C&m��a��� ��8U��=�w�,�x^��y:� 9��b�JZ9U��q!Jr�����+i�qk�ŷ���f ��Z�G��X_���T'�T?.�_�g(��+�Τ�C쮨[�_�?:���� a�^��DRY�a5����]�?;w�����`�5�9?��@�_A2��A�a_5a�R�ڿ�����%�+pC����vm����"�����p,��*���H�DG9�*��LK�� ��Y\"]r�(ӕ�;{�R�2/���D��5!��X���HXV���o��8����w"�OŬ!��{ee}G����E(����?�P"@d�O���r�	�+��޾�(��E��F?P�P2ҁ����ɺ��@�>��fnt�J��=��)!����Ŕ�¬�Ɏ�Y�&/� �jǐKi�p2��A���n��ޝ|�`�;�w�Y���v���5t�GI���R��]n�����Ҫ�_ ��<	�!͑j��6Xn0K��?nW�w@.mJ��ٞʣ�c���W�=��߳�|��Ӱ*}��(��2.�N����ZX;�+ S?��_q�^ִq�/E�Xc�qV�uU�n{D���:x�O�g*��Yk='�������奃:�8�#���/�:Š-�\.);�*��b��r�Sy�e����/�
��;xAT����A��̏�V�a���q���i�u���/�$:��G�� �1��I|�>��b)�ȯygx\��n���>o�ƌ��Pæ���m�L#�TQ�v�&���\Q��"�_����5��.|�m�Z��H`��jQ�����`KA����2*I�r������C��I�z���QثF�9-V�������o�m��qq�|����^�r��Tu�7���<��[���+6�5
�l�^�v�Gd>R�i��5B��}�5�_l�>�Nn���#O�ip_>sc�@�]8���~������U�$$N8�a(�Rˀ+oC7�E2M=T���b�R�����R��n!b���b�ߝ��=iʋ�TB�c�uh9��BjE}!0U:+,�P��$��]R���~���ޤ=0RX�f�E�-{n�k"��7[:g�G�#1 ׁ=k�l"��2[�6jyc��P	YX%C�N�T�X��+n��ƀ��g��F0M���C>� ��-R�_�m��T?�e?`�F�N��� 0��8�Gkk �.]�ʢ�pUMY���mƄ��Ix�[����ޯ� KL��,iþ&s����-�yh���q.^��Q> lʚ�F9�4ҢB��/}~Ϥ����ۊ��t�\a����beń��Ed��G��������p����,4l/��A9�F=-�\^�5WLPjk�Ip4na�+<.�ϫ�.ަa�<f	�,�#��^�ǂw��(����:�A9�WA���������6���k<r����i+�nA@��~��0�D=�>�~����Ҫ�A�n��JuF�R"�LѶMy�GL�tC����e�w���lkv�g9p>*r��v�=��4�jS��qğ<�Rd�s>�{�ӻ�0�'D�?J�H��!=R
�Ҿq�0��b�{s�]�]7�R*�����G�>0�<���D��1;�'"f̠N�6��{<�͑���B����KF���=�.���vh'�!w��{w���F���T��/���[ ל���Wb�i(��SA�6�����C���S:~<B}�_�)ii@��Љ~d�����,pL4{C�J��8!2YRd�М�m�S�Y$�ק�b����4"_Č����T:\��~�S	���->%��L���z,Bӷ�tY�a3����=Ss���gaf`w@��v�;�EX��ɰ -�c_��Ȗ�i$�y��J��A{K��)R.����{/u�Vᒓ��zdh�b�$	��$���q0��xR�܌v4꿣���׈�vl�,��׍X��O��e����¨ �$x'C�ɽ:E��O���a���b-��2�'�0�R��ҾU��b�)��V�j@�l$���_R-�=Zq��h�u�� �I�f9�T0���y�a҃�|�|g���°�~�5��-�m\\b��܄���v:4*!?�^\��C�у}0������Fq=��"C�hl��<��8��Vz:�KէV @���δ5Ղ!�T�*ZC���i�7D����e�p��mY�&�݋n����gƒG�N��O`{�M�	|��ȳiE����(O�%{N�1��s�2S.<����J����w#1�کw���WK�eX0?q��'#@�D�r�R��N�[Q��<��Z괟R�6{SS������q"Hx�@5����u5�hC��\�8�Y�12;tP_*��s�%�<�Aj���0�=�X�?���q�����1���ey��p�^��`c"�d�\j�@W��E>�Y�/��\��64[&Ig��9�n�{�f�MH`Z�d�<��6�y�ʔ�_���M�,TגN~�@u\�i�H��[��vيv+����Yk�_���4�h��7�zd1o}��̎���j��$�;j"�[LwBY���C�+ҿ({{u�&-q�Q:�n�9��� gg��be�Ͳn�	7�Y���Aj�+I"@Vl���(��F�%�ɹE�I������<�����6x��`@���;Zs�Zi7⏃y����=��%a��^}�w}S���x�-pCN�s�kT�� ��e�kb��Z��2~�o i�=�N~Xb�ղ�oD��H�2��ů���n<cÆJ%քR�]�C�$�Dٻo��b~_ ��U�R���<���*6p��q�ܶ��Ϥ|s���x}{͆���͌�z���u��.vF׉꾪�d)��/���8�Y"�4�6-��[*�E��Yʟ��$s�}Av\!��qhH� �����\�"O��,���6Yvv�AX#�ū�%���F�%�żlF���-&t�����S���}��.K#���6^���	�K�A���˧c�Z�o�d�[G�\�;��y�I$�����ۼ��h�A�s�<7�FT�� ?խ,���!���x%�F	+%��NW�Un��<l��C#�Zb�ϝ�a�������4�.(~P3��|&۔�֌��cN���qR��,����[c�U6x�|D��<�}�E*�\&-ڕ�Ɣ	`'w���_ ��_��g���i�rG-�n����=��CiT�ހ��V��q+���w9>R�hH8�	:�g
�
n�G�����e���Q�	x$P��c�9�A/�Fq8l�l�E�Tqߗ]����\B�6�6�0"Ԍj���Ӂ�&��x֎`*۹W����-t
��މ���$��:���EĹ��XtNpZ����7���)l�|��%�?p{Ĭ�k)����#��Q�����S�4�K���t��W�K�L�>m1��\]��N�X�I�0�=k����?D�3�k߅��,�_������\b6U��1Q8� !FX�m����a�
��H�gWYj��%�=m�o���`�B�l�8~��h�eN2�Q�"	�3)�:�'�X�)����r>^
��ɢ��JZ�{}�Gm)r~z���RB�p*�5�R�)�����b��ĝ^�8z��_4h44s�Ei��d�"��7kQ�q�_�iv���J� �@f�'���쇡��2]� �>^�T�%<�L�K�]d��&PE[h�·��j�HpJ�%��Me��FV���w�K[��!�y�,jO1/�ωiO���+"�-C��Q�z��Q�͔7s�C��uR*
�{�![�-���HNu�*nWN-r�����*�0��6!��)u�C�8Ǡe?ż������z^�����A�mn��Yb,��ۇ�k��T�����Dt09��/�Qi�ޛ(���ƣV�T���ፀ�|бs)0Z!�]�X^��M�[��d�c��v)�Yy��Dm�-/���(�� (�(��'������x����?(
� ��]k�h��
@�>��cΣ��$ֱ�57FA����oo1�d�TGđ}�UW�=5�!n���T�H����5$,��`�^^J��D�R����>�X�Uj68����hލ�
�Nk=^DYmم~�΄l�ܝu�:�.��d��� #��wn9�l��C9u6b�F��?�*mz��z�19������#�m߫\k�<������F���h���-օ�Y��sQ��F�5m���Y�1MX60����l�S6|Ű]{#X�ق�r������c��*տ\c�!A���U� =Z|�\�H��j��"��e�������/n�4h4V�G�n��"�0=�Y���Z7֤�0#�k�����8z�&�#ω��IZ�|p;^G�kE��Vy�<�w9ǬK9��ƛT	���g`���\BϯfZ�8Ԅ��.�=�д�t���[]����{��W�/�t��Om3=��{J�؂�0��^�ڿ����i�<�U��3uq7�m���hr�,�H���bdx���P����t�L	��8[��UX�#�a�k�'��194D���د�y��u�};��m�v�"�։��
����`��ǘ�_N����� ���([cz���b���Ǝ�Y��["R��n%�����@�{w�4��r:��]�?t0vc}���^�sdw�R����u��2z��%��+C�P��E�К}��r�C%��h��6���3pX�~L�h�D[�ڵM�(p�m�p��P�x}�����j���w��,f�4��E`f�"Ί,�x֋V�8����j2���U��z����0
�I�J��8�Ɛ{}�c�-���2޹}�Q��;P0h��v��36������$�����tH�u�6Ǿ�2�I$e=��8�v�س���.��f�R��_�0��s�����r�6��$&%�.ԌqB�\�F������3d_�	B��L5^�_�`�q��G��r�i)�<QA��^1F�*f�o�#� G�LՐ���e���C�_�&�s��>XC���\��b�`B}�k\U瓡�]'���L����䐥��h��D�W4�E�Vc?��w�(o��D�p�4����ś�;�<Uq�i�p�$�}��~�	�?m��o�=&~��aŽ�l�L��9�w{����������@	3���+��!�t�a5�J]ᴟ��#*�k*��N+�]ɰw�W�v7&D��=��kY�?��C�V�h�*�p����e�d&=�����r�wAi�k���5>"�hwV=�E�{�[�RJ��=w�\��9_!�&BB� �YP�q�r�4�<u��<����|�;ާI~��v�<�)�~�6^���^u<�s%n���O��bG�Ǌ��}1���@��7���j,���=��+	S.zF��,^1Y�<:���-P����#� �`�V�a��D�?������C3R�˨3-u��c�y�<��	��y7�b�8��� �q��+>��Z+�_=t��	���N�<Mu	�(1���1�̙��Q�nC��M���K��a�q��.��N���NZ�Ծ3 C\_Ĕ_((8����]��T�>w�
!��Ji��ܺp�q\nI�+�o�TSo�k�| y0��|.z�-�_��d1�i+wT�a���	�Zux��W�eն@�=�Cp�(������{��}��I�KBF4�ϴ��i����XQ�o��Q�\nc�����$j��B-$r��|�;BDz)����w�����M
�wg���$פ��Z&sգI�����>i�y��N�3��<�)7��.��H�N�{e�:�/ũ� ��\��rċ����6
�QZpC�B��7M���9��|���Q� v}��'vb�n��Vd<+�_����7oO��m�7��6�~�`�_I�U�.U�e�g����w���8���vr�<j7ʓ"ΕyI��������� ����OXe���������;�7R�ӯ��i��`j�/��q�kr��r��,b!{^�D���U����<'�h�}^@Jo��@.nI��Vv݂�$�Ù��d��?��I����5Q��mx��)Adq���Z��A���]�ȋ�Zu�|ؓw�/b6C����A�#�/_�2Τ�|�X4����Z���- ��Tﾜ����8+�g�Kg*��xQz5ر������j�⇐Մ,�Y�36H��t_�O�Fe�j^��7Pv���0ov<R����#҈�O�]�S�Lí���Y{�D�+���
%R��J?�)oWЛ��gg8"St?�5+�9�~ ���(�����7��dY������-�/�YO"G�F�"��~�K�PrG�)��:�z�$#`i��BoF���a����q���2��+�B�"�⯗��0�?��U�Eܮ4�m�ջl�!6O�����aL�;f���[�=�sh�-V��P�9���j��A�=4�K?�#]�+	��'����Z R�D�n�(h
rI���D^�Y��u����"�B[����[���H����Z�]�r ��y�r�m�:���-WV?q�^���5Ŭ���Xߒ�=��˭b�i�*Xy�L�W�M=m�B9.�$�H��Gm �7q�./��+ە��k����{ʼ8��^<K���k�H�p�n������0���z6콛~����/V�nz��Y���;zG���{���d�'������p�ko@��1��Ea� �������7�ՄkKS��3�r��.O�t��D�h$��n����i9��v�$��`��z�Y3艕�=�)6I ��[��h�+�c���Es�ws�C{ʶG�{qؿ$P��~I�~��䡌(1��7XY����p)@�R}ԍc�_���4m��}�3�����M���6�����jnz��m9��G"ٛ�Y֜���r%\��]�'�O�\��i�t��Z�S%X����t�*0��_HȂ�-ǯ��о/�w5�3fD���ȴ�+���2��j�����}�M���X0ۉ����x���o	�"��E:	0��F<�tWxO��|������w4��POM/ص�2C]�:M'�c�a;X������H)���(Wf�"��#�RQx
i ���j�GO˖29w�F���J"�9�J= ���'8m��I[�?���a���,A���s���$����߹���d �Z�!u���47P��`R=�,��v�r$E|܎��
 ��2��_����mv���2��m42��h������O�H��n���o�
�,]�����l��#m�fad��ݹ�����d2 �i�
��,��ʠ0���4�R��%A2%K�H�a��԰��T�J~H���dJ�bv�E_=� �6 o��}τD�P[�:���;��V�Q7�q�� ��٭g��?�o�6��ms�̀��s��l��S�������GJ�Э���b�:���"�w)X�yy�@�٪+���R>�$O�[��Q��Uޅ�v�&�7�L��_�ٯ�D���>.�7�!b9��]�p�E}�������KG�ϼ��aQ�>/�Ȓ���3kBSqG�~D�7����#^8����+*�E�X�74��y�ް���R�~�?�?Wˈ�k�� ����`��LG�*�ԕd��!�@��Q�Ç*�Y'bL6J�l=s��N��K�����6_�}�2%����`��]�^�)d��Őu�dc����v���}�tJkl�+�/�~�����-^q1U:�m#,�ޠ�O(�sb��a|�����<���eGDt_4�]�~�sW#����n=�x4������ߢI�%k�c><|���ƽ*Z�� �c�@A��ʌ���� �	�D_�B^~Lkai���Lvܠ��I�F�}���HL��1�{rq�V
; 3ضSb�c��o�@	�GgsN�@��q{ګ�&(�UO�ǩ�_���C������cպ�x��@�:�^��u�9���ڧ��90s".*Ǹgj�&�c{͢�6�T)h��.Q���*g���ɫN���F�A��&Hp�``>Q+�.���c#t�u-��Pu�E���}n�q�y� T=@�5�����P�G��0ݑSGD5"���Y�9������TO�3	��}�6��!�`�TA�@ �7 �_�9�)�6܍��iⓕp���^��Y|5ٺ-���2+^���؄2^���P)b�)C��T_�L�F�Qm`��7����T�42���:��Wn���SR�Y��#�M=��O'�/G#ulWB�9���y�т���0n��g���läﯕ������V��Ee�I�A�����M�Z6_�ZYSa<D�����<�.X1-`C�U��D�(�'���Z'��a�q?jwQ+���R�Wޤ�<	�hVY^��p<PX��lj�I�yJ,[;p =Co㦽�;vR��L��}�E��@��xL���Q,��� �E�s?eL��ܾ3Jb��j������K�KA�h[��Y�~��1�~�#�iʒM��]K������^�}�.�B��HeB>7�]TC�;!�D��y���r�
�^m��W�ǈ/ߊ�o�u���E]Ջ�p�g)�J�@��T�����V�YY��^4Ԉo�ܚ>7}����8k?�N8������ݦ���ʧE������MMn0��P��Q�|�W>���.��ΰ��n�2Z�� �n5��իˍ3�� iFtM��;Y�m��PI�O��b,�O��
sA�v�}H��_��)��0�6D�T7&t��O��$�2z4��5>���0���u��X�N������T_dΖDzٷ�J_���5��`���G*�0�!X ���OA[��Z�4g��x�%��@�q�+�~��^�@�VQ~��Y���e�2��h�  �)�`��{�2LY}�����6- %p�a�?��Me�+�Av!��W�K+Q
���7Ս����'�$n�Gz��LS'��8O��g�o��5A@�G�}.�b�[�M�pY�*w�9Ijd�&<�Z��ŸR�4�o4�VH���̵"Fiݩ�mA>�v(>�����e�4$�%g)�1��	��h�w���è��i���k�'������a�����+bC�ZO&AU�cj~S�[Cت+ɖ�8^uʌ)����//��5&0I� ����T)5���C^�q?�_�JT���WN0��1%���oSYir�/V1��Ve^q_���Ë�q�gAko�}�1{�D���IvKo�"iK�rTXW�_7��Zz�CI u�p���qJ8��w�d�o)|`\3d�q��o�E����\�i��\��7���T�b��D�/HT�6{ݿx;�dx��E�*l˦�%Vw縿ct."p�ZP�~�r����� ��W0B��[q5�q�*	��W��<��bZ��ǰ)<�K F��|��rN�2Z�4����]�~3�
\0�<����bd��:F1_���,��_O���}�Jm�ւ���N
��r/�5ГCV]�-QF�[#�!0I�r�e����px�@��w�c�l�<;�M�dz�+�(ax͘#B��ѵ��u��aG�T����C��4���Tz�4x�^m���<߸�h6�}
��u���[��Xx]Mh]ӛ����A�[�uE���Lλ2�_':�&G[ۯZ�XLB���dZ`L~�
�.v�fGz��0��Ї�8��3�yOT����%7J%�#+��%�	��9sr;�#jŀRю�UK���&�QY��fkQ��e������#�ɠoVs�KW}���A�[1�X�8��:��U�d�*��\���=�KC���'�u˽���ӲA��Pa�v�2R�CȇDX�nꑪahRu��ӕ��(.�OPsZy��wix(�+jr�?�_��R���w�5�m �#�_�z4�P�W�o/ᥢ�Tڶ���/�,���$�ta*n�@�+ϣ֥�X}�+
 ��ƌm#/��&�RT|pM��s��wB=��������ă\�L��Gg���[C������EX��=Ulh�-eo�yV�bn=�^�j���ݝ{�g�T��V@k���}R��t²�?Q���t^V�!�o���?=�����e�Ua���^�ve�R,��l���&��(�tJ("�0���)������k�v�I6\�L\a{�)���ڰ�E�}?a�lпRk�
3~���6�����8���(�4i+6pwӬf��\q� ۬͠L�'k���n��'T)9��ן������Z{�&+�-�П��)4��ş{X��*���!����B��U3 Ѧ>23F�� A8�'�I�I�!�� �����%�~�(:Jڻ
�4�j�u�3=14�=I���r�������B�~��"��d�J�x2�Їm}kY���I+�k��ػC��EiK|>֚�w�=[g��R<[B;�س�B.�Mo�!�P�;_t:.���R�F'�}�,4[����k��G^xx��,����b�$�J�D��1��Qe��|����0lFt˗KO)��e��0�]5��������=�$Ȼ�ͣ� �f�����\��w���k�xg���+�~�WYyQ��r�����(@Ȥ��Lf��Ԩ �$]p����ă�ҹ�N�T�q������A��-�R�	�?����t]W�v��a�R�Y1�u�]�����'�<�T@�C�(WQ�k������ǌw�P�C�_�!��fޛ�ٙ���r1�,(|�݇���U�|��]�ښ�r?�X;�e�H_5	�Y�דl��p���( �F.濹9R�6Ą��ŝ��\<4�@�Ǆ�^��u؃��(��fq-P5�7@�m;o�&B/e1,ä_��R�L���&=s�1�[�0*��a%!.��s�f��?�&�89�uS�4��/�g�mg؟0tC��~�H�Q/,�P�7�6���}7e�+���D�<0z=/}�x^&���6�~g+�6���E�E{�+ m5⊙�{ȧ?s��r����w��t�v����윇�婤����Œ{t�Xs�B]�����]��_�HBI�,h�@��
�i7
��j�H;��ސ�75�)6�c9{�HT���~��
�=�婆���Iy�5�c���璳3�����עa&FRd��1��-�U����z����� xP���߶.��>bd4(��̦��I������������b,1�A w��^�Q��r��C:O����Fp���)�fj��D�v������7�4�$����@�ޢ���F[���GK�e�b�+��?���޺��kA�j��P�T�np���W{B��	$�j�a��k��N�{�� ���i\
x�,��ΟЅʋ�9T�s�G������*a���� �
�}�0��݌�w�R1&��=�)#ѳ��d+�~�- ºu�cEhYr!���
�i���!J~g�J��$��h�]�[�~�E�3 �"_�c��Ʃl:r;N� ��aNQU��|�@o���N�m��_�RX��n��-|��!i��֭5I�Gc8J�d�_�sZ�A0�.�<	2�äߞ�܄���Y���x���m�4Ô4-qok_/�d��<�����g��'��� ��i�#�2�W��}�Ĺ���t.�;qo?f���.G0��C&�&�2&a��4��š�Y%!�vҶ��}�#�|J ���kh�z\G��Hd�g��C�d�7	�{x�n5ifĐ�#\wi�a|�C*n.n��m={b�0�M�s�p�~$n(����c�	�b�q��������I�=L�9n�m��-�UG��攰�s�1��a'�N���/}��|HWl��7�j��&��>���������ɃBw�.�,�·��� �|O�����j-w�A�L���*lK��������wϭyF۽K��75���@U������X�yi�������Y�$����g�{\�2��E^3c��<~9� �𡈅���'"���/)\;��jtӟ�缽�U[W�
���m�T:�V%��.�9`�X"�{�����Πw��~`@�풧D����Ux��I�ՋM{����E�ǖ���l�ߜ��DL>0��\g;���ߦnT6�}t
*® �y�"Џ[��l�D�-s����Vv4Dp�^^ o{�t���J���宼v�+�e�C�ƋT�Iu7@;MJ�ZȈ��(pZS�Ȣ��;S1��I�*4|�Ei(�\�a'�GF��,ҥ�h�ytk�y�c��C��
%B�T|�-HD�o�X7�������z�P$sq��RCQ�"���'r��j]Y�����v�7a�)��qH:VZ7��H�KZ��G��ps3�[�����[��(TQo.Vמ\�P�tj�7���vY|1!M�m��r��sP��9%k�~n2�t�`E@O�C��T�U4���S��\uF8�#�A�ca[�G�ȏ�(v�͖��b=o����ބ/[��[,�N[^y��R�Y�l�q��7ȜyN�`�ڔ��ѣ �b�qT����{�l0lc��J�G���7�%�U��:$M}2T�X��|��G
����n��m{�U���i�������ne�� �W�2%���6�'��KE
�d���%�L�����zJ�>qMÔ4g8�dl܍E�1|t�<)�O �����@����bW�Û=:�-`]et����72~*��}�zB������e��n��f���q�U%y9������� �Sΐ0B�A:��;a�y_F�1�@#^�m̾<�0���yǣ!t��˷&B��R��]P�:��w�$�F|&�x-3v�:���p!�!��K3�S-rQz�G/K�}��@7T�j�>��Y.+dg6$l6�BB�H>vv��^ɍ�<U�4���NV=_1�1��C��J�Ps*�
{<�WJ} ��vd�<���(N9tV�K/��>�H,��q��_e{�Cn�jJF�\��UG�u��l�vDCL0]�2M[��P����K=x��^gN�V��o���M�XI�ϑ����?DS[�7��u�޾�����H������<Z���g1��x��0��ۙC~���<U�]b���dC�`[)z����`�d9��
,\;�b����gc��6G	?!l��x�_ K�Ŏ��'���;�_����f�8���,~����z���q�F8�`��5�ZV� �	�WX�h�É��F�
"�Xq�z��R�J*7~=��(�ǈ}y�=)⭱�Drm�)-�i.ɟ�6������+�ͬS9�}D�O,`�EV�~�3]-P�(N��t����G��At��נ_��0ֲ	�f���t+��{��"9*�Z�d�*�Zrx��\D��#[�yf+i����؊��ku����� �*x����U_��Q:?`� %�ky�CPE:&��� �E��}[����r�6&�a��O�W�᲍�C/1�w��D��b.�(#���ǻvar�*���A8��M|h!�3L��>D_jV;�jܦ;ʀ�lY��M�-������v+"dW]ɥw���ٷ6�؈n�:7�X�=�_��i��Kg�/��\�hB	���Jrl�g����Z.��TV�4�����5��n�S�����FE�^�^�crV���*Iq/	���u>��Y�eKE�!·�ߞ�r�0�A�Ƚ�ڎ�xu�ua߯Y2f2~�밴Q\���?j)5a��u"��R��Q�pXa���3��-W8Z�,-5"@�i5���Н�O� �"t�m{s�xLfV�A��}8����:+�,�OrW�	��{ذ�|G�%�ǀs�Ĩd�
����^ U�&[n���ʘ1pג\�!��[/��q�z	@����P ������}�-J�@�Km�N�w�\
Q$5�j���
x�O K�(�pR/~�d�]�F��+ʁ�ٴO��+9�#�ӫ{��Q�'gX�?j7�B	c6Cn}?(%S���"�\p��$O&*a�ֲ�t��΂������	|�c"�Lt2*�+���x����y�h��1c9�׳�;()C����yn�S+8�^�(����k}�gs�<�lb2�Ap�n���l�X����= s���Ǭ�"������65X�J}��/�2�:M��^�%�E��	�]�D&�Uc�%ș��%W��/�J0�M0�݋�|�=��B���;� �Y���1|ʃ��:�N¹��V{f��z��B�tԔ�[6~:��u?(�o�O��~*�ϧ�v��m(�NU���T�^�@�dg�p�����2��V�a��N|��P�~5/�S!̔T6�x�XV��7��y'rJp��8s�����%����:�N-�h���0��-��qz����FA�9����k��8��uA�����:����[Ǌc��f��e��Ky�nqEK�b���"��sb�/)Ѧ�d�8~%�c�h2ܜdP tt+"�
�I�� ֒V��m(ޞ��B2��y��6sg�YZC�[��o+���F��:D��09Yɔ�ǔ�<�D�BNC�y�����l"fOL�}u3�K�/p�#H6r�$l�?)���]�����y�HJ��?n���"PA�=B�ⴞ��9_?�B:64�K�y��NY&F&��EI����a~��N/l�u��t6u����T�	j˨Ʀ���!��o���s����+Cz-��*�l�"յ~4�n�fN��ʌ%{G���<�"��w6��iS���_!���c�}��Lz�`�AӉ݆&F�6��P�:��4aQ6�ڛ �,1��Z����O�"!�(�N��mgmy'�3R�%�}�>�f'��NG�e�K���)lwPig2���������*���N
_Ч