��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�@��x��QZH!/h�0��i'�M*bH�	��#��V:�b�dR�\YŢHq�ث�gHgG��N�6��&Tz �J�t�����13��T�>P�w��b ������o��γ�y�;�����;�A��ćV˴��1�"�8��u�K^���V>��
N\��Xy\5��=N�{Ώ[r(73F:���+��G�>�cFt�t{�
詢:�>��u>!:��k�e��w�@���&�(�^�i����'�-q�v[�,���تxr�}�+�T����G���k�d��;+6a�^��t���j0u�Ŋ@��qc� Ȧk�Ƴ��><!�\�Җ�����Y �`UmA�D�3�Ȍ������;�jeW�,�e6c�����>�yp
֐J��ο� I��ΙKCf��-��i��.��ʗ.O��s�8�dK�'2�+��Ɛ;!
n�	�~���Lp�Ѣ����-ϿW�)�ו[����_��O
SUĈ���u�1 ��3�8bε&�H�Tx����)�׆�-����E�FE�xQ�닁�n��'!�R���SЊ#b��ʧ�c�9�AB��x��G�H��(�)�i�8��Г���X���͙23L�Z���S�AHܓF3�M�t��'�ϐ
I�Mb#����q!��W�6�tz��@�3	0����Mg�jT�D
zgIC��<��r�0+r��=������:ç%�Ӽ�ϲ��g��_�XI.� ���GزΊ.\�	��*c��Q�?�-��;5}:��[A�_�C6X���?�l(XW��M<�u�G���/@=ڗ�F-���J=�i�`�]�6�]�Hc��W�[	�%�Mj]$H��K����wqڧ�ς(��L_��8�$ �Z�$�d	�k��_ѥ�*�S�z����C�6�@��,�8�=��r�;@\lVФ�]�����g�LϖY3����f��|!��Pf�J��<`�Q�ov�D�Y�vO�_�û���SuD$:q��A*{�^������P���vj����u�^>��,Dȉ��{���ˀ4Ã>�HĞ�z��H���Q�9yŮ�.���i�i͹���:�k�0��)�(�����q�$�ʤ�^d΁���$�x�s��ܷt�>�BP�����8NJ��H�[�T�U#��iR�b2P"�Z��X�����h�^ ��kH�"�rspq�X�h�0�pPt�i��aflޅ@�;�B+8Oӭ�S#:�,����v�aK_�B�x�Ԕ)��ӊ�ת��$e��g�,�?�y?��)�l��e��t�1`�<��L���%)���⮥o.~l�����)�K@��[�{{�TUJ �)&����=� �P3���
���љP�q:��m�Aȋ"t�rl.H��!�B���V"�����=���n?&��J���oT�T�u�+9mD���pG*�_��(�P�;/�v����Y�
W��߯l$�y��(�/���f/�S�]���b5����q>���7E��k4��t�d.L �a�_�M�T]�`�J�G��3��VA^��D�j�;*/��
��d�+P�����uޜҹ��A[�[֩���h1�����⍛�X`H�::�3f�r��q%���r։��o��çֿN��P��p�MA������*�9�@�o������D@�;�3$I���؉�. cMҽ��@k�J7Mq)��ѹ8��)��!��MHks[�o���V��|Piޣ��*	�k���xu��!����W��jJ_9��픶���Y�q�H~&��<�h2�~�g/X��-#Ff=�<����X�}��awv|�mO��5���Y�/I<�a���J2�eM�̂�q��<�Ʃ�T%!��7|�FlTg".O%��n�5�U���{�]�ń�~OzA=��Da]�\��ACL�>��ڼ|���
4�X�C��B�e����ĉ|՗��o�y���pw[��6]6�Ǧ̀N}*��K	�]�_a�Q0�tbU棠��#;?ղ����]���;<��஦���FTK�7��	�'���&�n�q�wV��^��VF�"��)H��&�.���?Q��n���B�B�q�y�˻�٢k,,�������<�73��	�F(�j�ҧQ�vU̕������WA�,q�M�iL�g.��HiER�h�AԶ�����3�\&����F>|� 4K	��4Fܑ}c;�hi�Rh�T ���u[�:��\TT��g�.�]���0�S_Pf���I���k�}�S%{�?l��M�#�g��\�O�:R1|��+J��3�k�t��6$����#tȸY3�5�H#^hJ�<C¨�P]�
����}�v���yJ�C>:�Uu%<1y��ᑁp {p��;�hH�fR��%̺QXy�.��� }
6�'�4���Z������U�h�0��t���sNG�x.?ݙ	�2��h����sq��?֒O�[ǼI�~F�_�7�4Jb�gW��M02sx;�Oh�ӳ����+m+��-N*1\ ^� ���%$����'g*��O��$/0���t���$ r��g5&JVr���F+n ��[�t��8�Y��{���Ϛ�S�CBTX�as�v;�����6'�{�R��� ��5>#Ñ�1����zi&���y����f~C���	 �	���;���9��Z;{ ���z�A��tZ�w�2+EN?xʄzA��`۽4�"-��t�'�	u�A��A��M�(���D��w� �"H�z@�id�`<��vjSlr���z�5�8!O��<���0�����s��r��z.�!��a��|I!�.v�_�M>g�?s�J	ﭞ7�g�[����Yd��E)��5l��%�7�
�������o�:`�����yXj�B)��;s_����Ć$&JX�N�ۋu�]��-M�w��ɗ ��WZp�ם[O�T78{GB��G�*��?�j(uħ^�r�=Y�Ǖ�^5O��>.�O����e�gR-�]J��pl�z&�X�t�\�\�K ������)��#9�.5�ԟ�B�=����q���T��"~fU�|Q7M^]�-��I����l���oفt0�xA-y@m�Ӻ����%�o�[S�~<K�To`l��k��}b�"o����{�sH2կ:���?�sbij��E���|�:�<�8ծ��FbC՘q
��	r?�i��u���evH �|=����Ơg���Q��x��uM(�Dv�?[�'?.թ����Zg�vS�孟P�٘���Q �"��\���U&5,�vXz���Jt��I�S��<:9Ѥ�k�T��]+ۑ��b���D�,�u��E3�T#�D��R��I�[��Q�x����G���V_�d��j&�{q#�C��!�j����~�)OG����&����ZL�D�m�ÚW��V�~�L4�V��7����x��M t����g���o�ꮪ�������n�E@�j��H�~n'��I��ر2��Xs���V��k�� �k{îB��Z@|x�w9���Y����AU�n��ɗ��N,��븐�e�sƶa/����[T+�knI������	4��?����[�2��nx�{]���Q[iC|I&��H�Ͼ�ߟaV�h�����w�+T��d�IV�΍j��P������/�?��Z���&[
}��D,�d]�S���_�?鴹Y-Qsa�ׄ�*�_�M'�D��A��z�ͼ��h�	)����̏�z�#��������~�9���_޲g�b��)L[���l��e�1= M���m�3FW_��2���W�������& ����B��y$6�{g�/.��~஌&���]�/l!�A"�a�Ae��� h�wāc>]p�5���؜;�Z��Tt��,�5l�0��_xʻY�9�bYW�O �����dK�`	/���a&b'�l�����a/�{���T:����T
\���/�|Sq�ctA����e e��;��Ki���7��ν9hw��[UBobnW�O�n���_��y� ��9B��)�4E�mA#��e�kHT�^4�G$92�(�yH�����}z�x��<��w������N�E$/
*I	������o?�����rP�ɰ���~��f�cK6��C&麢����ί�y����2֭���a�w�J�\���� �;P����eo�ڶ��hg�A��hY�rVYd�m�R
�E�V�X�}ek8D/T�kl�$=��ܣ�3�߅8y�\�ܮ�h�����#|QE�E�:d�4Ӑ����	?���i-��L���	;]��W�G&��(���� B���:GZ��2����}[8�9	�k��M���r�؁h�tG�d�0������`M��&������(����3D�a`��ԹǦ^�t�{V)�pզ(�H�uE��o������t��m�	�tk�a���f��׭ox�j��A������1Z�ї_�|��\�CE` A@,I���\��ɔ�1c�
5������ʌE��9��9yu+�n=�M��X�z=T#�W��8(�!��#��Iܽ���v�?�Hy���܎8��8�� y��qxt�n��م���(�"q
rɬ�ΊC
V����@�$G2Jń��/Wgk�����8�B�5E�|��]BLAǨ��h=�{�q@7� 戦�D��0�f�D�V[K87*����l�r�z^�=C�]��sc���� ��sm��WU��tv���8��V�@��q^��US�z��+�$	��ڊ (����,60��f�nCg�㜹��V����Yx%����ʈ�q�rA�+�5ɩ���*���0���� s��M0��P7e������d�_i��-�(D�
�{$�P~  ƽ�Ӡ��� �m��GM}���.p�L���^.���- 0*v���/Ͷ���t��:~�t��h��MY�������D�ȶ 6m����dϓ
Ù���3��0�K���PG*cS���
w��@���0�今�`9�U/�|�����0��9�˖�1G^3������c}��?䍠��~Y��̄�o�<}9ą��Cۨƣ>��L0��`�'L��oUΈ^a�Qq$4}��9����K��{��1�I���ߢA,Rκ9o��+靡�y�I#Lg&��⟧9��Ŭ��(��0�����Q�q���$+���x�Y#�dt�e��a��g iD���a����!l*E���C��f���P3��(5h�8j���x��u[�`R}t05&I4�.�Q���%i�Np/�R��|�޿n&Y|�kt�Oh�m�6�4��D�.�i�l��E��8t��I4	�ZɌ�A/M���S�Lw�G{Z/��3�����d�������
�Y�怍�b��F�Q��~���s�������a|�
�v)Z��o�Y7ف	��-1�TRd]�u�&f%�52����4��0�ȑuM����BV۩�*{{��>�H�^Ͽ\ᓰP,h�M{��S�,:2�W�?Qn�k�S��P	ƳV�"�7��/��%����o͹p�/�"��c��F����B�̘4E�F�&�ź�8;��O�%2oU����%��Q9�r�����%1�S��Z��b�����f�)��OS"�X�5K��@ɸO�"��/�UB"
�WP��$�
A3��� >&���[��(��G����N�5 +���v{��y�D��5&Zwd���~��� 9��g�C�Jz?K@Do#w*ͩ���.~D�Ϗ�8s�*c/�����Y��z�3���Y@���)�>0Ճ�ݔX�|d
�Z�N�=�1��ա,�זk�Lƶu�uh��s/?�x��^C�Z�l��տ�u�|��ׄi;N�O4���I 7�ujŬhtO����5�g>ZS�zm�#��fVn�y��k�ղ����P��'�����>G;Sg�HX$fނ���[�57��(�_��,Q[C���S\�ި{h�$��ޑSŢ�����Ƶڻ�_�hf�Z,����aB� ��< ��gm{q���Cg{��7���l�E}"�<��<���E6N� |71w]��)f��
1�=}�G<E�6.�4���|��(~}D2 �q�����|�SfTigb���>İ�a�]@r�yس3�F\��^��)���A>fGQ�UɎ�7�B�+��I���S@ƍ�7�i�"]pPjtG/Ƽ��e]\)���I�C=�gIw�n�nA�`)��|gD�<�2^�[z��e��p��}�Sx��Y!���7�AR'���1R�]���P↊�Wh��y(/�*[`/��|{���S��=(s
�=������=5���PP��:���c^�ͩ�"8���՟=ؓ�I���♾wS��1h��������iP�̠��5����b�-��0NXx�đL�tUpa,�45�O����n���X�^���S��k�8���D� ��T��f�P�!2����9��E�4S��ފ�j��cz>2u�6�ʰ�!���M�B�/�@r`}�y~����,����dȟ����fj3��&G�s���_�(@�G�#�����!���{�v���6�%k}i����x#�;u�EEiC�X�z��`�A��ǜK)�8[���6�����EYp@tPS�&Ρ�d,�P�$��{�ػ���<��U��h,�d�W뤘{�a�_ʧ]�W��f<违
=7�sǑ��6r��J^�����h��i���u�/J���y��R	̛n�:�����`�8>�AAUs�����H���ؚ�����>�GzF��͟�kiOⱳ �v��T.��/X�@��]������v�NT�!r=} /1��ػ�bV�ld}%I׎���� 	bmy�y��%��S�^�l��Ġ6�w6��n~b�Ö$�&I�l/Y�����7���ܐ$��(us��	Sj��s�]Xӹ�&���E*��xs����C�鲔ã�N�/��h*�ފ��(��r��Jq�T�-u�Sn�՜Ib�N�y֙�����%)>xGy�i-�87�|�� �z\�7� cGC�׉Xץ ����Z4����B�֎��&)) �D-��i	+H^��\u��{��N���|q)��Ҳ�'�&3�|��f�DbHkg~/�M�I΄	2�Aiح�}XV�w36�~�Cq�4��p���t�R�p�Ѫn�|�+*�̡՜�+0�Bm"]�ᚐ�O�P-n�>D��h�Xg���_2Q�p<�����S�$�@˹)����}����ww�̜�)}*���&�bχ|S���4�2^���RX���"����.3(vH�P�5�fj�рsm��Z�L4��r�"]���k�m�QB|2��J���:��g��(��,�����z�r?�he��'�(O��8��F_]�9�}B�UC t�KnT��y��E��N�{X�� t��p�^`8�NR�S;��j��'@~��Vo���t���,n�\��&F���	`�ȍQU�ɮt�⩊5ib^��OM�P5�x�w�3��L�w�s&w�)�?�w�g�ȑ�̩s"��/��@�� NǍN����>���5r�as���~��1WOw��3����v]9��bih�]��ٜLo���1(��A�S�Ϙ�Xok���V�v�L4��{�hJ�bM�k��œ�j��\��p���2"����O��}Svo����v�g��F�bJɧ��@+n}ﵠT��l C<V�rG�s��jv���I��:͔(�U%�K�Tm�>��#�	Y��	����-�rx�~����m�!��4���+s���Y�}�q���NN���=�/n���q�p~�a�~ ��5m0X�K�0

~�����I����犫��=�L���g~���Љu�<b�H/��a1�A:H5p"��I`.No�0��3 J�J5�繴������)ٍ��pw�T�X�y���^H"Pa�%�o�ڑ�'�2>M�I51K�]ne4YV�������gFW��dn�"E�����6iR��Q~˭��0��d.ܼ�X�������S,A�9bE�k���C<�߇��eA����X�ad���++ܑ[�j����!�����{d��T�5ԣ� 57�m}��K2NZY����?��z+rc�m���G�����Ç&ߞVJ��dD8oD��	}�����q	���0�ăt���(�8�"�b����k��*6��A��Z"<��d��������R���`�����G]��< N���ԙ��3!����D�v��9E�V��:E�;s~m�f��e���.���!�,�~Ӧ�'��v�[5$CD��B�E��̂8:F��}~�eύ�@��RYm�ȳr���o�4�����hY�X�(cඒ��f^�ɛM?I$	C�5Q���ds��3�ځ	}����E�H���)ǰ���N���tdbo[!� X-�s�Y���sE����P�b�ق!����������W����i5�"U�x�F��b��6?��y�c�����0�[zEym�v�c�D�n�ż�g��~e
�vZq��
WO>��-`������7��\{B�k�ߍ����K�tq�e��p�m��_)�