��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ����Lr�q/���6�ƘɌ�eBS �:��yg�������,f��<~B��2�� 0���~��m_�P���g*E�%Հ�}�|�}�x�ʖžȠ1����1�&"PDH�5�({PX�9N���I�N��MJ�$�=�� ��k�x�)K�hs��F�T1ӣ�6	P��;��ȫ!I���և�;�@@ulS����Z`����2sdsJ��v��E����u� 鳗�@]R�>��D��wE�}gpS��4T��Y�^^�ڕ��;����Ǽ��;�YY�`]�!X���������]=;���<=� 稲���ܦ0��[@�'^�z�L��P��ȥX<"2�ކ����U����_��y������t_���v������1Ӫ��Wl5��$�4N�q�)Ҷ�e��Me�^a�Ɨ��@9y	����ִ=x�*���O:%��L(0!?���&=�)����$~���U۹�>4L��!9�|���م����#����6{U��Dɡ�Mbѕ��� ��5���"$�D�l���^�OjՏ����M�C������H�Ԗ&L��+i7�����Z���iL��lm��;U�matS�y~�ڈ�����ů�-�a�ڡ7qwT9Fp:��IxSČ�&�#:��q�Z�]Բ��V�������"Ӿ�m�Cj6�,�m�L}n�>�ΓI�\T�a%��VL8Zm�����8���xڅ݁�F!M�>��o�$YW�vPa���p�(�����<�1��"j�M��6�w���Ap�ݛ3�&Nx�PYO}_��Aq�h�-,,��&z �O���%ͅ޷�QQ�\*�1�?MCD�x* �+��L�F�+��!(�\5�Ͱ\��b���S���3��/[I�C�i*w�ր�{hqzXX��Wq�:�k.��&}!��2!�C�Dʞ���CZ%�<�t*o������O�/�Br,2���+������?����t�~t���] &g�k��K�i�~Z���ن�Ub8���De�BTK�k�G|����6��M��q%Si�w{��1�� �A"�?� ��=9�!(��~�����-�\>V�2��9I���P��%�fDv�Γ�r���]�.	�P��գ���>�,n_�zl�{h'?��bg[`%�R��7����[��]a��t�v�z��#�g�aeP��Ru���d��w1һ�M��f���"Є��Uƺ������hT�0�_��Όx!.���f;H��C	 '�hr�G-��,V(�4�}�?��[�ct�8�Ǜ;}��� �L0�4夋�u�)cRQ3��ՉdX)4BNn<c�B��*�1/��h��m�NQ�V����9���c�����k^xJڼAt��*����B�,��o����߱[5��������Ϝ|^�	س6�i|R�V�J�Z��,����7)ЏG�L��K��T���Ѿ��E��0tn7�cΓY�>zE2�� YOM[�R�: �d�}��g\@
=\s�����@>g�_����,��+p�/'�S�F��L��ϯ�V��ގ��r�Ŏt��p\��׿�=�����+�l��g���³c�m��C籴�W��O��#,m����q���"*��� K����Ҁ��FM[U=QV ʏ�'������,Sh�[i�H��b7	�	2��х�h��fSz�V�g5U�&��hǖ��⿼ ��de�a�?���3M��0�-/�.��v�?N����j׫��%��zM�e����t��T��r��*�i'/�	���rC���.��'?�G�@.@������w����ܵ�Lb7��N])Tb�z�6̰b�(�FwLd��w�ί�Z�\f� ~P'�ä˄F���{���b��K�
���V��f��nEJ�q�WF�Mt,*]2?����(x��h��	Ϋ�-8��Ŕ`J�p/�ؕ��W%PY�����H�sgU.E��SFzC��r��f��4>G�z�x�Zuay��B4m�9r���d�f�\Av���i̴z����O��|��?���d$�>m}fs"�����'� o��HX+�=�ao�g�˓#�W��f�)#�O��n�B6��Q~5JE�����Vv��1�U�і,+Ɔ�,�W��q23��S��l�9��`x�7H7��I)S��){���$�}#k�9{�pg��a�~F5���F����Y��¿��\�����Z?�f�&o7����L���P8.��_2�I��Z=�y���.3��@-U̹.Cwwh�4�E�W\��.Q�����e��X�PHK��b^W,�^�M�QW�j�KtҸ"&�tܫLk�"���=TZ���l`
0MH���+^'�����*x\\=���w��S�d`���A��A��`K��3�Ee�N&���ݘ�(�^D(��=�a�������j�I��T���6���A��L�	��J�6��"	3�GHN��#�z������ړ&�!���󝑶O��s�� ���gd�a�p}�e�gΐ�����c��A���fq�j3b�j�-��q�&��ǳ�Ƞ�D� B���>'o�u\i����6��˼�6o�+6�h��� ����b5�i�6���6
�Ƶ����\�����gp4�U���%UA6����_е��x�}:�T82�r�f�����*��Ə��6�b�ݾ��1��4y�W��rw��ŽKluI�����B��:6Y�����("��k)4R�21^f�fM��П�!����l��/�$̥�JR��������dz<�z�h�@����[Sp�Mq�/����9|M�P�z���o�h%��"���ϺJ����B�p`�\Q��CI���a�c�^;��~�$oНEe��"L
��K!%4)���,�7#��Y􈂖����%��#�����>͔�>��RF�z���v�f՝��������qk���9�N7��3���3U �g��%�%֏�j�5�VX��:8���p�4A�ߤ"n�NA���Kjv�zT~1Xc(k�� �!�"��Z���̦��n��K�.l,z��[��&_С�=_RfW�|��T�M%�$Ţva���|�ҝ�%:�@e������X��Y���ٶ���n*�L�4y�2ܐ����jw���2�y�"���J8����m�2�[�����Y���١8�#�Y{dڠ�^D�Q]��k�6�/X]�ڠ=$��j�a=��K!�{`�q����Ϭ>���W���a}Vuwg^9.i����Ǘ�����F��+�fU3���y�!B��:�R�Q�A�%�O�Q���E��K1<�}ץ$���2�?�}�1�Ư�q_c���q9�&�Wc%��L����Pp�<�A\�F�݋\	�
�9�x�U2���5|����&;�uc�
�.��]��R�1Y
��P�N��Py�D��R#���CN;V�+���l��u���wbi潽2�a�?�`�^�b�x���-�4�Z�;*�X0��~*����I 8���� *gA�G� B{��qFQ0e�{њ�J�/b��	��_�DE��s0�1؁7{7K�U)Wh���,�g��u��d��}E��o+N�da������p��`{�A�<Ȭ�J�"���ȝs��q���O�_�9V��MVZ^�u�E!��-�4Yp�)�9�������dR�	ρ��#9�H:��^�	DT7�|�>��`&x��y.�\�w�Zr��Ť��Ȃ�����g[�Vz�����D�@�h��Dh{�0P�Z=�D�=Y�7�?�<���Y�0O�IU���`�K,�&��@{%84Ǭ�m_�	L�z�ΜnQ�!�P��	
�G��\%K�=w�F{����NEy,r�؆03�|�cCz�ʣ�Y�v��)�s���:��#�0Mj��Fo����)�*p����=r.�F�ۼ]QB8��9�zq�#�:����t��n���:�ɩC�U�V�Rx�.�Ƣ?���.�	�FN�(�|���|:�����5X�Q����L%�A��;cj���}�[:ג�:���u�5��3[����n�=��B^u��ϼ�������vcMPq��Q���i�7��n�ԥ��^|j��I��
]v��i1��؛��X��g���@hM|F�j�H���K�+�~��t�Y	������J��lu����:�p����K��ŮF$[g�Z?T`�)&+�����ޜ�����~��by?���5Cxue���%�^�C�+nӪ:[��m�z����'���)_1>�ѹQ����P�=�.��RH^F�ތ9�!k����_L�L '3U����>�euS=��=*"�x��=2Y��� �d�ُ�e��fj���i��R��J dѳ��j#J�0�Q�����`�d���x�� 3.��E�?�S��꾐S4����FK\o�Ī���_�7��蠷Ɯs�Z�y�3����eq�N��/��_�c��3����\��1�TB��Љ$�3�{��H0훽-1r��p�n�.�fB��J��q«3ajJ�$��M���ֿ~�	�	
�xA��j`ӾF|�8�pkZa�eLu��?�^�{�P�2�V7��tDs��" �)��+ٰ`���YQ]շ
߁�ԫ�3ٙ��v0B��h�)&�KS[b5��vB�ʽ�i�YHL��-R�h~� �[ K#�=��Fы�fRn��kz!'q���b�>��*;*j:����+D�av4@U�>�+xA���K�|�����I/C;VԽhە�����D_��GP
���w��C�n�j��f��:����$[���X)8�X�wt���i�舮��"�,��P�����t��Vo*݈�鲉�1nj������毦B!XE�ML X���.;e偃�U�Y׻x���$=�Cd���{�$GP�bh�zX5ض���j��~����C�G���_;�C�Rxi)�v��	E5[$?���K}����/GF������!�U�����p`���5���1��5g�`S�ϝ&gO�+������ͧB�Jngm�^qc�����DI�bpTo2�,���9r�Ϋ�v��p�}ǒBD(���۫��l��$9�%�Uu[����=lh"zo�J\Q@���0+Қ����b��	+��4j$�P��˘�kk���$L�f�M��pѥ��A�ThɊq�x9��w��<�Q*GR���7O�OvQÏ�,DV����L<8>�z��&0K�hD�I<���[�Y&�B����Ǆ�H(i�	A�T���&&�Fs�_�xaL-߿��	���䃌â�:�H�ts�$�E����<�xtp���?b��ċv�x���U�k�+�9�D�@xڗ(y�ǅ9b�[A�X�Rw�� �H-��<���q�xy)OZ�>�5�I��]��<����:*���i'���Y���;�]!�>��Y�e����nn�v�Ay ��_R��{0�	���3-�ǰ[$����7M�o�(�	�1\��Jyl�P9�@�ϓ0�u�x�qYx{�`y�"4R� ��gp������=��w*�
�����MdY�e$��ăv!(����j?x������W�B�ְ�����;��]�da��p����Kw�D�4u�!�C��v�m��&�%Z�l�á�%�@Z'�����`�H�6ÜZ�_�ȊtQ�����a4�aۮ�\4�usM���i�8�y��f}���n��ʛ>pƸ<�#�!����g�>���h^���d�:I;��,I]٢�}<��wG�J�gICfO���]�T�yTw>�)fh1�EUq�:f�x�cC��EXc4���g�m�'0r�#�:�K�}Jɺ#]'H9�8��HQ�p�ȏ3���M�MU���ǡ{�ju]�u>�r��]D+��P[�v��߱i��m�������3K���Q��8����J9ҭ�o-=���`�7ǀ�
�L�Z�.�yFx��8k�g��O�XCWo��1��ܬ�Z䀒<Q$i�
!�<+��
d�S���u��$P�|�ܖ$i�t����;�+-�y"~*bSD*�`i9m�K5�C۸Cz`�f=UsR�O�e��+��p!$焑�-i��X�8Dv��շ��c�����C��M�[����[8w��ǻ�..=�K�䞢C�YY�$��[2����?S����l&�Z�o��
f1��R��b:|���Ѷo�����2�P��ww�ڸ���o/���+�	c`z�7KrĨ����~re0c����8%����L�o��}����ǀ�}��4*����GS��@:��[��ߒBelrS�-����*���M����_�{zl�t�*.�{q����kyٸ�������/Oڻ3��>�	4�bl:����9��NI)F�P��cob���$2O%2U0�F��H�"(2 b	�l�l� gdŴs�Sڎ���p�5VY`M�:�D����ɧ_�^F�Q�3��׮�B(�e��*���*n>%�/H�i�I4Rf�s;����t!HF6F�P$�<����`����~����l�_}u['Z�ƈ��U�� L�꘮A���]Fzs	��_����n�U�əI�f����-�T��ZG�R�.j>;���!՘��fc�>֛��ꋊ�` �t�˙��6���'�ABƿWQ��v F|%:"�`,���-pn���U����"=7������-̴� (a�� ?�
��xY�+�^]�0b'�0���m�u�0�"Iu�~ฏho7��̡�����<��ɨ[[4�l��wdl��!;B!q\b���Ѓ�c��QB}�`U(!�q�#Cj�� A���2j���%����Ce�	���@�\���Ԋe+a�����b��=Φ��%�>s#�rw�t4(`�j|��"�5����=�)���$9�GI���m�^�<�LwR�6�1���e���83Td�����n�MZ� ъUzdtL��I	�?�eKq����ـG���B��J����yW��Jބ���Z�*�sor�t���c�`��>uS�B*Bg���*�(JѰ'����;���7�AxtI�u��ś�%!�������?���)��:�;=�HmC*��!4m�M�K8�R+��fF�#���y;~y�����i�^���޷�J��Dۀ%�G������-���x$���=e1����*�'APd�JФ��~4�%�����3��J�:�>nJY�?L���BP���c1u9"uj@D�2%X�s��§t��x�F��iPbYf����#X�,�9�{�������򟚎C���TA�u��F�:�ج ��m��&��I�!��!M1��+�-}�����*=u,���-����ɲ�m�=U�8ӡq�?�����ɏ����O��#��b(-U0��d2�{B�Jy��	�eu�p��ɸ��I�_������8�T��9��ww������Eɇ2,��q����u�NR��m�L�����\��f$E�������L�.�Y��;�*>o�$�WIƨt�1o��Ynh#l�*��9M5����\e�չ��G�&Z�qV'>��(�9���/��0[�j�,�ci��1?�E���z�9ծc�R U
p�߶#1�v����1��m����0-����"�*g�C-��D�"/&�r�e�<	M��8�"1��*S�������T�8ȗ~x�<�vjY/���r���E>�H�6�s䈶��Qj3�K*�*�·7��$~�>����d@��v֪�9�*����Z;cuЙ���s���z�s������U���Fz��(4��I� (>�>��{��%uL�t��*[7��a��,�՜lYRѳnQ���W�oMm��5�����Ϝ.-���/$�"ک��_YB@�M�M����\���hϏPʁl�W-� ]������dHA�+tI�w���v��e-�����~��õ�I�@�ڳ��tdK@���R�lihf�����Zt��M��SZn	Z�?X(����S������,#�i�" �%��D���|��Ĺ�|R{��E�ͽ�D�n����\#}<&5�0,hJ.9�HXQ�Q[�v����X�'��53���K�����!�^�f���фGй1�AZ��ʴ�F��4���� H��y-m����q{ȍ��_���A\"i���qb-��鬒м ;(K�NZ�v�����Hb[�;��j %��z�"��TF�kd�s�lѐCAʔ�p��X&��a�����-�Q0�Fg��=��t��J�a�`y�1��ĝ�0x�c��U�5�So�R��K�(���ߏĺ�x�4�	B=�r�,���>� 
�?-ܟ�8���f��2"�0a���>��U �r�A� T�Y���O%����^�� �J���'��}��I^]`w[�<�$ř�������Bi	B�Q	��1&��MB'^O�<HK&��I\�9#�<j�^��(�s�79�x���􃷦���*2��z��x+��V�9$��㌣�d�'�o�rB[�~MA���z�;�����u.��i�|h��r�9ޠ�ܜ�O�yK��K�S���q{�#���c�ž�v\�y��M�7�� � ��g��pv���K�j;�|q��O���x��^�<�	
X�j&l�2
���]0�����K�&��"v�e�V�<ڊw���Ӛ��@a���\GA���(�+{�S�zY1U9{�9/K��?��c�<��:��ƬP�F�6C5���UD��y|���g��ueC|�oN�q�ta9�%��v�3��;f�V�xmUy�Z7���I%�o�Ƞk�B`�GKc�!���Ƨ�C5J��Py�k�ݸ~]�����E�����DD����X,���Z���ܱf�Fͺ}��r5�1�IAO�Sw'�I׊�a�KE��
�l�>��PHA���ӧ}�Cl����,u@���&CL�x>��C՘�ڏ��y9����s4�x2�$����l3�ک�e���Ԃ稚�&�L�~S��\F�~9��u���$O���:k0��8�I������!�L����b��caF�
*�⊕��hj��{c�ˀ5B�0�|�m�7�4�,F6�y�N��r☴�AhU{�&@[t⟻�����<&��Z>�;dqLcp�.���5$��E�O������A��@C��I��u�e� �Gx`O����a��ǕS�V�V��_jQª��Ie���
�mA���K#N���C���A�T]S�������7M�R&p�M�Fȟ$�#T�X:2���<~��׿�^��Q���c�³bD��XJ!�+	�G賚�Y�+��9 �x?�z��ߟgWޘTH�df��[cd��L��w0�\{��}+��ۜb����K���di�뇐�9���9��L���X4����uBu��d\�v��������|D�R��D3�'"��Do.A���	�������܆�Mׯ��VҳN�'��Ԥ��J]��N"�^L@�����tx�?ͅ�)2H�OY�h��gB5�6�2'eް9x���<u���s?���ĢL��3ldI2�O� LS�L3�e��R�Z�%�!��J���
�*^^�$k�R���~��6�	K2�r�y��D2gx
Ӷ�T�!Ţ%�^e��mp�7kK�n Tt��/�cw#��c6&ل�P-�����[��K�/A���݉�/B���Y�k����8$-O���Ñ8S�9���h�3GIc]���<�\"�EX�� e
ʴw�e_D]q���QbKBnX�F��{21�
����8.���c�I4�z}=[E������D�[�tv��n��\�Mˈ����.�FW���fr�a�����d�s%�׸'���&Sr��$(?[�'��T�5�h@�ⵤ%"J��ځh����څL78�X����x���u���!JF<ݷ%'0��Z@܇�0q�s��ȏ�ɥ���	��"4.j�h8�#��r�g�Mq�:9�IyB�(���m5�L߷�?i�՚y��i[�o{b�Q"����H愔�PB"ID�'i�2 ,���:{:q%n�D-��V8���/����L�Ml�	BR
��(�.wMb�g��V��f�Y�q���,�+]��rd�V�T����a)F���{H���+�O=�i[Z.uPz���6��$P��J�X� ��C:��	�� $n:{LPN��<]k����+$��+�&����YN�?���E,��Sz�ּ��y�~�����@���Sm��!��|��[Vo��4�B��w�fx��J���k{-��.q�#]Z?->j�q�vش��CaѪ2�\$��Tʶ&����]�|!D#lbH�N���]C�W�
�x<�5��~�mo(ݕ���C���k��..���g	�M#�2��B�P�f�� ��Nxá�P�-J����e
��t�ŋ5�x��t�
q�n�i}v(D��.$^�:�(7�>�؆�Bb���ځ�B���LJ��?}i:��+ܷ���[��x�`$F�� �!$��eU-2k�
���{���vM��o$���SX�m���=JDۅe]B-���(������ �"���`�qJY�助�����`}��,�� �_)$��l�W�Qw�I�Mu�d4U�Fbą@������b�->B�H"p"J��C�,0I^[֭̋��c��}�'ѸjX�O��ĥr�rg��}��`ߊ_���t�x�)�+k���܇��$Nj&�����Zm�s7薿����6���&ՒCp?�U��)X�^q`c�,��E3�b�|j����;"�����$U$x������i���K����� ��8���[==�zR+_`QM7�3b� ��F�Yxy�x|-���h�3ʄa,kp���2���gZ��Av�>��-�^2u���;}��#�S��J526��Z�&}Zg�M�2��1:���R�>�Cu61����4����̾1ĽܐWC�L����^��t���I��?/l6��ݗ���r���m�i�^�q, z7Gگ~�O5�{��\)&�A��ۮ_��憔�|���@��)!r*��;���\�^�&�[��sz�����@��������CO8�w�a�)IIy �<lGW����c�c|b��^O�ۯ��p�<�S�i��e�ʀ�\�����W�
[Qˇ�2��X<wI�Ԟ�Y��@���@�B�_o�6���w�5�(�m���,pb��Am����A�N.;��3�������'�-8�`�&��Տ~[ V��`��$��۸��o���o5~0����E��i�g�q�Ġ̏_�����RA���f2�$�fR��E��	�Cw4P�<�2��}�ɫ�U�Z� �=�$�˟�z�^���s0悇L�����3H�0\ټ�Ԓ�l/qV(����}7fP�o�{�k?`���c?�����g�V8�k���{9+z1@^�[WS��f %Y��
�,X0ٟ	�,����!B�Y;J����D��bgGʬ؎��Z��