��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk�㣃���z�Y��G8�SB��@��<Z��^�C��R�=�};Tv ��Gh>�vc!���	l(�ߌ�,���R��G,V&q�mvJG|�:/II�pu�R3q9�1��q8LLyW��kq ��K�֯�s�S6+�$_ƨɅO���G�D��Y�T �-FS~�Je��
�.�d��h��EQ;`�O���Ԍ�#��?�nѕ�t�q��2���՜)*ҋ�	����(7�4SbkH�w:��w�O83��Y���+��&ŃN9��&VQ�y���H���7�R�������@av7��(d@���O8��cgN�,*'���̣��i&ź#�ҹ՝
֖�2�"����z Z��G)s>��Ew)3�F.�Vr&O�u�*E��t��V�P��� mG��5g���!>����~V��ٔג�@L�7�+���ܬ�M��*&T��{�y����΋�4�B_6���:�%5p�h��n��Wm�@ǪܟXH����]mݮ>�d�"鬔hHF�mk71$_�볒�8�1�o7X�5���4�+��¿�C2ˣ�}��]��J3��dY�.'���Ow$gS2�k��N��g.8B+�*]}f�N.��크��ꖼ}�$�5tS��s4���-ET�|�n�S�m<���O(�R�0�R��Qk�2waD:F�tƙK�oE ��>�8�4����2�9�&IZs�֓���o��'���Vy��{D4N�7�F)m�+�^O���#I�Tb�y�ɿRS"�Hr��]����qc�AEgM�pWi)+����J�rߒ�\ڥ�%FI�K6�;�(�ۇ�K�o��������G2n|��ݦ+����-a>�V�g�eT�此-��ǲnX�K/��`l�V���|��Q��0?�zK���t�B��:s~�Y���J�|�]�R$�a�]>��^��D���(M�|�<�0�؋z/�بu��7)�-���T�y�;���
88�.���� j�)��>�<΢�b��ǐ��1�����%z��ar�k$B�%;�u��O)k�'�}�9ÙӸՍ�&̵gK�V$���!�s[�o,Dt�0��M�+U���2�+O��k�1�uX-RQ��s�8�!6�r�tB��o�0t�����+�Q�F�3� ��=I��#��_��3��q�u[��ML+q48u�	b��u�lj)qZ����?�!��� 3dcq;/�9+X�b���#�J����#�.�cN���q�O�x�q{�0�o4�T��� �����m�m�6 ,�>�d����͸~��3?��7�Zּ !ɱ,��t@l�e\����r�y��H����'[p�3�ehwX�/_��J�q&�>:�Y�{�VI�4�� QFtGpf/�E��5.��=6>t�u�3R1O.�F
�s�S��/`L�#H��!�q2��Ҡ�B56|�+��	��%�w_���X�_]A[����נ�i�L�q-3�da��t�n*�(���m�	�w�uwV�j��L�N���*�f|�1 (U�Q�ŊˤGRuJ�X`ϓ��\XH�m�.+������f�Ӏ���6"�#��@&0��:P͝����{�l
r�YM�}J�:a|�hUy߆�C�k����Vet�oCۄo�P����5I��P�c��-Կp{�+ǐ�,.@�PD��G'@�	�P��H���g.�r�96�1#���Ƣ?r�S]q3��5A]a(6���2��$�#��9I�:�G���C\1Lwț5��v�N���8�4bnҿ��c����މ���
ë�ۤ<�齒�
LD��;I̺k��ȩ2-2.�E�ڏ�����]�t�x�<���Z�����Ӎ�^�}�{���P(;����?��>��ca��%�?֤�Q#�K���^)�z��ї-�����S�_D�K~:���IZ����3��2��n�;/�ЅxJ�~"pύ�~D�Mh�ٰ�Ə]�q��7�&G��3��y$���H�C�y>�"ɢ�zW�]L���1�A��x�~�>�\�/���G�#�#F�8�΍�JU�@T��3���_W	`���93�#����I���8�+�����˨Dzi-Or�Ƞ���7����|A[H>:��^�%��n��9�q��'yǉ�_�[h�^L%�X�!�U�� yٓ�`LOgLūD:�=�D,��5��F� �؋�Hp���c�<Qz;>9�����������]n�����?�c�R���_��Q���������]��Vs1��ȏ��qP3}c���Ԩ�.%7�~,Yz���߂�A]^�܅�z�������Id��\ݮ��r���=���N8����Z�5]��qQS�3�����	sPh�΅,@h�؋KKֹ<��/R�5�~u���Ő��m���*�d��&��أ}���0Q	 ��"�<��}7�`����:�9co8�Zl��B�Kh�-�7VA��w�3��ne:� cX�6��F���'S��w���_�����`RDx F<�
F�M�`�Y��p�<�}��y�<��^uTf�'�ӥt��Mα[$�*�<o����-RC�[(��ꣲ�,8!<\�Y���ܤ���)�0���Oz^r�u,�XT��o�R4�@qh��ߘNP�!�Y�"�:)2�o8�� �%5�X��
~PǊ���غ?�N%_Q3�7R*Xi�~�}[���m�t�<���?�k6�n�P^�s���L��\��جyQ;M-�-@<�H���gtk�zv�+�K�&��n�.������vJ>Fr� V�\�����̧z�U_�iQ��YF��yb�.�diZ���f)��Ew^D 0�I#��q�>�%�}>�EM2�+���0�2��,��.�%���]��~R��$Vo��Kz���Lz4����~4k�"fV>G�^>p�a z@Q���}�Ƌ�`�u��NQ� z���S+ӿ���m.���|)K\[D����ŋ�q��#��bW���C_�S��/Ѿn��/���o )R �y��+��+�H�Re��h�\a�����m��DD���o��A�=���86M�$�}��&Ӫ�}�X�[�6��
H;D�:�P
FM������G�!����'=�,+�� �l� 4����
�o�6?zik(���s0�\�����u�7�ꀅ	� �H�j홿���x�-W�	�	.�l�5�$��k�鉼���&P�2=65�\�IȄ��a�\��k/����{-���P�yyF���
h#Ƭ !�(@I�#lU��
�HNJ�Ĵ�K	%�m�2�_V;PL����J��vdxw�(�ms�$],� U�du�W��b����'��.��\~�O�8|��B�y�ͺ��VX7J҆>şp8���Z�N�Hi[Uk'�����\?�MʜS;t�	��Z�-��"��� &����XE��N�4լ�+-q��.�p��<���h��݊on��2O��}�%)0���(͒�ͥ���T��u��Ώ��V�i)�"�T�i�M�Y�t�
��~���t`A=�K��<O0m�O]A�vE�P�	���Ӛ�浳^,S��;�45���QX<�'��d��%/Ժ/��E�uƪNau���q:�0���Ȗoz�aV"���b�ԋ�wp.���]��.!++ 59��T��4����J|7������t�(0u+Ĵ;'g��|
)�t�j��Zе��!jTZ[�|֩���	��"� L�+o�����|���v(��3Ki�kT SM�V�������;�u�F�TUV-��$�.�ݼ��'�U��	��V�W,��7S��i$���t"��懙�\��msgKe\
7C\�2^��|� +�)|��i���"�g� ep鰅e�$k��vM�#�PC�������C�y�Q%R5�0d,@�݁ �.��#���\�.K��
���L��@JX�Ⱦ�n�<���+��=[4����ip���6L�=N}�T���������v1��
x ��u��}�L��x�4�TԳ��v�z?��+@<�p�5ď�q���s�����ewgO�{�e���r1��TZ�e�kEi$�hr!l8�g{��~C��]�,G�-�ş`��K��?Ͼ��e�Qn������VW�FFg�F�A��}����ڑL{���[�Txt ��u���b��y婺�K�`o9�*Ξ�T��5��e�o!=	 �皎���߃�Z�Uʤ~%~��D���������d��VB�������?����RS�2R�rI=~<���P0���A�!xoҒ�4���MWEk9�`�X�M�����db`e�U���m�L��Zra����~�LҎb+�f��ʚC��?�	��%=�񒒵ټ�&�Ł}�{��A�Y�$�S+���[�fZ�$��w�')߈�E����ОU�߄rX���앛
G@���B���aܺ���Wڌ��o��wW{#��L�kw����E�'
,����M��T�!QF)	�S�N��Y<��������뇹��E���EM�i���;�s�:\~�����~�-�W����)�m2�@�t�h� �����t��q� ƾ�<nm i�$�� �mN˪�Nh������T��Njq{�Ŕ8͜�4���me�?Ǯ�UN#�&���U�߫����il4eG�6��.�('����C��_�e/��� � �q�-4||��|Z��}L��U�����a��%�R��G��G_���͙6�P��,�k�M׮�O�H'�DyQ*��+=QpH��^o߲�ri���u�ܫic�b��X���$⧢A��R�Z�WF9�8�nh�t�=�9����FZ���������9BT�����As�� ��-t�C&>��3< �9՗�z����B1����g���qZ�;��z��3�Yu!�����6b�c�����K��<��1�����.�?��-�,u���J�D�ւ)�f�i`õ�5�}�Ir"���"?	M{��Y�|1�潨㲛��m�Q��!\4w��n?���&n2��R,����L�5��U��fS�ڈ�q��^��P �y��l]p|�+{��ǩ�p�S�3r}ϻ��<�q�&��E�Ч��+vI���6���'}"_�IL5t���R�k�s���^^��@6$++�����D��TK4-���*�"��#c��̳�<��[�D�';K�+C
�f������D�2�6U�Z���ej��V=�{�˟#��=5]��n�&�Sw����n�$,�t�~Y����oA���rּ�
�����]ʹ(N��p��h�*��U�iS��-Y2���]�ȣ��_w�O	�r�ppY�:�9�q�O����6������8���6�h�_���8ۿ\5��66I�� ӿQ/sf]���K����������_�vߕ݇2���������5�ʒ�O��ʕ?:��*���h�f
� B��!�t9�Dg��*i��Q�ޛ�j�`�sgW)�F�f�O�2���u�cW�M�u�n�I�s'P��>U�ȴ�!�|���L (�E�_2[�Ê$x-v>��'$�ͪ=fKgSF�`L
'�j?ڶ�P�:�*�Cs׃XqA�����`f���B��~)��ab[9��'H��s�����W���LwM�|���΢�ȏۅ�UD9����ʘ������_���x�N�ky�u�U�ɝ��v��R�q�MqZ��`��w����ֲB]�-�Z�O'�4��h��ˌ�+9��ۄ!��ynJ���G�|iP� ��9a�e�4�G�*���rJ�P���KWP���QU�3P_���q��P��G�A7�쉡��׻!��`c�4lǢgZa�wk܄j��R�����@�q_$/S©��O{��߽���h�,�C���C�Yv���ү����bw�S_RXI-��Ö���g�y9p��'i���H��̿�3��
�>\_�~R�{��
���{b��Xu�WI�.�Z"�p� ��i�[���=@,�5�u3A䰷v�a}�t�jt������^�׺^l��	������������N30G4���n�xӛ���
� h���r��[�V��X��j����V"�9����nCg13��p����1�%����v�5RK��b�{����[գ[*e���Q֢X���������y���h #��McG��n�!��'�Z�}�T,[��@:�I���أo��Ea�V(�e�Cb����y������C~i�=`�ω
�LVX�Eܤ��]D��a&%���9tL'��L����¾R$�U�Aq���E�{]��y~��S2Yvֺ�<$�Bd$5�����Fz>�1���1�,P���v^ҷ��`X�מQ�=bQɔ��zdC��7�&i��E�L�公s�'{;2/�8�ɟ���̝Vϕ�6?`����!6�N��G?.A �6�xs��yE�W8qІ�����H�O�!��$�x��!&|QlP���q��e�|��%�8�G<����w-?'��\	fe� |ɽ��ʜV>�=:���.��b�%|�0��\і��+�8�T��@J��A����ہ3:��>p�Y�:�^^���m�+�X�L�X�
��>5�½2J�~94��>�I������2d�"���h���X�:��ǵ$���T�O���7iإ�Ux�)��A���!��9�m��}�h�^t���\���>����w�&�(��.RH��PZ:�y�"Z��n�CA�O����U�������;G����Q�
�u���I\7����k��$�P��B�E�l)�W����SZQ��l�w��߼\i+V�@Q*�~�����ڵ�Z'ge������+��2�e� L�Qlrj��ڛl^G~?Z���c�w��uW� J'ў�&�#'W���9���Ui��$,�")���@IQ<�*j�i�?Y���u6�%�L|w@��6�bD����_��m���}�ӻ�c�P�w��vo�݌�s)R/p�.$��D�f�#��&
ѵ��^��2��j���򤋮aQ���}�fO��[b��ьs&vs� �^%�8���"����)�~
M͖�����̥����4{_���|��)���z���(��:�L;YOb�q�Z�L3�O���\gJx�_�K�*�@[x�,m��bfI�%*I*��8�ʗ���jN����s��w�r�
�0bΦ�@f5�l��:0̔us#��3�a��αS����B�JJI�)�P���Wň0v���6���N�T�3�gk�C�J����=4|��-��������n��;7pd>�B��4��q�TN��BY�
wW�On�����.�E�5��2��h`�F��T�	�����(��,!rZ�S�h��W*�C��'��W��3��7�{�G(��E������V9��:��څ*��0|3��/�X���k-I<��-�2?��{5~�,~���VH7r�~�d�GTx�9���^v�L򾽣} gr{�yygO��)�=鶧��Ɲ_R�Yٜ�g��A=�okeK�Q&rv�S��J���X�%�{��jJ��#Y�۬l�q�\��>_*�ʆYS0s�=�$P�[D`��L��}C,����t��fI�nO�2y���ǉ�ӄ��z4��w�j(.�l�Ji/	+�܉�"���ִ_���/A�7��3����������J��^���q�`d��Z��X003�m��}/u:���g�
�1�9��������y��LAuVH��ũ�t8��x(~�i�� N)�BR��O�9@��C%$��g+(:���+�J޲��$ݫJ�K�k��Ȅh�h�F�wF�����9Q���|[��.ir*X��@�TC�%�i������I��tgc�a����F8��˭ea�X������m_�������9�кK����Dh��R����A��j�0�5Q�sɁ�'������T��������Y������Vߔ�����rksY݉�[{��_�0s���s�����u���AH��fx..�~b��1�mt$��m>/CU�r茞��+�h0�	�����(�%޾gw5�d?A��VW@M8q<}�א}��I$��k:��`�?�8�Eb |/�{bP��!)�'�VQ$p�	q�;],����Hr(E����J�1ymv~	����2v65��n� [a>�=��͘�����gg�H����%�����Ŋj;y��`�U	4��D퀐�� h�ކ"�%��pJ�����e�2�Gں��E
b=�;�E[}z@�n�m���m��T�!U5A�[�IE<[s6��� E䳊�� R|��v iR�M�SQ�ŦG:������O��Ǡ�E�ڎwt�g&򲲰��5���O��^�z=Q��CN���*�)�#av@"SD���l��F�2P��腆j�H�IK+���hL��M�_92$33��<
�	a$S�\�˚�م?��N�O�u�7�����{�bau���	�^�V�Q��y�m��(@�K0�9��kHn�,p����{�p�����t�fg��.O./�tǙ)�5��m<�0��h���RD-���<�"x��g��2�7ڲ���8���KD�d�<e�ڔ�ħ��$�t��!���?eaj�T���������2S]�>˧�\�����H�B=�����>��r�X@��陘Ig*���.ʢ������ڊ�h�ƣ�?�|�a�	 �W�vF�?����m����N�/$����|�qfX
��I=)��]NT^�q����P�Q�}��<���.#���¿�G��zF�����)�C��>fIN/eߜ��1�����t�ڏ�f�J�	�x��_%Hb<�4$zz;*����[k`��AK��\{�>��<j�Y����)� Ҍ�A���p�%�C�SݘF�_lNp�j��PΏg8M�ؤN0Ҁa=�ь�w{9>�# ]�2���s#��b-��D��Q
�ˎP����?�M���Fio��7��NW��~���7�Wˍ��H��Q��#-��R'u9��g�'rۿ��M�B��W-	2,�Q�5;7�vd�����լ���B�6��4���m�G_�&Ԇ���N���r����@n�-�O[���f��7��I�����Ojsb*
Z�5��	�t�LR>�m�W�ry�o/�\B�p�?~�S� ��G�]B�}����j:\�����m����\��Ѻ�:};uL�I�=G�uN�-e,~"�%�� UNn�ݞ~��h��@��
Q�\^o��E�
��^�Goَ0�4�H2�2�p������M��ܽ3W�d��giParhF��q.<L$�2O��(�L��:��T/^&�)��8B��5� ����T��HM��R+yg�x��%������:�:���ǋx����[e�E�����(L�i!Iv���ѽf�lv��j��%'G���UD�v~�29�Wl'��uXL��l������Z�m#.�-몷��?���>]�[k�xX�09AӶ�{�Nk�����4t��T��<A�׵>mo��B/U9&1p�ag�C��Y`�hd'h��~��dc	�aO�.x�~�0e�9���>�z>1����$������vl��#���n}5c�Pw��@�X;sD�MYT�P���nΩl]�i��1��˒��V���ͭ��/@�ϓ�#Yx(�3@r�1qi�R���-��u�#K���BHkI[���J�d�� �L�1���p����&��*H�;��#M5�8�����$K[)�5�[�-�b��<̮�2�x��Q��j�!$�z��1�0N��B��̂e�j��[��C+���c�p�/��l�B��A38�*�n�;\ix�7;{�|�4 ��g�v����mN0͏I�.J&0��Ma�a�:�͐���'���C�T�߅�wَOs��WP,�C�����?
�|����2�[�P&'+�@�b�(U����3 �n6�mƉ�5�n�A�,�tc����P%��G��?9Z�x1(0T���=��Q�3�*';C)V^�og4�~��E����W���I}@��(�U�|.j%������w�	B������j��V�@�nP�m�����9���?�D�X��Hp�+�/_f1����0�?+6֯y� ���{)c���岼�;i8[Q�W�/�Ы-C�д�5:6L����јysE�h^�L�Į���� m�z�ŘS�4m�V�X�YF*"����z�gXV7m�\@;�3��r�8�(���0�0�@Tr�&�����*���Z�E)�Q�[��_,'��[��t"���q��e�B�?|0��A)J��!W�����F�%ڟ߅�*���J�pօ!�C�M��VY�d���ڏ!��OjR���y����>��b�jdLh��;:��.�5�y��|���z}2J7���H=�IGHK�[F�&P�4&y�n�ϟ٭��*#��ޅ �9� �h׹)���]����Ө�ё�jР�Ĕ>);w���_-��;J�PcA��z�	�,u��6��{����?ن#���.�x��hi�<f��at�����P��zxp�r/y-�cН� �yBj��{��[;�,�?��p����{��V'Թ�P^�W��h�:�aO%��2�ia�k�{�7��\G�.1f��T1t*��<r/���g��)�I4a����r�-fU�}�.����9�����$P8�������`�B!�m���O�"� '�䵮��i-y�	 ��qD68Ԏ��bI���_�ě���y�r�,[G �}�]�� �˘���PP�``��U��oE;�D�!E(U�D^a �9C�$�io802[�ࡡ[�[�<oe8�C#9�����1����5v��6�|R�����w�������3K�, �s���Uܰ�Wc�O{ �����Kв Ǜ��(Cߘ���X{?8��Ű+�*B�/�J�6u{��N�rj�{��UM�O�3I�>Sɀ?���=l���Z$KGT��V]��/�����
ɇݔ?��y*�:�p�6G~�/�-�F������D�t�E�����n������� _��Ck�_	���T$Da`�8��+ď���\Y����{у�E}�Dˆ(3S���r��h�M��[���ّ���qv�w��B��|A���&~�����
ύ��֠����kL$�J��Wi�7�BJ�'�v��Tn��S6�PL�03�V珗����s�h�2���o"с�G�,�?P�͛4��y@��l.��W�C<f�Kܝ���J� ϶!�5�L#���t�����Mńv�&���.�-*��S$���s���I��Ȋ�i�_A�6$�}��ϥZI��U�L���t��1l�_o ��g[WE��ͱJ�nl}b����p]�m|9wi��c�	�7����̪^�Sq~���W��@���`=���y )@�Sy�TMG������ܹ�*�\y�b�]4�&���~����y���f�&9ᗐq#Sm�'HI�T�6�%g�����Խ"Z��y���Ԅva>���!�5�RxRgG���Z�W�{��U �i�:����A�{��9Y���Q���$Y�'��T��[�ɩ\)�+3w	�����MtzHY���N���&���6
c�l���bF�\��ѝ����hS�v&��"_���'�fiD~F~�'5$��NQ���G��  XU��a�޴�$�e���G�[�+�Qi_[Fd���W��0�q��y�5��CW����nR<J=m˜+�k\�ǽ[~l�j�p����-8���A�}��DC�ǚ7�Q�1p��QI<W�o]���R�q����9��66rFY�.�?/Bf_��M�(H*f�ؘ�,�@�fz#~e{��0^yf)�xc�._V��#O{�%�?���P����l����ij&�A�����@XI�s�A�C5��p&?3�P�^^jOc`8'��h
>�� ��_�J^F'���a�?m�d`�B�̬�]DEW��!����og�8&��q�ݭ���q<}���M�zK����u�,�l*�2Z�aZu	T���CqWS=��.��΂��<mD�+���[�N�S��hu��e�p���O�(��e��QU-0V5�`���	�]�X�1�w�:>#�ް�U�=Q�������J2�A3G|�`A^0�(H	������&F~�����Df/�m6����w���$�������5�O �]��۞��K1q��I�wVǅ%A>�v�x�=����/V$xp+H��b&Gh�\��K�Y�T�Xv��ʉ�y~��{���H}�z6Rg��F����U���`Wj��j�b��]w<�$�9�ⱈ]���^��DXǲ�y�1�E��-�y<n\)Q�:o��\������1K	uP��)6��U`��>޻����ƛ���:�sƪd/xi��B��R�p�1�Y[�9�{(��I��+a�Lc�����R1 Be��-7,�&���?k�9;�����x_�9��e�� T��=���QeN��E�?��)�����k(�k��n�){�(�W���@Jp�W0�=+�rsp�ϋ@�W�a7q��h���n716�y�zL���P=�UJ�k�N��2�n��3=���"��Gs�oI��f''��ꪽ2�P����YB/Bë��v�K���*���m���[,��������k�e����c�y-Wl�z=��B��I�� ��"���p�_#E���M�r�O�a����s{�\U_�bQ�׀�xXFY�N�J�w��Bx\�ؑ��`V�>��+�hG��I�|v��O��]<�X�O
����_�b�_8%C�J8�ym�G������\]��X���/�_�*�i��ݽH+���m�a��{�o�s���e�wjq,ad�~��!��OD*k��
��C�9�����'N��d.��	��U��,C��@�qfT[44��ww'P�~bC���l�$�����ւȭ�En<��;{��dC�*5ٰj�wMՙ�Gq�<���u�� �Q��_E{M�f�[FmC̠�	fe�o��D&���?4������y�-����Aж�J�>F�z�7*��N7|�6	�/��ܜ��!G����D{��4u�KX��N�	��z����p3��2����qU?��џ�}|�]�+�J�J8yD-	����K{Ǟձ�b�Uuk�M���wܗW&����ؠ��@���М=2|[깨T}KS�GD�2醅�!vy�}�Ǒr�T{�)�Q�4�}b/����j]���)���$�I�i�E�Z}�]��r�S�^�2:b���W�&�w.����'�7��;�~�]�?;���+Q�x��� ��L�X�_�.Y�؆���S�h��[rd�> .��g�Ĺ�(��IÁ+��p��#�#�k�H����q�
��F� ,�S ��}W�����T�y�Auh��o���h|
c2�A�E�j)����v��F���L�8���2~h{�I׬�=��e�JЅ�DEc'��_:?7�P 1����������Z|�K�������
M9Qpw�RK_���X�gg'1b����9�����PE������0�����K�0�<�'� �Kz�!�/�\%��CAE�p��țq���
���j�82����(��x�e�wB�*sO��/ӊ��"�}����r�xTV�{c8#-�_�&��1�ï��¨�I��YF��]��y'E����
-; #������������>4��4��=G���|o�f�b9:c��wҀ��`���v�E�cf��M��~  I.(� ��cӴ���Q�eF^KuC3l�K���M�h�PQr�]j}�@�H���:7n�Xr.p�j���(F�<��;�,�o���-�<^��HK�ř8#�I���]'��H��8�Ȣ1?6рl��i�b���SG{S�?�X�e1s�Q����!�vZ{$�ķ{���.0C�Ɣ̽jH�c&��sL��@����|�k�e�7�.:�a�;��_ ��^P"T"��P
~�f&T�;]	���WI1���RW8���f�P�\�L����~cZΑ]�V�:(y����w2��F{��U����� ��C?�eQq�D۞��(�%��Ud���mWdZ𥦝S�)��Δ{�!b���߲��L�yVrr_�o���$x,��m %�mʇŞ����X> 	w�`:u1�S$����U��$x��қ�7�,k��I����Ԣ�=�[� [nd;�R�O^�/���77.ģ�p�#�L�b� ��EJ�i�[��C�	:�/�ՠ�Z�֥�c����at!�Z��W�;��$	Fb��Q���B�2���� 0���ګ����PBf=��l5 5��]��y06�]d{Oc$Z�Y�X�v���@eJ�P�s>�@��^]�6Г& *�#�&�F�U�VK�}P��ns�p6)��Y+��\`� ����*���v��E�����t�eJ�O)�p�(��[Y�AƩ��`��m ��~О�#����:3|{I-T,�Q�m[�A�Ǐ�FYX�Ҳ��Uz1�����2���-\2�j��4J��~��4ߵ�I��cSI���N�w�ch37�*7O ׽>���f�����*4���"s3A�>�7v�K���K�27���̄��PjZm���M�x��g�)?"�vy�&���T��*^ �`5t���*��A��r���k^�a�8KԗzE��2��t�K���R���g?���"J�U��ׂ^G�x]>7jA���83YI|]H��JR���p`5�����Q�A.�.9�6`!Y�M5,rG�b����W�3w�L��
M:q��,=�6�i�E�{σ�}�]���1;�w���v�mSЮ��7rkY��"ާ�����u�e���ڰ�@j�5��-�]��X��׋�f���S�	pꓐ3M���<�w��cP��,����l���c���6E���[�e/���,&m�g��@ҢF�N�	,�\�qCǕ@��<��cZ6�UN�
bm,�g�KRk��D����*�DYw��vc�o���K��-���F*��m��^z&�+s�n��`*�t,���[m8�N��<�y�G��Ӊ�>�o�xg��6�M�.MB;�/P�+|��R<��l�E>�%���T�*% i�S|T�N�����VS�}Bէ���A�}淨��!���ͬfC�j6��#�N1���4���"��h��΋%G'�g�leǘ����s��7�:�m���;=E�}�6ig��A�����{Cl��+Ιh��<=n�y�g�I]��*�~縐^�w�P���������Y2葱F�j-����p�C/�Q��s�5���d�um�d��^������6`.��Au[�!&2���
S������S*�y�v�#}��w�[��&�-��%LU��Wy���*Vx���#<$�7ݮ�kU{kY'"R��Q���WlA��Y�ό<�M���^�;�յ�A�ëK`�ϳ�HFڬq�,'�8t9f�����Ѭ�[�*Z�r�H��YF�瞃+�x	�X�D�S��sR�?�'ڈ���������]d�;d��}�I�,�O�f�F�2|���8b��������b_��ᬺI��w�>����L��-�iQ�{Dy��� �q~$��W�A b>�r����iXY���g�i.�^o���x9L���
~�n�4�+�g@����V�n*�6Af�����8�4�f�����U�v5�O��P����O5�*f�U�%׏I�Ego�L{0��ޗ�~�c�{�,zt+j��f���b�u]h>����?w�#$�Ϣ�U,��\���[�QL�˷.���OdV�ob֥��JRox{o�ԏ��@"������f_��ɷ"ԏ�Q��I	�I�b-�6��}�.ۣ���'x�A��FX�V�kY�tU7��7h�Q>P�}�����/�N�b1�� s�]KX�f�)�Dm�S�Tۅ�(p�p��t,U�'47�Z�3�g��V�y�b:���ޯ�Z
8� x3yw�����-���{]����<=�A��/�cP;���o��Y���OS�����������{�}ڳ�ɴ���=���T.��@�r֑����:�2n̙D	�d� 	�x���c����s{L��Y`�Tαg����'5��Ȩn+�����8�*e��r��"�ۏ���sw���V��wJ�_Z�iC���Ŝ��B�����W�$f�#��8�tU:��y�cT3\���dsS?����ȝqS��VNBi»?�|��ȳ��=*^�I��x���K,��w�n��T1|ٍ�vQ��I�]N���0�X�i��X~U����!}�_hK�>��5g6e�X�{~;Q������3��� B�T������+v�Kw4:2%��3X)cR�^���@�3��&��Dʛ�.�N���������;������<�eU�qZNդ�6�Y�h��d�D�y=<e�&T04 B�"��K+�N#�\�DӺQ����
�=L�dфh�q� �Ѥ[�nd�Q���{�vx�k�".�c9��n�
��Qm��`WR�ķ!��%?<]!���J�����'����}��J�zW�C��q{j&�R��A�ĳ��F��L_�g��du��4���){��\� �@�A���m�H H����&E�۞��z��t�����O�}i�a���?`cY�uiU�-3Ub�Bѡ��NK#<�UF�R��������"�"&~c1�]�v5)3��}n��X�]���N�8GlA��%�7�aj��������:�	���5�%��0�Zaڪȥ�W�"�[��U1������Œoe���Oʖ�Y+)�d� ���d�p�b���%2���G���^���>d�������I2�U�W�p�Q�r1X�x���䓗J<��/!>t�c+6����k���z	,�(O��C��O�1�!���u�YO�[��Pg��|�1A�˳١��;m_�����K~2���X����AR�t3<�4�<�m��1?[02�YLa�w��F����JZ)��������T��Xu�'�\���$@9��ւ��&��gǙ�)��g�ʶ36�^��1�"��p<�X�s��G����j�\����츁t�
�5T}�����@�D�}8���mo�ո��Np��Rm�g%�qqBlE��P8�jI��r��gӳL�c�����v́<�7��t�8�X�N�� +�ʌ���ْ$��7Q ���^�,�&Twm�u�6ex�g���rg�q7s�7�5�%UZ� Ͻj��ןf�Մ�+ ƻm�Ϭ��y���5�0�Q�t��Q��s�f�v&D0�.�w�@1����2N!S5H�}��L�dx����
�p��DPV�qh�
e��:�S:�K �R��+yq:�_eߩ�%�K_o���,Ɵ
Qv؂d�'��$׉847,�F��[�_�t�m����^����o������Шj�2��s%ȯ4��h�2�E��7o�B�o����y����rDG�2���l�;)�Q��-NU����g��"P�.ĩ���e,E��+�$X@�+8���ƃ�X�����d���O#w�~�O3sg���������	J�2�7�\�6�O�F13���ϩS5#G'��.]�B ���K��:�{Y�'���^$"�wڟ�XS�f�Md8�`���D�p.�u�B�+��^cl�O���4��R��ORj
Z�OO�����"`�$'���i��Ik\�*f�����'��!$ȅ�I*���Y�ѭ9m�7�I���8
.5���@�1��O�`�k1�S+{�rH�$i���km`"$t��A@�_�Vb���>���NJ��?�<6X�����_���ޓ�n��M5���Q��H/��{��� ��cTĵ�t!"��ʐ��(h�|�of#��T	Jp�߼�6�a�L�b��gq�B����5��Q\��s��ME��Z��\��$�nx����Lx,�
Pb4�i�t����_�$��J({N��R���ef����O77�R���奇�S�h��!�x�u&uٞЋ�%f�Αt�e+��rV�1>p�l��*p�t� ;���'Y^���ާ��c�-wH8H�)���E��h�3�\������?76]��ch���k9˄�m뽳��4��7��\'�y�;5�.fc�f�m�|��R2���J�A���WL�"_i�S�^}z��w����%���\-K�{��G��Qf ��iN�6�[�Q�'�z	�E�܆��4[����ƜMT�Qzr�&D�=�^zܓ\B�@i>n��HH�z�� N�bzh���/p��"+�XK�O[4�a��\]���Ce�(iF~G�#�[�D��4��&�D����H&��
�����8�'p Y٨jw�E�駄J/���C�?�bc�/e:�|���/n½�"�⢹~��Kcp�a� ���~��B��jV�L~��rم�ǬO�7> �x%�Ԙ�r����+4�n�����p=ȕWX�a0���ق�*���ճ��O���#� ��O�8�Dn��6 ��hJWx�8T����j6�]�'���Y�a�r���F������${"r�&�P�[�P#]o�{�Jʒ4g^&9,|��2}��{je[�"�f>p6����v��>O�ٳ޵
f��G��~"�������[3�]�VϺg-�~L������`e/3�`���k��vVI�#�)yK���W������#�}d�S�fo�`�!�3�P�/t1FҼ{ۯ_;X�FIz�bg @@pT��?`}7�u��yխ0����x	n-Lơ+�,������F$�ȸ0�F=	�(�K�i���ĉ��nڜU,ZK{#CR�dcP5���єV�eC��n���e��<����6����V��բv@{�H^.���(�,��_��R+d|D8�,Q�2����Qѕi:h�9݈f�Pd!<a'q���τW��Շ�ǅm�T,�@�]k�:���H"��>?�V�\B�(�2�.i��~�Z�(���[Ǒ���G������;k�:����+���v�^?��EZ�N�w�����<��B�/��X3722�t�����76-jCd��*h�{�Vv��jJ��4W�g_��&�Ӂ�¨���a�g4IZ|� Ϲj���q�p}�R	��T�����!"w�89<�U|�1�=�4�r�=a7�(.��]ԩ4��
D�,�#�5n,�����k�V:�c4�y&��4~�Fk�]#$k�>�J��'����B"��֙��23�M����<��}�1��36]I5k�8Z��V�X
�L9�D/JK��y�Ii� ��^�ߨT���K^�U��&Rѻ�Z�E�oj�:��p�F\r�ZB�������A�O���̺=.��7�$N�Hs�"�G�?jK<�9�~%�ը��X�����D�X:v5�?`Z�H�q�b�z�R�!���
�~ȕ��`u��z�?2
*��
�:��gz	^/����g�r7f�e�o�)ܫ���ͣ�Q]�u��mS\W�B}�5w`T@�5-�����H�1{�P����ވ��"ԅ�^�lKg�M뤐���:��yBɺ�Zi���(���^�i!�@h�L�z9��w�I�����,��;���Ww�.ǵڜ�"�b�>/@7����uγ�T�x��p�5?r�Y�G�'cn$_?�d�%/�6Ú<�0�^�d�����q�D��.��s�IU!��E��xE��'��ɛ���U)��紀�ϖ�צ��ҏe��u�	}�<�����Q��
"�J��]=������!���,���N_x�,�L��Q�JI<�5�v��Q望"���5����F�O�>@@��3M[f~7}�O ��ٿ����.V��`qqRʳWO:���*SlI��EJF�B����-㔅�K	���5ߋ�̧?7�\�WT�}����	��:"ޮL���ZB����-@).p�﷦��r;����=���t؟D"�}��J�W�.m��օ��Ps����,���6�yDV����I���$�Gh�E���7ʈ+�;6��j�7N=M�2�4��Ws�V�!�|��M&(]�9��S��f�|�}�	�H�p��dֱ���w���>�.�0�4OlF�R�bƕI@G2&��K8�C��-;F�S8���a䖭!�$��27��6Y��&R/�=�~߮4���
�Ctx+�,��};����LI܅��i3��e���������׫� M)ҳ��e�����	m�o>����W�U�V����.�+(�_��c��Dr�A���R�m��"l���2�T��_N�1��3�R~í��-=�N4�
V��Dv�Bf]�?x���/�Ed���kb�W�"ׄ"�@E�2���\�
_71����K����+-,�K+m*/�w����,B֮���X�}1�n:��fq��e���Ƚ:<�.;���!��\&I�+vj��5:�p��i�l��=��H2��WIӃ���.*�Rʪ�ްD:t%��M�V��c�-�۟��!�޺2A��o$P��
1��J\(M天0Bׁҥ�=8Q)����� ���w/zz^c�&_��=V�Sp��e���*�&��ѩ���F���\/rf���V�
vIMoMT?�&� 6>z$"�����\W��8QCb��y��y��漪v�\Þ@a"{n�_�~{ԃFj\l��Y"H&�-%,Y��L��N��e��T��B��;��u����B���]]޳�c�[�۹ec+�8��6oӴ
0W6T427�(�������T�#���G��kc+�u��y�,OＨ=N~`���LP�y�ٕ%������m�&Y!�X��!w���(�i71�A�c.ۄ���i�|"��$�������*>��� AQ�E�B����y��B�J�:{*T� "��t�"Vh?Ey8c����s�]5��գl]�:�k˞=�?�ƈ�����G�:���[���^�θϤ�u����x�t8֩ʞ����H�M�Yø��⨗�ހÿ:CȐ��:���Jk{����ž\�3��鮁�����hh^o[F*� �FE"چ&��?�@$�Bp�ꌞ�~����?\!��|P���XC�8���>.[W̖ �e�E�ΊC߶���Y?��=�.��g�\�p]��K����n�v�ѣT��1�\�������]�c�Z��{�a$!��c�o�(����#'�ʣO���1��f�W��߸��J�u���E�FԻ@��[���K�����B�H^nҩ%����Z
�k��[�N1�q��i�\Y��(]~�K��ހ�G����x0�ہ�A��-+��r��KK*�)��aV���$	N��W�\c��l�ҽ-���򒽚@gm\I3X�Ʌ����'%�UOl{�y����>C�?�	tq�2�*��6x�dl.Lդ���J�$�~T}5 Ӎ#���ʄ�ƀPG.&�̦ODZ�N���J��Yp/�MuP�LT�_<��C�\��u�r��T �yK�s1��g�t��&i�������5S���E�7�9��澛X��sB�ɚ0�3����3&a
���	�)6����Ь�;��kC�zaК�S=u|��	y0�1�F4b��q���}�CC!�Y����K<"r�~b�g��t��/�&�8 '2@�(<=����4jbH�US���i֖���{�<ظk�ś�S�5�X�I��R{"����#�\��O}��p���� 7�^��.�U��1.��r��0�m�$2�U�1�Kg��ԏ;)s�$~H�	�n���?�ME���-_�� 8J�H���|��M]E��e�:�(� _�����PU��JIK��dg�/e�5~��fg	�����fYӟ/*&R ���������U�GD�Onuxo/l���Np;�9��GPd�y���x��]~��U�Y���
�xKF����5,ނ+�ɋ���ȕ;�/�׮B�ί���G�֫�$�L堅��}���Z��A�q
�`|0�\�f@�9����w�������Jp���!�92�>�32�(��PI�Y��h�C�2r��{��P1jk?·0x�N��1�B��`K��t�
���xK�`�6I�����_���v�"���J�6���P��`Ø�8_F\0�7ѡE������Z��qُ}���w�'�%�]����O��rB�&%R�� m��d�sn���P���\�u�0P;�]�m�E���&m���T�X0(L��,{a6\^aU��8���7�}d�>�D��R�5�����C�,٥]ã��X4�w]3fa���]��m$[�RNT��vq�ŋ������ I�XH���Xf`yCϙB�ͻ�nh$Sv�����-c;AD.��LlVF��O�ɴ^�^��nA�;`aW�k�3��?�uՈ7��Wtv9�B�,�d��EUi��)���|���e��'�N(m��N�RK������J~g5/�w櫬=b�S0�q�4������ɯ�l�{��, [cC�WF�Y��G[�G��x(�1]��E��f#S�8�J4�>���63؇ȷ�@?����T��`� 4�Iz��K58��CǦ�$�b(�y I���})����h�r`n�� Oz?�z�Df�P�ke[I�۠
�1ʻ��R���ټKJN�;�Ql��~*T�ݑ]�݅Ԣ�O�7#J�B�u�վ�p�_�3�M�R$q"w(���{��oZ�f{o��,<�����I.�L��
�?λ�^�{ꐱ���Ӿ~�����T/p�^vr@u'D ��.��8%��V|�`W*_��E+��c&M!r(vy����>�9b¡���,�lsv���\7�"���������n���RMv���lj��[+�BHͥՕ�=�M��<�	ix���nH�������T���E��1͊j��&��&-���5Y8D:z�čY��X�1���f�-���<2������E���Á��h�mR��t%�����f
��G~�U3R��C�kbp���?�d/�ZTS��s�;���@0�lz�T�w���D���{�Ej1OG��qV�������+����?ɭr�(yF�&$P����#�Y�i:�����	�&������s|Pwx�i]({�J�>��XFm�3)"]H�\��k�����QՍ3�.-�V+a����8P�*19��yn�m��iE>����qb�*�s�i,eU&�&�(zmWj��
���Cq��������{�ͳ�7Nt��c�*z>�1�bXB�~]	�i����({�82TU�sL!C�]�#l�W��s�AE��qv�=@���t�z����#ַｵ߱����x�L���P�[����٣_��_iSAH��lg��j繟V�;�S��/����Mh�����V��F3d�
�W�>Pp:U���I���[�Q܅׃]h����T7�,�����y�ߒ}T�(�Z�s��\�:� ͨ5v�P�7W��XߧD�ԇ�������-�U���H$��͵�
ɵ��N#��p���-�U����i�t,���!�=���
Ӯ�#f$���J�΄��]�-�����L���j�����#��t?�;A��N��
�7�ꨫ�9��@l43[����'2���q�b���V'�fTҰ�l�zyQAxa�	:��К�ВI�1��8-ع��K�i��?��k숥I0�X ��t�"8�̶�T߫�2R 0;j9�!v����Νy�����+2�jr�J��ڦ�
Iz�*�V(}����KF<�Kqk�;���KH����#"��������ᛄȎ2?��.㛻* nH'7���CR=���y������N�'%>�?���
�d�s
bӘ-�^d+f0Y�<o/�Ut�f�	 �?{A$C˧w�g��ʚ?�.<�Jʀܰ���3"��46p��քy���w�����8�b�.�TG�P	��iϽ��N-�)&c�Wf#�)��	��F���f��ǃ��̺*�J��k����mN�E�V�:w���p���&�dR�������V|fA�cg "c�uJ��{������T��̃&~����|�0W�&�<��b��p6��V�37���v%�Z�윇���C���ݏ��9�����)�#W��a݊�����w&�S����q�������� �.�$V�J�f����u��l�!�E٣F�p`��#��^��r���;d(���#Af��<s�Z�[�M���x��,E���bq�F3��Z����\Y���8 �����f�A������z��К��zDjGӲ\P�t/�@�A]?�*��v0���&��0Mc�#�[�����.aN݇v�2����+��f��Ď��+���N��h�Hj�����l٧G����>!�Y��e�}��ahL���N8�6��T#�z��$u�N�ᔳ<����m��z�ͯD���nH������o�����9)�ۅ�fܭ��o�:RvN��4ټ�E<��j�]������]B�x���a�9�Hex�$�"ښV�"AW�h+!&N�����EO����c
��0����Ħ�P-Ҥ���z����°��\�rl��7AE��22��p'-D��ھ,�?���/��k=���d�ic�Z ��s+k���bwǨ�-��xz��������O|M��?x�O+8�I�	W/G5dv� �L�@�`� I�">;+��4)=�me�g�
�<�9%���a�l�>AMa����B�C�8fxt��/�Pw�����t;dg��ƀ���B����4 ־V��ȾO�Ŷb��s���p�A˰�,���	aM�����W�F���Y��.T���!_0�'��L�� ը�����CX���j�d�ύ[׆�N�9.�w�x�CNA�|�8�S�I�����K�D�O6�Ar{��srJ��H�ғ�H�u�9J�5,�Ǽ�K�~�#��13j����f7s�j씆Mޡ�3C˺�Q΅��0!ʦ����(���X{�KWo��襶���;�kڇwz@�� VUC�3c'�����d2oߜk��J������S$�,�VJ�ðS	��|�4,Z�tNFù�v�.0�O^�Zx�]xv���׳?(M
��E#NI��q��d��e�n�}�n0�؃z�-=���I��
�H�kl���eT�և��~����P\p�PJT�����Ӣ��V�	jz1n�޷}��}g	��5��?����\���'Mˢ�M�46I�i�<�!�6^b|� Mn��):����3��M�t4.���rs!)�V�x�N������*�OP��+/�����`��<�*&X_�y�����~�<����O����|O�M(m&��`���r�B�FDb�K��T��=��n���}���˺�k�v~�1�w�>E8�����)���4��𜄰�?�k�'/��a�>���&�SY���@�E�g��0����V�>�,�λ��8*�ݬ�~}��|�G�S�p��N�7��eP�4o�᎔e1*�1$C��xW@ȗ珬@�r�o &L^�Y����}��Z"����!��X�#���R���N�ă����jvz��9��7}�i[j�S���GI�[���__q�y~��q�/�q(ã�ϭ����,{7��yH�y���Pٶ�;�`�)t�5�8RH�WP �Зu��\q��¾�RQ'R|H*dJWo������1Λ|A�e滕��M�5��J�N�G� ���9���4�8v���1��r�zW�A2�(4��U̷W��$F����4����ۀd�<�f�O+��BZ!���֖��bӚ"�n\�骡��
 ^���x�����A�	�ѥ̝3A� 'lؗ۱S3�p���q��zğ��NB��$y�p=>�xp�f�cT�<���o�,bʯ<�%�B{�J�Y�٣���
�Q��cS�7Lހ(2�8�S�;�;�R����8�����P�����2C�mvI��awv��?��h�l����S�a�F�9�s$Vln�X��#������k*JI|~�;��mP=|�=��y	�.82��j�� 5{0 �R8��C����	�:8<,a��~t�*`�5���Z����c�Md�L���]u�c��/��
�~� �z�Y��"5^��T<CM��$-?x@�ع�jL��万�W�.����t�Ú�� ^N�����wu����n�����5������G�$�=��4�'���s,��
\���]*Yح{5$cF�׽y�֎Rv���S��E��H�-���A1��O\��O|z��Hj�b���/?�(�B�Fw��4���c����Tzk!��ׇ�P𲊃i���c�-��F~&p�AT��?�����,K�>�v0�b�uO�ۅ	5�w�5��jKso�[p�4Tu���ˮ2��+�!�^��i�.bנ�)�;�[pu��\��4�,�*����?�]u9U���L�+
�p����k���2��P��qA�� w��m��@8���ide~j�h�z �x賺qKCM?�F Ja��XA���EK���M�W6÷�]�6�m-����W��E4��˥Nv]�&����D����<��b�����T�B���}�s�k����h�ۛ��!�X��M���+��u�WT9�^�N���TOk�D2���k .�cz��k�}�p�2Ϳ]*�֢%�`���,�"2�O���,��n$��2u�񹉠�~����
O0U%@�0w�Hխ~��3xp˦R�G����b;-�]�<o'w��Y/C$7jv?�ڢYU��:�-{��&&!l�}���\����J�s��]{x7��G��4^��Rc���=+]���l��L�<t�;�'�������G�v��?Q>c�z�CC��Y~R��z3z.Qf��Y|�d_����p$p�u84S|E���_l�7��m�z{i,I�:�9�ȩ��A���
%��?���=,�q/���07b�t(d��x�'��]xΈK�ֆ��|����*,ne�GY��סa��m!���n�ed�oV���~//�>����UV�(ɺ3B"����6�[ �=c
NY�K���t�a�HUBh��3UM��c�Y�h��W/O>��%4]Kj�b\�7��$}��!����[���C��|C�1!�~'��ƴhO���ø&�B�tZ��K���?8d}�p�b%�̂������|*��ަ
d#C`8?ͅ	�ɡ�\���{c5��x*Y�ZQX�!��<S����{S��OC��s[l~ؔv�?Ɇ�脰�^�����J���w�I�G� ʉp�FH�q	"].NwU��ũ���#��HC+t��)唞��2�e��xWp�)��fA�ZV�o�e9B��,�����;��x����'��V��!�2��l��|5L"Io�hjy�,G.��F�s/cA�S�ɓD����v���tto:��D_y�DL��𗥋nv�Ͼ��زH{��c�)>"	������4�?[L���b�1�Xw�j�{���P��Y�50,V���(��f�e�,�s=��C�>J�#����o��LZ���K?8��vv�`�8)�=��.��k�Z�:�:hN8�o�ը� r*h�7��Sv�Jqb�e��&�X�+w

,E�v�����teiz>�>̠6�$�0^ߢ��r8�ֱ��b�k��62�ZP/�v��|�Aǵ9E�ܢ�D��o�*�����T�^RSk��t@p�_Т*�ۙ��{5!n^�C?Y$��&Repg3�� (�s卞cX�B�nIL{�~}�Z \�b Ztx<c�`��źE�X����~+8�V}�������#$!��h��@�}�jF跻��÷��c��k����EE�p;����h������NYp�Bm�� O' ��� �n/�����<�bZE�ұɵ��>��Fy���[��ҏ�?���zC	�
PB�92����WG�+��� ����u�q�]>
��O쭐��O�O�k���W�+��uJ* �F�!�	.rQ6��y��QY[�r\�s�,>�}�ޔ���ѣT�	 l��xw0���ݨ#`X�bj� �-���f�8<̅#�:�&���4�b�N�8r�`�9��8�g(���u�_S�x\���A̽�l�s�b��3�*۬e�tr9� �mL_-�]�/0�am߈�>`s������-Wd�U>F��O�E��
�@Y�-�bO��dL�`�嬉�}U	AP>�VǶ���6R��x��D��p ����e��_�9�`3���kS�\��zG�r4�����-5o������DyB���u�ۥ����[�G�7g��DOo���j_1��}/�!�Y��[�!\{�ğ��E������ە���2�L̛�*��_��m���0���h�*�9ԉl�+��¿D?��کr��KY��>g�h}�Ʉ{64O��Ja�̟x�H�o�O�p]��t$��de���P�:з��n�$�7h��7V��&(+T%$����(�׶�ѷ�����T��s6t�0ε�3n�-��d3�O�* ���j$�՟U�a�Xh��^(*���O�0�|����[V��0�%��nnf��x�p��Gė�h�	f2���R�!o�oGF@}�L�6�$vKĵ/M���5���dj�Ɩb'B�r��[P6܉q����������dp:�Y�kw�9�r1aMf~�Q�O;�4����~�U-ٷFծM0��T�����Q�{��Ӡ�1<�`��h�h��^)n�������$��<�1o0~_�^g�$�J�6�Ә�$���bCߣ��]��#|��^قtU��^j�d��1�۹����z-�Si�fL��a� Yy�#lO�n���K_��u�p�G��� ���U�9����r܉�6	�R��ٱ�(N�?�-`- �Q��b�w�-��<N:�:�����Vc[N��H���T��j��m��l�u��[&Hg���
~�wq4k�14���	^Wp�������q�"��i�=a��zG3?��^���g���pd�}��f��:Y堗c��T�-�=�
�w�GP��4��	��0�iL�#�����,�&�\���=e�F@cS�@�}�֞ ��u�$�{K�ņ�%Ƴ��ݸv�پ~%FڕUwxY1�6��U�[����-�z݂?�9�c.���vF[dsDQ}O�D�P���=�s�hP���͢�۽��K�K�phR�E�XKq&����!����k���ϕBvr1'=��%�G��#	��7��,39 U�蜏͗��	��_ ��Ձ:�*^�%��F�+eNV��I����*%��V�8t��X��p�u��S���B�~����K:U�w�;��ed�7���h}�+�l����NO![��io���V
��;|!ڐq�q��kk�-:jw��,��i ��A�qmԥV@��˗�}�nx	�A�d���|�|å����sw]�b����`��R�J���KУ�i䢋����Ƚx,�~3��b����5���M��[I��[5����J�6��d%^y��	����P�i�)�|R�b;K0͐s�1P�����`xv����h{�4�.&lu�z�}��`N�fE9�T���T!f����z
M��Oߕ����r[����j�J�*"F�m*����1%N���T = kT�����Z��H�:����*X^L���-{n�g��^����b�'?�4j�m��aE��]��V�,��3K��2݊�d�&<��ҷl¢`>�R��3?�2�Q*�� 0ðP�c2{�|�� 2
��K��n�i(]�d�F�j�<!���Md1�F�+���/��H��!��:�x`�1��rq�e28�"�
�
0�O����������U��z����ß�N|X��������:�l�U�-���]L��`�5��z��>`�"��9��Áv��W5���C���������e�ou�����&�A�$E$/��zn��R!��K��z��v���^`�ĺ�]�p����gew�T7����@���v݂w��@P�y��e耦}�5ށ��4�(/�,�v�җ��K��`E;#FU��t�n�"�d�0�� �ȍ��`D,x8���ԯ��:5����!�c!P1�㷺���V����F��%��(��8:����P��x� z����v),�y��f�B��<�vrC�K��^�0�����a���Q��(��<z5���VhM'6z4gf\D�9H�B3�H����37�>��:�K��~dgo п�f[��[5��Ms�0�FǫWޣ.$%�FC�d]��u<����-P�qLRj�z1�<`�.���$2Va���)d
@J�)C3��'8��M*��7���oJ7Lt?j{���sS�F�X�q�����}V�J��n\��R�7y�X�Fu`�V������3�N*�7�h��0��c����8���;2���2d������Q_!��gn�o��u�i���K��nN���^�vt+4�6�A���e�q��0)�BP��𤀨Q{�����7�-�(�6"�	w��P1whX�hV}�o��O���gy��`��#�"&<eboQ�]r��"ƕ�WV��d]�8[٠��)_�X�:�z����L<~�5	��@x�=&�T���ܘ�a�6c�v>P�/z(����N�H�*t$��6�>xCw�iҐޅXd�E��s8����������rR��kR��Ccew��	��k���`^zE=ʋ9��?��#�s�o&-�����D�м���p����]}z���+*'����Vx�_x*��uIU��F��+n�}_A���	~*�����~�I�aCD��l[� |8f�f7��Ď�nY���&g����i {�q#�^�ʷ.���.�v���rM%ُ�D�<AB7�8 2߈p��n?��h0=�=?_E���+5�v۶���U���:m��u2H~m�x�+,��x
�
��E�]6����i��1d�u~$5�?}��;�9���;Z��࠹1!�u�#��搖k�Y�]W�w1��)�P_U�8�i!�%yu%K����Ү� �
�o@)��p�ŦMJ&�YtG6k7u�Uz�6L`�X�	�e��0�ȭ��r�}��Ðwg،Z���Z�;�g�6Y�z�D��\d���+ܨ�:�S#�s�V
���Y�v�@'g�u��. �G�����V2��z�G0���U�?Ok*�Ό��]xzקx���@>q�>n&���l�U#��ʾ���b3��h�X�\�峗��J�/v��I��
G���l��-�2�
fwL�U]s��H�"�(VP����C*�|��2�=,���A�X��B�g����5}O(�p`�5r)A'�?�.	���9�c`��;IӴ�Ӛ>��(��>��üsJU5�EI|�NA��ld�s�}���7!)��.�V/��Aqŋ�"�γi�$07����(u�v�>�S2:l�k�w{2�F<y�X�Uj����ߟ��-r��.��`������Tʀi��
\#N!�d{j\W���8�������zې/��	G��lT~R��P�6�f�}&^�Go�1�<\�r��_1l�V�	°/e��IA�^�U*�h\=FJ/19��y�r�گ&�S:�j��<B;/�l�u|o8Y�m������<���Mx4]��։M�'Y=��*Ϫ��Zs	1�n)�����K��A�����py� �T�!3J����1e�'E��Y.������\Ni�_�i����a�W|��E0����X$��Tn*��;ʧ!3,aC#.����1/�W��;�����M���-@i����F��~��o�B�yE�K�\�}_�'���F��вh��R"�:.��}�U�x0�yA=s��*��e�bKHK����e�j�BgF>x��x-��*܎�/$-"��T��߉~��O����6M�0L�-�����.Pĺ"�Oz@�m�74��d8��g�Po�=�]��^+��3O��RB�szH����d��������!���.�:h�Oz4�Z�R�xf���Svҿ;+"*���%�cx��7�`�C��l9B܇X���a�d|Jg�D�+M���� �@7|�g�\�9�;����+��f0���j��	�}��D�+&��� �o`.�U�߻t��s�Zo{�9H"G�\�Zoվ��G�K�����BY�D��çC�oa�'�.�*^O����%�:<��1����{z~K����5��
�RU�,���:��V#`Ik��8��� �����%���?�2G /,��
�0���u4�Zpc�H��>�C��kXS$�H��.�7���\�xT�>
��]�"A���⫋�Q�|����'���.SK�Z��Cly.���&3��x�P���Z%q&!o�v3�?�ڂN~<̉d��Ն���� {���b)BTж��:� ��H�h�[��Xb���Up5@>��hQ������Ү�˙'�˚ȯ��#�j��8G�4��
���c��5	�{;񣒅�N2��Ik�^}�%܂�ۊ���nr��/6��s�~Hm��\�f������;�=+��F��/�)9Y˄�� A)��Ci�9\5�/�\��o��2=O`���s� 0����֙�R�V|�r��hD��p�=�t��;�����Bg�ڀ�o�j�QZ4��w�r��F��]�Q��R����y��B��6��t�&��\�s72=A��O����ˇWP��@B���hYIF[&���\@ų5�ߛy{�E,�Ze���)�0<8O�l�6�;>�Xc�F��}��g'eٺ(�@��S�G/5���r%g��L��Y��rƂ�$���w�-�M&P>���x�2�c&�5����Q����U�y��X������"�1ޙ�)�z��`�,s@F�l���qٰ���|dm��	��D­�<O�8��Ny�W��X>녂;}�O3(����EK�=:�0�Je���¨ A��
M�j��;=�]���\|�)6T�V�V��F�4��dY`��4���Pۉy���ԸC�>`
��������'� 9���лv���㞳�m��sŤH�S�X٨�{b���.����W���~~� ���6�q(��<��?�U�ߴ�E3�P���@�E]�飃 ��D a絵�`����Ş_��]��D�o�]��υB�6� �9�E�NI��qd-K?F7� sg<"fmq�1A��%5��l��.$��fL�S]}�`��|�K>��su!�C1Y�	�2F�W��\�(��upp:�^}��w�˿�W\Ez�x��/��YYbζ^{ƓSε��e����������p	�w�c���)Ty}(#�Z�}��tyA�����K�'�
�uٝ���"��0LE:�dQ�n���Nca��|�U�Չ�7�q���{K?��T�����^��ʲL�� ��������c��-qk�\��D�F���5uK�
���5B�r�W@��~Ֆ�'�?ܷ���2��"< ���Vོr�����@= y u�x��p\.�؏4�艎�;�?E�پteU��v����i��r�{���/2�Y{�r���t9�Q8��KB���<��k��g{K}1yAf�g\h������ܰ�3lm��m���FR>�����c� �UB]��u�.������9IVX�iU\_�8�����|��si7<�o����=鯄ݣ��Ȼ�l�)�d����r�=7�R��^Ǵ{i�W�}'hӑ53Ui��Co��y1��pr�Y�`��x�� �R��a���g62�V�����Oҙ��x�J�䰍.�S�n�@�G���-Xn��:���N�(��E�E:p62:� ���4�G�|���ܸq��=}uv�������$Lf��"���9��ٛ������?w�B���@���q=(僄wǐ�:���o��[��$D|S:�+?�Sc&H��.6���M��5��Չ/#��*V�J'������1��7�����"t���9��s(f\��I���y��T��qqzŽ=��0.���Bn����8$�~����e��C�vi:��v"s\�(��v��I+�Zo����c%T:t�Yfy$.�$�ˌ��Ǥ�2� ���-e�.���%+�3��VV��o�8{����̓��Z ̥ ���@�ݢ@
�ڃ]��E5�ז�s @0�A��ց�h�&ߴ�ZP�����w�,	u�_]X��ԚC�	v�s9i����ަ�_>���?nι;-G
���|+���{�c�.$j�l�0��tDd�=�W�V�V��a��`y{VJ�����BE���Yj��V�IE��$�ʕ$Z ͳ�)�h���]A�w�`��Ɋ���}-�E/��H�jOJ��H����E�J �^Q��;�����#�_��Z�D�֖x=���LY�C1�q��@D��Y0uK3�ޣ�8���T�B�I��_�J�y)U���&�|�C��*���X��#�)�:6��I0o����1�G�Q<0MMQrh�x�����p����B��z+r˥�G�Vs�-���P���m��M�ޱ�i�$���xը�.7�J�ə�/^N�o�Qfv۠E��l���R�99���{�:�ym�>�;�Wf�����L���{n�W@Űm��3���ҥ˙��-#�v���糤�,�/�䨻?>���2�o,͌(%���=?hdR�n���M���h״���t����F��ψo��g�Vl�߀f��;9.�>�+�\;�F潕bwF2�^D�G�^ΫSXh|��;jd���OY���;i���!F�h����k��7
�BC�%.4���/�?�$Y�cX���]���>�0��V� a��n�cO�,s;Q���ɉ��8�Ҧ��¤�K!'�O3�@U�\��7���3-��tr��:������E��A�6� ��:S���"g`�[�]LEη:m�]S�St��x��j�iGK�hȫ����Y^-$K �Lٯ����8�z��P��,_T�I����N�QC�N��Y.yg�<B͵1�KCl��t�D۩m�I�����^� �R �*��\ߚB���p����#%����6�=Y�a�6U̔�aG��=�f|߱�,�ӯ9&�?�r)�����ͧ 7"ހ:Ƥ��@�-���Y7щ�y�P�������������X,ڊYQ�Śn��g��Au�BYч�i-ك`��d\kt�:�.miJ����W?�Ͱ�Q�����ٴ�fo�����,>}N��������q'&^҇&��8rdUc�cb�m��Ġ����{X��[�AM[_��L��
g���7Sf9��,e;h�O�r�e�0<�g�_=96��=d�}��F����2�>[�%;d���؍�`�`��"��u����Ȼ������U�T.~$�cb�6�&@��e
��k�R�#n-�z���y�.��`�!gU"=�$�s���%�1
�X��&L}v��@�f��!7��"���L(�fK&��|=a��@�s����������-.���7������p����J�r���$!��6?�>���v����߼ĝNpN\�*�hf̅B����\tZ���J��,�-�p�Z���"<�=39�J2@`��C�qF9����*ΝɽN���	z핋4����=�څ=��������'vA8;n�`��oZ�X��
�T����l��:�|}��;��V�o�b*�}$�����i�*Vʍ��u�W��Q�'9�i:5*�C��OGVT���G��Ha�Ċ�C �|~.�dxU�~Ȅ������>��;,A��@�k^|��bgI��Y�	`_�v�߂:�9��̈́���Mf	<3ǏW�8(�Po�o��'v��+��ɍ��(v �ً�/A���2�5��M�9ϲl�~��{�q9��	�bRG�i������Fzs�� �'�b��3q�O���8���iC��\&G�WO2���h맪�/�*�G���*\êy�PY[܁.q��"�߻�O�R��OqQ�d�K�3s��
�w�ͅXW����i7՜UR��UާC$Z�$�s��~Y��f�=��~9�W4�OH��10��%<�$FK�D��l�6:�ىBv�5H�@R�U�1aQ�G0ޭ�Vx�9�Kk�>|M��^��u�$s�_�gr`��ϯ$Z�Z��L:.l(	��yZ��4�k��`���0����8RϢw^�] #�� #�ZXgHTg|k��+^  �t	!�m�x�j�>���q;ЦI�3|B�N8F������n�,Xe B�
	!]�"=�S�!���l
�g��lh�">�(�
M2�z�����:eP�~�#ۑ�������P�Y�*����'�6*�&��R�X {�d��E�������8C ���~��Q���&���7�r�`��/}P�w,�A ���kQi�0��Ay����f����3�a5q	�.��!���V?$�I�V�e��/@D�
g�)��t��SEn�kL�����H�7!
G��)(���C��$#@���hv�Սu��F��G�i^2!�t��<���qp�����R�{&)�bi����DzW������[6�+\��pL>�m4Q�����A�e����PJR��^E�����R8��_�%qB"��1p�2�ʑ1P�����`�Ҷ��eǁ��!��)>`"���N�BTO}�G9�����lə����. D�#��pT�X���|��2xJ��G�d�ʿ�k5UF	s�l��X]1�
o��X����6��e2,2Lq��ʈcA&���N4����,a����VƺF��9�3�=ힵ41�ↀ�N7F��\2� 82�~��Nj��,��{��3Lױ�U�^.�H!�0�y~�r��E]�ԙ|�9>m���E���hv�a��5���9��KB�QcȎ��>�T(D�m�������#�@�T��H���֢9|�v�M��H(�Ѹ�� }���
��h0������D\�
������-�s��\��C_j����j�L�$.@�qL^��_!{�I��W��u�_��U��d��|�
��o�96ef�0\����-��+�����r4D5���)��V8���\��QQ�E�� O��j�]8��l�褷x��`:k���p�e��'���>��2��v{���Z��aimIr@P�M�F{���l��=���T��ȩd��/��P��1�� Ȉ����<�=��n�)A�E��ێ=m��~�Af��~�=�5/݀�R�d�$�K�����\ty����~�7m��Xo9FJ��E�&�ሔ94��u^P����Ydc�����z8����EEO����AI��B��^ 	.�bdh/���k�r��2�)�VA/sd���D�e���iGhl�D��=�ݯ_5�k�A���<[zJ��1' R��@f�&s�>�	��Xǔ�ݳ��r��e�s�fȒ��l�����1��r0��0��0�D8�=a��xвs��10���(�'^U�R��&�Y4ms�@=�2rRΈ�xT��.�J<��߇�,Tl�����:��O��2]"0���كݗ�.�Gq�6��[+#x�N�K�wFͪ�B	�o�_R�M1�;�.e��cg�HI=� �S��|�G�0�q�YR��30�J�S��ہ_>�R��w_�v�<DoFց)��~�W����0�+�<�ސ^P��0���i�M[�W�Sb�8�J὆���4_�IȾ-e�/g�nW�X_� msW��!��sZ0�%�!G2D�Y	��D���g��C1kR� �By���P��6}�m��L�}�	����b�C���6�+f��R)��k^��p�iva���M�FN�N��s泵��n����4~]���kk<2S2�J~���{q|�[͢�㭏����д�*�\��1Κ)!p��-8ۨ��EJ)K\.�����	�mmZ2��V^v�j|��*�������|�|h�I�����H�cQtj_^��ڤ9-�B�#]�1���7Je��	��ickT�2V��6�8�� ����1ڼ���c��y��7���Q�V�z��Xͥ
�˻��{Z�WA�I���]2]�nB �6��=��̬���]����Q���������E������4��0j�FEr��M��&�fbW#��M-�\<������e�#�૽|�=��.O�%2u���i�\+"�B�;g�$9��R��Yx���Y6!~*w��@K�-�8� �j���^to�+onWB8�� WD��h�D�n�G��w�B�h�@�&$����Y=�f��DTnm������Ya�������<J߳�l9nAO�*G3�:d��筙��\s�<׏�K����H� ��+9��6Ơ��r�YRL�ŧ���'unOo�bN�`�[��%:��r�l����_ƷM�5Z1^w��z�^�?r�]�m�%Q˶��FC𛀬�D�K}�g!���ʭ	�;5ҫ����9U�9Cq����aR\�nD�.�� �ý�9H�}���P/`Mh\p�@<��M���8>�f��Ʒ�A���_�\�v�m�����.#�b�ѓ*����U��?���9)����L��^N�>8���~�b��N���"g6D��E��*�*{�NM�=�K'��+]��u�"D&\_�/���_�9�2֡7]%L�E
���\Ҵ�^�s���dmN��llA������Ws��9i�
TA*?�>|�S�F�Ɋol�H&����8-�A0��Em���O��3�	u�7D $���MM7��a�A�%��8}����P��A	��[~>|m�D�%���?�x�~\��Li�0e�/�d�����nkGm�g��:;.E\j�P��&�=�O�ܥܮ&�t4�#����k��CfD����JJ1<�"9�4߯S>��Ppwj�ߜ�ѸȚ�G�Ko<v���2Y�L�l��u��|v��~�3�]�"|&�Dl`���4��>�!�eբ=O.(�ǘt(y�u��Z�w�ہa'�� -�Z�� ��p�v����!�R�KT�u�)�ER9ڐ��$��,yPn��	����N:j(
�raL��}�;Xw�����$��� ���������e�hI�`5��K�K/�_�����D��򜣗�ȍ���$Qv��,��Z�vR�'��#̵X?�.M���t��+���
d�¨^4�7�(}���K�q�)��j�C��ݰ�zJ<�_��� ���Ha
����esA!�X�d?COT�e��ý��
?������Q[A-��טPjkH]	����&��h���JQ�@��7>8�W.���+a��~=�!(uK�2��D�E�≖��kK͌�~K��A'�9YHc���� �b�e�$�K�)�k�ܐn`BT#P�U��4Rg2z��
ov�,]ϓ~��Re���Ϊ��Š�1�m`+�VfD^$"ؠ:�6(1� ���sI/`D�� �m���9Xpc��r]�� I��k5לEz�	X��(AǰXCy�Z�����/�<�,h��9�N\�7��=��)���q����
.jA���A��Z�I�M�d4�m�8@��k�����c��|?�8 xb*����P���9�f	�&�>֗Q�A�\����aE���G�鎘�YU��J�O{�E����a�g�b��B��r%�� ��P�v��m ��F�40��r�a-���@H1�������X*��b���V�_<52�<���%ާ䞻+v�U�K�'gc�p�@j��t8�O�
@�n(��+­(�^s]P�o;"���bR^DI�$�X��+ ��v������������z�/%J�T������t;�'���Z���LZ�5k�76��ǉM�)P4F�,p�k�F����ɢ�PO7�W}���xJE��~��oV�����((Z-�X�.�%�f$P�:F�.-`�1�HT��+�J}cf;�	@�oSȞ^ (3�_)����2#w�>u+���qXA����,��z�������k0Dje���G	�r��c�%,�~]��YB>A��3�T�F]���7�"�$5���X���Y"}�L�e��"� ��\��?X��L�N�KpB��N��z��|�p���n�릦�ִ�&O˹l#��'��6?�������wwa`��A� �̞���ﲇNh��W�^ �W���Á�v"�j�c��r��U0&��5UK��Z�F��dceh�Ԝ�^15Ym��	�)m�!�Ke�	 �*]�
��fo�l��@�����C�dS�1��$L{�,��m�����3^w�Ng��Q�2��V�jV�]|�De��|�9�[;9� K���윘/��e�:�md�@qڱ�L56���i�k���(��q��������{4��m��T��]���o�@�:K7��L��T���~r>Ձ�����n*@d0hPΪ�~W_
~�N[k�n��iA�i�C�K������tl�hݘ��7dL��r��Ͳ��7]>ߞ���VE�x�g���TG������5������q���V��!�L�8�e�Q�ә�ea�p ꘆ�t���e�7�������ô]=#�� �e[Cc*J�&S&� �Y�ܤ7����Z_|J9YF���'����vKjkSUd>ͺ��6M�ڤO���u�{��^�\J��%�WK#Q���I��T��F۽-�;L�.,w��~�����0B� ��I��{yT�&�v���L��q��P�3��<�G�l�>x`,�|`C�b�� �!p�@ls���w�i*�����P�i�.w����SԺL$��F�@e�v��N�W��_�ZaBK�U0*���2��Wz�Ci֢�0W3����'��[2Q-1����=��hi�\���jx�kZG�H'�����6�ႬӼ{�g��9��i����X���&?�E�r��d5���ޔNe���܃��U��!x��ȡ��#t[� mk�C��wY���j��K����W������f잇��Ϩ �4��ё}He���NT��9�=m4	:*���/�M�2fuUm�q��/v����
�SN7y�.�Û�*��Н�ԜX�"����=B��킒�dŎ�;=`'kՐ��Y-�O ���y�f�&�~|�lBH�ε%Nlm�E�,�d �D�`�p&yC��*�_��$h���0�'~�Ec�#��[��Ax��7���Q�m�`����g��L�+(b`�AᠱLN�{q54�����������ga�L�T���ʔ��r(�p�!����JF��w�j�f���Jpߨ�ȍ�:�����N�I%#��7(�7�vH�$�
�� ��s����Qy��C������*`��Oecjl�L�Ҷ����o��c�>��Ӏ�˃�w��:9�b�הٝd��/��V���|�=�n&%���uSHs٬o���g�n���	z��:u|m)@�(���J�wc+�����*��◚:+�o���3f��E!x�z��x-�عǁ�%�%�Ҕ�l��锺42>*�@{��CqoƄ��p��G�����QL�w�&9a�G	�o�~�]=�	��c:�w�C>�m��q����$��4��lY�_C��,���qO{�*+�n�5B5��ח>]���8;^_�Zys���o�/A�Ԍ��w��4��aP�v/A��
^�Y
�ؼ'�M5T	ob1�98��3�;z(B<ֽ$� �o�,ԥ�6VZ�H���f3Q
ћ�XC\�#~��:N\���3�,Z�آ�N��^����o1�-]�&X�Qx��(�ϾҲ�#�1���FɇqSs�g�S����?I�i_��I|گ̻\ O������VE�{�pe7X��;��/T�&�x�q#�
��'�*�^�h���EX�C5^]i}<��m���"*y��u���zG���~
~0EH�C��%�)n!��V_Ǹ0�/�۠��27J��톑"�=�qj<f�4��p���q�;"ZG3�����ʹ1:�'���n�G����D��Q���g,x2%�����Ӌt�a�b
h�4ao����z�x6�`R�LVzM�i�P#F``�d#xhsw�v`�-�����]w֙��<aD-����q�}�~�'�w�T7��O��|���}yu�DG��|��'k��)9#xg��z��y�{�3��%C�w�˥�eX����F��1�O�Tp���pA���*����-��d(���V�g�R��aL��5����� ��/>ѵ,<�L&���0!�xF��Nb��e���M�Gmk�k���W�����o�B�j���M�E/�(@�9��ia�pmK���q>D����F�"�Ǌ�7\\���A�U�Nr;'���m��&K+P)C��,
�w#'Y��ŝ�M?�u��f���}� ���oɻN^M!�D-]}�L�޽�ujR^t�i�"������ʪ�����O�{�_��3"�!)�Ev]%b��! n�K��o&���]��#H��mM��v,��+��*�\[�������gM%�3�J���w�Fy�c��ٯ�S�,��P�Ca��%���_�hWEN�������L�/[`+��n\�A�(ka�����/\��扢��롧g��pij������ԫ~�@ ��́��5��衿��C0�S�Pt���!\�*�B������pm��Hk򆄙G�h����Ϙ�h�{�6���~S}bh�Ԋ�+i��y�i�ŗ���lAm�Ѩ_�<@ �JQ�L/��>��#4����f�ze�5_�zJv@�ܤ[����)�5���uV�a�G��\����DS�;�S\A䎌|���L�H�lȼ��9nU�z�s�̫1J�_ȯ����g�_��(C�\���z���s�Q�Y���yH�%�!���nGr�L�E<�����,�O�(���u4)���Z�;�	���*B����-�:w	�����@��x_�����6���� ���"�ѳ��}+�[I�� �te��'G���9Av��\d�>�����-�Zޭ��i�xp+���m@.�)f�m���鏫�hu�ᐦ^�j3�5�6�g��U}�J>Ʉ�K%:��fV��k��)�9����kf�aOC셓���]ٌw���9�Z}֫�.Ht�c�1T��Sm������cX��N��xTLS�����\-FG�tF ��U�2�u'Q,��@�ػ@|H�Y�j�q���0��n������������2n������� o�ߘ�iG4��?\WH�!���d2����;p����+X�9o�-
�f-"��*�wZ����GUd�V�̭�m�RD�iZ�� 
>���L�J�;�w�K_�Y���qZ��ť��� ��mP���ޖL�2��G����9���LgZZ¿�����"�>=#k("(ѱ���h�	`ҿ���yTQo� �k����!ɠ�#��(5����*�Z�f=�u�(��a��9F*�A̬�$ׂ�{�o��Hh�f%�9�����U�
��$9sV3-����M,���a�����`=�5Ә:]�UI�R*SfD����ya1LAMW@<>
9wp ���?j<��Ho��=/Fb�ǒxC*�^�d�QZӏ<̝�2���&G*\�U0�Q�n-a�[R�F{��B��0��lq�*��Z��6���'.��3�J��Δx� ��Yz��/BC��1�Nk&�T̪���Of�����M(��l��J�;<F�,Y\�����V��*�D+SQF��!�:�i{h���מ��$����M��n@I�Y��)-�sՂ��Bv$O�3oS�Y��0}�%�G������J��?"YS�[p���5�.�A��%1-�V��0�޲AI�8���������x�.B�e�3������@rg��	�~ٸ^|^�Z�/���0Ԓ���X5a�Fm��=�B�ᕴ [��6y4���%�~� ����iR�'ՠ�~�07t�ώė�~�:d�� �Ľ��D�3�.6��w�dr8�Ҍ�h�݌A(ek-��b��xz�k�q�v՝\�b1\��HF�5:�ٯ�ڄ�A�����<WGAdQ���5�������޴l�W���~HEA/�����q/y�$�XY���4L���[�WN+�d�q ���],.��Io��O����L�]�	wj���ol��>&�3MƎ8�jl�Dp���Kh�'Z���2ס&���U,� ��Iߑ�,4u�7!J�N^#rQ;4�n�lw��?�M�KGvv�ZWC�*F0iX�+�ǝ����8�y�&�����#qn��-���φ����龕�%,�Sc!�YA,��M��i�@�<>�QN\�T�m�\�7Ό��`2H�<j ��G�6��Ϛ6�s5s�K������°����`V�H�b����]%�}�?�]��	?`mY��eӺN�-���tc���/)Q�@��E�ZL�d�� :�i)(��@�E����Z>#�1U����B��l� �C]sA�������'!_���3"M�iM����(fzh�Ap4�.�I�����[�!��&/yb�!�%�,%W&�R�>,���<1�V*�x�=���/��2Lݡm�*d	{�&����=&�]������`v�X��]��c�y,%�f/N�����P��C�uU9��@�M��Jh�飄�Q
��y-��@Ǟ�Зg����E�p>f4շ��Ec�}��@�^Gc?R��g
����.��,���[y����u] q�zYl'��4٪��#��?jy�xl�Cڨj�6�L1�a��}(�;��P�!`�ݭ�h�K4�Tf�by�����p�Č��4���\ݧ�uq�����:�F�h���p����hg��S�����I�����^�v7�·؈����j���i�9���Tq/{|n����C�^�{O	ꠣ���vZK�K<��OS�BӺ~� �'��\�/��ۜ� t%	_���{�;�@�D�&�6*KF>���S��-a��r�y���0�������Y�:`c􂮗�SR~�2��7�)� �܉-k!�����I���h����]Qt��YP��9T:�����$ r7�_Iq���n:�n0�DܔZVzr��3	�@�o�0�Z��ʸ�BU�����l�N��_�� �q3R�EB�|�/ҵ����Q��h�f��0xbUc�4��\�1�	a��*��[/! U�u�^�
����G��M�1|v��G5�����o���^��ngz3~�E�X\�Ջ����~r=���0�c�e2���haY���HF�w{c�V�]p�C��%[rCZFt�c�p ��!:Ρ���P����nѡ,lB���Rr�70f�0z�/�8H���j$%FԪ}5���u8��/��Z��@�of���"S3���Gë{�䑜i��|��L�(�3�QE-�%�_��n�<P}�B�����zKwA����sZ��O�?�0�kP�Z��d�Qk}Fw�������ݶ����B�0aR�w���@DÝmH�m�j�[���sѽ d��MFw�M�4�r�-y��p��}��E�"�@nJ1T��'�&�؂*���L�m��m������L��p��e�}ظ�$@;��z#o_���?����,��a��!�ݣ�|����?�	Cn����Fod;�p<c3��,�Ž��g%��:~!��b+��l�����WRU!Y�\Eg�Ǥ�I3ty����I��c�P�
ƖM�9�|�4i�sZø�amz�K7e*&��B�i%�7��	��i|X�=��㙫�ynN��`Wju�p^�Ubm%V6�/�˸�k0<��ؿ���`)�J��hsτ������"B�Yv�5Ի�5�p�1xWYAc�Vh�Zq}����j�5Q�����dblF%(�``Z�(k#".)u��`���o)�f��� .��۠O�}��W���H�=Q���/K�޻�~��ʁ�g���k�V,�6��m�z�ʒ��ƚ�IA�7#~�[d���m�q�s��zp�U^5�w�ˣ`�_�����J�L8�3���xs�U}��@o���C[/0y{p{��-�f,�D��/�~𯶎 s/,nh��5"s�J�l��kK�ê}��L�)n��oT�z| M>_�A8?�~��|e`��������F�=|�*���
E����g1̻�zAn�� ��T8�c ՞,���Jb=	;��޾}��%&�vi1.�م��G����rgQk�3Q�)<��j���F��P� �z:�=��~t��R>�%����ۓ�(��lc�"ʦw�!6�)�BN[�
'�&tTn6?�$��Ek�g�&�I0s Ӣ���`�C��Nn�"��͌���%]�)�*�wȿYE�����=�V�HΪ�7l�i��x�
��L�N�S�J].iu��x^�V�\�_0��>."e~���n�/	!�'t�U`�ש`4�Ɓ�1�V6�M؆3ͭ�h�m��3��7,�q���H�Ԏ���s0E�b�I�x�9�B�I�HJ����t4j!D�F9�k8�y��'Ā�iif/X�	�SNd�"�:��!$�(���8��N��V��_"��1e��0D��d�9B�0��F���Յf>|<�@�;��y�3����i1��"��΀2�t=�2G�z��ҹ�FS�/!�46��s
�Zg��Fb�q�Q�`Q*״F/��'�8���Fʿ/b�m��3\� q�
����C0��
Ҿп�̡�]a���Ly>6��>{��|��Lަ�:�l�(����kh��c�x ���]}Z���&�Wx ԷZs���C�t�p/P�����2�Gr����Ԯ�tZ��:�!�3ǣ15���9�[�º���ѭ�b�)�ǭ��MX)s'�r�|;T���Nw;*�
:���?�[Hv���ց#�?��l�U`1�MGc�
�xW ��1��z<	�M����,����<%���f-�[�� hP`��]��4��L�u]oZ�>T�XC��e��E�+������ޖU��᫹=��kcʌGW<�!���r��㱸<y�@r"��~���h���s�I�t5���x�Vj��y{��a/|?>�ۀ�}�.ħ �H��ࢩ�j�k����J?��:ST6H�)6�گX�`�D�!IXJ�m�����-g�����h��x������cB���+�e�O�)�5G�潖g���u�&�C�$�[�4?#�SJ~����co�� bB���39D�$:?��%V�������S��h5��WO�Y�
\�v����m���#��� �nǼŁD'�hZyO�Q�ȀQ:��\�D�F[4 �C����O�!�d"&��!�f׺�.ގ���x�bl�X	�8���P����Q!�5���6B�b�=�Ѓ���}�H�r��JV��I1���H9��S��z�r��#���5hwn ����8���%Ԯ�\�(	Љj.�v�P%ľ4�}�0ȊX��"��OoZvg��|:J���*���
_O�ﱳt�wO�t	�.���ە3G��mt�0w�$	D3P
c�������9��-AXsy0�z�h���<}GU[O�I�x��џWH9-�_��bn:���[xH?芸{<o��<R�뀅�k����8#c�����HP��Yp�[ ]��_���
��gȴ�9E}Y[ʆ�Hn,	�Ct��}&�Ɯ0[P�o�!~&�jZf����3��������m�	�맓SJM,ɶ�5�!�0K���\�Q�3��bʬ�!4�d o?�WХv���X�U�9�Eʟ�+ZU�^�I�� ��;g�:����E�k��Կ��{�t�1��1UORx��~�L7	,t�V��5�Ev�t9���w���nM�Vݶ��\H�/A��P���PR5�D`Kס��O��N���;y��������.IA�R2L<��٧�9�D���L~�6���|�������f�P�����y 2�����0;BE������\@>Xؖk��C�H1AY�M݄�⼀��)�%K-7\+֓E�X�26�+��T�{tK�j��q5������9�+m���?���Gn�nq���vesCWm0H���5j���}����!:�+������ON�XIp�$RgDK"��/���  o9I�~o���#F�qGJ�吕���6AԠeH��cTQx�p߶�CW�xg�IUr�\}��~���^>@�-�fi�S�:��q�=pى�Ӥ��c�JkV���b�(AФE���}k6������88�S��>�7v9�Ý���Vi�?�K�V�^������×�I%�㵢+��q�HM���׺��@Ip���_�I���m��|W_��+)�=��2V]h��e�[�X}`1��r��7͗D7�0���``�8�b�8v����E��Y�	/����ώ�E<ۯEp�Xe'O���1;R~z�����Ʊ�ӛ૩Ƣ�7+�b�m��R+���$�F���?J�t�ZY�.{%#���*�����=���20�g�l�F��\ػ�uIV9y�H�A�[V�,Ex��/���D�BP����I��^m}ŕ�\j�<2V�$SV�����ٴ���M[l��Tmԝ�\�kp��w����>��٤bK�Zn���_��	����)�,@�<6��D@RKA3�m�t��/�_G�~��{����&�������?�a�N�ع	Z�M��H�H��� s"��� ̉B�w�=�T`yKt������Z���:�4��������%AOE�,�j��x��F����f&|��g%h�H@�����<�-\�J����D�e �wh��������vZ�:tu�u	�+5�av"=`8m;�����-e��lZܫ�l}ՉD��|L�Z�1BSUs�G�9�!O�f�-j�3�mӲ��Ҙ��%P���MU�Nq����3R��|:�!�,��-�b���jp�6+YG,J_�8�ot3��r����u:�<�3;?`�S~)��2ȩ�����@*:���2//�h����8���L��'�5�������YK������[g��fpYsA�5o���]��*+t�cDB���O����ٕ��ZKG2�+j�a�x�[`|��2���0�pBtM����:�\�b�]ō�;����}�A�S�3q7i���kH5�-{X�}����?��#��<X��~�������'}��X��0�?b�f8GD2��~�ʼ� >�,&�S���\g
m)Z��i7��G��$����,R=Z�����i���lg�s�H�>tO��Ӥmo�'�W61���@6'Q����r�4R�_<I�'�ͣ��F��u~��f2�*�|T޽������v�<���2f���`�N��w�6����̼_��k��m�O�q��ğ�rq���T��㗮��4O��N�EĚ����q�#"��ٖ�U �Y��qg�#�a鋙�@�ר�����!�,��t�m������K� +�B���q�xJ%�K��(m�xsR�ӏES<�o-�m!P��f�S�B��9`rG����Y��R�<��爦�dh�ƒ>d��Jo����qCRA��UB�Y�E��5�����j���J`a�rE�\�d��A������ȃȄL_4� �'�1'7	���r�O�8u.a"��r+Ҫ��p'���pk;��tr�~Ħ�h���'����B,R Yq9�ĶW�^�V}��^���O��:QRWV����ؚ�u�	��_D�tiW��~����"�@<a�A�»NM�yt�>���G)� XX�:�4��i��+>�?���n��P��Ȳ� ��n���MP�����R� ���C�����ϩ4�ؔm���}���K_uE��ݨ�΅��𒩌��8;����C��Yg��9Ni*�j���4>;�p��#�-����riGw�S�ƫGWӡ-�v4��B=�<�d�=��7�:��,2��M���m�o6:O�E���>7���8a�L�� n7��k腗�n9?m���es2y]>r�8���ABD:Ӂ7hz����ƴ�y�m�ֱ�|��t�3-F��*�gP�7�_>��9�u��Q�]g]z��x]�9��~aA����Ĕ��W���/nG,�5��۾��u�qt;k�P��O��<�U�wi�ej���?�f����_��	o��%.EXh�Bͯh��4���c�7��s����~�k�J6���F�e���fX�|4���Ou����33I�~�Q_|d����'q��I��Ŕ
���z���M��7�>�8蝺z��`�Lnk��K��\Ԥ0t��p[Z������P�k��������cSy�,��|�h#`�a3y	-�L}�=]��τ�m�>�V���AX�9���_Z�s��!{=&�"���9迴!6��	 ��)�ٛ|�����u���d���y>>�5�es�����+�M��h��qS���v�iDM�Z�g��%�������j���xŉY�<�߃��6�Gu��ʫDT��R����n�ʅ��j���?+�f�>��.T>!�����m	�E/�+/��f}�C	��B�4�w��ȫ����6h��yP>��F2��'���y�p�MP6Ri$P>�f�Bf���H�&�� 0:��_F[_�������AY�N������Pgr��x�4H}�쪧g_�ѐ@A{p���&J��x����LŲ,�Z�M�r��R��6�n����K�����m�m��;à]��^��nm�s�JVshW<�Z�t��g���!_���
E-zS���g[��Z�5�Ş�O��Cq����-F�Ӗ���V.��L
�� s�Rw��x͉�\�[��)�z1R��sj�6M��0Z��Ҋ0�����BhV|u�	�ǥ���iӴ\}J8�:�/Qixh�&����P>l�<u�-���S
P��j ��i���5�ß���A[d����/�7��� �yf~ܰ��-%�.��j.�i���F��0(�U�b� � �^(i���)���`�M?ѕѯ.4��D�i�,�����*,�S�So.�!����c8��3�K1�n�hiy�}f���2>wj^���.#E��U|S5���|�* �Y��1�ĕsYA*pG�}����h{� ��eG;�}�A<	��r����J��9��VtY)�E��_�\���o�-{h�֠^�]� �ڸ�ɖ��Q�DT�#S�𘤛k���;�#����>)y~3&���%�d��a��>�弣�q|��9¢�|�F�}���ݎ0D�VWC�4Z�<�M)��NYCm沨�gj�uǌxt3Q����ZF�gMM*���%�e���}��-�{p^Ҟ�=��}d,6��I?+h꩞%���H�Y7mA�H2����\'���ǃK	Z�m���[%��ܭ�k�/�p�1�M=���$2��~��|S`}�K��LB��oiI_�����+�Q�XM�zvo`	5�Ѵ���ݺ(��@�X8)���S���f�w�����q�t�e^ϩ>��"�<��P��������/m�%C0�2�#q�����lj@�\ X*�Θ L��j�	笶�n�jaHqˋ�$r<V��KƖ�W���W�q����	���%�FI�Q�2�N�PF�G�|f3�h�Y7=��� ������+��U����gm�$a��_�����Z����5���&1�=���(x��۶�����.ET�"��Ǚ[�4?тR�\�El���g���e��2��L�Ug�>՝��j���4.jK����=��)�n12�il�ӟ�zC��J�F�(����`�������ل!!29��I�Uy�u��G8�.YW'O?$E�f2�)zǐ�M�ê�iI�Oҿ|J�,�_�v,#�R����	pd�m�C��@Wc �����tzt��N��Q�y�n_����b# K�\�r�^J㐑�t���y�������2��F�O��*��+m���R��^z�K#�!�,mK4��[Y�V���!R��ML �oG���G���6�4n���KQ������Npffġ��)1�P��g=C>殥���'�?Դ;�K�>|��x�t<�[���Q�լ�+{��hu��h���W�r���� �TcuX����k�$�W�!�k��v�(�����Z<�Z�c��i��b��}�*�E��o�qÑ��(�v7��$���^,���@�K�f�����%�WV���Κ���c�쀒��I!;<0��P1��K�$ъ\tc	(l��3�[�iDI9 :9��Y�p��72.�8n�|��D�İ��q_�ȤF*�Pw!"97u��헡Ⴍ��~3�<P�<N'b�og+���#��@���ן�`~�m�8����ݹנ�r�\�W�Qj��S����EՋ�৸<�g�v����;!�`ͤe4ک�]b�&载xQ�j��ZaqZ��ͭ��y�����m����chĽ(�B0�IK �m_>�`e�C#����GF��f�@���0��q��S��\M%�%U�]�=�����p��b��菼C E�t��\*�e(;�]����]��:YU8u�p+��|+�1AD��֔�3	�V3ے�1D��%*��Z���UTw/���[�������vRO֪ۻ�M� �I�ʺ�  [�r��A���i�.������P+r��HJ��s��<��w�olmZ"��<��w�.)=��(x ��@��[!���`j�Z���1�y��'�:��x������rm7*Z|�K��2NXRKE'F�l��z�|�%��6ֻp����yr�F*�\l�[L�|���-b��֪��(�8�">5A���b �[�E�Ժ	:B����<E��6��	��l�[��m�������'�1���Ψ2)~�΋����(gؓ��H�a�]r֛4���s�ƀv�*g�r>N|��ξ�&������0`���0�F�v�j���;����\I�m��(��r��BԽ�7F�'�
��1�1�YqK�Fyx��2d�N0POf�#��׮��8<]�y�XA�C��(����tԢ�73�ዝ�����(��ò�U�+�R��|+-�"eP� t�ݛ�S�����j�4�aeOmDK�_'݌��1�A���@Ȫ�jv婄Z�r��/cAy��b��7B����(������O�9�3|դ.$P3�sS
�K9R�uS�S��L���dZJ��2AP5�G�ԏ
>�R���!��+���m�j/��_�Z6�J_,�{�?V�	���F5[���M�D=Q��#��.�܃%m�4W�(��1��@o�)V�ڧ;$4�͗Ԉr?\9�a��4���K'���N4dN�q>��n��ȯ/�����v]$�o��jr\e^��c
}��i��,�6������s酫�k>�a5��"!�"м���ܢ	��<'�c/Q5�J��UQf@�������BQ���5@85�}n�[To%�L�,�Xk����{��$ݽ�Pa[ٮ^��x_���Yɘ�Dz��x��^Rj��zo<8��q���\j<�.��A���^�$-q�{�����l [V��>n(�&:�p;K�:`mt�4�&ֻ�9x���6Q���Lv�m������ьp�V��AK��7�P�]�&�8>/����i?͝/��I�]��7kMb`�sGc�W���p �%��wW�eCVG�#��t�x�P/��0�����,��gb�]ޝF1+8l3��Cư�Js�qdN�˨P���q#���LW�ș�N��]�Tt�6�|^��5Y���@�8���\��lX^̓��dň�#֨,��Ь.�ݪ�D��Ң:���a��Po	EI��?���78�3&�Ў��t7��4u�t�=[���kaI�Z/J?�����=�����>6���oJT��G��� ���<}Q���\U��a����:#�[�ڵ�5i����/xf�MaČM(#Aް�"GB��z�Ƣ���`��P�æW�_ć�z��s�b�Dx�8��Ӟ�w���"��/zܘ�93,@�Bv��T�w6	���W��C��%�~�,</H�!�f���^���V��E:��ٕ�Y�ь�\����,�$F4��9Js=�����xܽW
a�%E��5�1��[c9�z���N��s�T��g��]4��tW�oov�T����:_�"��߸}:�{�w����@H���):yy�:�C�P�c���}���s�ˎ����#/�����ZX*+�GA&',_h_�]x6�H]t[3�%�]��c�i^���I���2��R4&��0��j\���,�/�<4Rb&���Ն�HQ��
O�XиN2kpv����2e��EX�\F�>�Tt���͉���J<�Y� ��`x���H"��&�7�q�k2���y�Ů���Q+O��<@���^�� 3�6'��A"��g�R���tY,�ߏ���3�P���3�^LN���C+.��Q���1K>���Ĥ@U=]���&�q�pIC-r�$��b=�i�W�|���-�G>OlP� 4��J�����̇`Ͱ/+���s��q�N�6ZMd�D�r�-�˩����+�\�������q$xsg�!p@�2b'��p��IW]-w!�$��@Ε?�b�^ru6�$�X+}�)�Z��P﫶��[̷f�"_P�r��2��r�\p,!��[Q+sI8܈>܅��PR$�+���Fx��Ҵ�+��T����hl�eiM�l�@�2E7
�4�,��Q�g��-�@�N��0ї��wּ>oV!	����=C�s;g'�t�B�{�R���>��4�!_^m�TiM|��l��r�cA;=u�����M ���[�����H��
�g �|?CT�}=��楓+B&��կ���������Q�j�TE�O����M1����â��z��H/�OƇh��\&�D0�Ԍ�LU���
[5����t7�<�?9���w`ػw=����}<�6�,)��@�R�Ȇ��ֈ���<�R�SXc����ZW��h'��s����]��������q�b�/u�C��c�B�n�첪K�����o;�(�E�������l�6ii��n�|1i�`X{�#Ttk�O:P�V�xC��m�+�����G@\Z�v��qg�;:Ѐ>�Hˁ�)�l<erO�]q���]2(Z9c��mݻ #�m^���	��4�n�d)���gk	.�M�]��y���B��v���g�R�|�q��^�2��\r����|
 �7"
��b�
�΃D2�N��La���CLc�X�'aA8��QNI�(�.��Z+k��gY�Ơ">H��X���B�hb�3�(��8]�����D]�}jzT��2	��ܠͤ��F��Q����Ƃ�9����8z�y� "���t���Df�o�z�t5@���e`R���Mol|��ɵQkJ��Y54�(�5)+��+PEE0ݱ>T0��Bg�ㅌ���A�f��$9{�ϯ�䯇:����MNh�c^3^�g�p���?���b⠊�UӮ���`�� sG�q�n�/G��U[m�k�-?I���U��1=<��C��U?�F�Eh���M��`�,m�ּFC��t�Q��[x�@���u�z�P� U��FSd���\>,$ɝ���бm����~��J�;*��<�XD%X��a%J���җ�ݼ
���(r��$��'�3���9!��uЮQ�)q�U�u�T� ��|���bW��ǕU�6�?���b�7�Ҡ'� *`��x=�0�+�[sYE�"�Wt������I_ق,
o鋭��QDd�+�����@\ݷI��u@��|X�$e�
�Ȕ��a�T�3�P]B��C�q�Dte�6ɪ�.C�嬘&ӿd��K��Dw�瓢w�nJ�vBf��`2O�}��5{��������8�4�gf��0*�3�/B�Vi��p+a��Ͷ��l��\3�>˶�q���*��.�(^�*˓|Uˇ�6�~o��;�E&f��D�ݦ�5������bm��q#1d1/�݌͙�7�𫶧;¥>�d?~9�� ڰ�E�4�-��ig���A�Qy��g��8R	,%Q5fɐ��{�㉷�?E�R�j>�`;�(�T�]�*�$�S�$_���n�]�U�}g�V���u�+
"6����fK������6[2m�CK������,�,�s�����Uw�bo�X9�)�S�e��
,82-�,?��k������D �i]��F!җ3���&꤁8�?�6�k� 8C�u(����@�}C�{INHۧ0��������T��uN��nW��0�-|��QZ]t��V����1!;�Uf��
�^
'�7{����#
Nc��9������3.Y��� ~:�b��nix�P�����2k�w��Ol&�ف��KV|�P�P�
��N!�����jR�F�چFK�Q-�cw��W��*�a�Ȩaq�rr3���l�I��A��-��������L�����`}}�$a:���{���)h|Sb21�����'����Ȋ�G(Q���j�ن~6��o��:x�h>��H�"9U�|Sȩ��T�Y��|稍��]�4m�/�������I�І�7\�<�O�-i�q�&}?E�7 ��H��#��^)���,�� ye���� X�v~��+d���|�rU�h�10���`���Mx�~�����V$�nH{.�P%v�݅�-Ȅ�ۤIј5HࢊV+!�+����臨���OA>8�@�w�6�w5xG���9�X��<�4o��7?�7 y
9sj5���6&fӤ78/����eɢj�T�K��p�>b/���%+X�AdxL�j3��pk����ŗ��9e��Ì��d�-��>�YMWT� E4���D��< ����\�O��ܧ�,�vZ%mqR���\��UDv��Gr�M!L��oY{;"�QʚB�((�4��Eճ��1�&���]�{mNr/�7���\_l���]�"yo��\�����3�/WC��|�x J�y�6�h���?Nu�Kz��PW�rDӳ3H�jH��L ��Υ��	�S�xԓ��Q�=~�:f��{�
�,Qe��7����V��Vp]�R�#�c��t:�����ح��&.f�#�{z�����KѢ���4��Y��T���NƓp����?�q7�0�D?� N_�B��#�o�쪿���1�k쒓s�������4OP�F��)~㶅��%�f��m�SEffh�I���o�I�2_�\���r�{�c���C$ ��;d���a�R޿���~�?�6�ȟ�*�w5B!�*�Xv�R�L��&�0���Z��u�e�S�u������6HtIi�s��)j.ml>�e��&���A�trʯ���3K��K�K�D��؝�����h^Nk����:Avu9�e�y(ߩ4|ɦf��uǨL�J��z���Y�@4ʹ�qU���0Z��EY����ΖL�>/UC!$�{�l8��G��4m�!��
��G��2�0������]ǪJԲ�#�S�Rg\�k��ʮ�e��$o�lAp�69��D�JG���k�n�ϓ� �g9��'��Zl��C��t4��CfXF/�],~��h�RV��H����2���7I�ua_)j�[�~����z���ޝ���ĕ��j������qH׃�=m�t���?�#s��>^?�W̲�؜�G��YM�ts[py!�Л��l�\`�-8b�::��'���d�>U��b�qE��G�8	�m̌���n*uN�6C��w��}=>#�P��dǒ����d��<{�, �٣���"`JV���Fc+E/(#@K���Q�"]�D]Y���Ae �J>��Ғ~��9k@5à�`8� c�Az=��s�:7����7[�7��A�W ���`��;W�;U�K�X'��nZf����.���!��e�p���M��1��]��k��MS2T����m�oX��Wn�؃��!�X�x(>�Y���8�Cd���=>S�u⍬�.�#�D=�$�	���A��K��-@���Y�w�U����u�Dy*�6�dd�TA���D��2�ަ��~�`f�'������A���n�ٙ�3��%�I%G�9^4M*g?��(j�J/��P@*��M�)-��p{�@?��YRvu���:�Tͤm���}���@)B6��N��o	?���_sI��Ծ� ��	yPY�`��_\dDrX�A��8�<��B�~�"���S?*N
ђ�?'�H�ݍ�5��GԜ�Ce\����f��F���yH�j�Xړ�)<�a�����EɾS��\�bi?RG~���������_ƕ���T}���'P�����-�hB�aFf����m���/7�ˮW���δ�ڗ�)-ڣ0���;��c�C�1.VT�c�'��\钬�H@#�k:���i�0�Z+Mk�K�fSg�s��OD�%�7��������ۧ*d���#���>�A��#��iv)��ZJd�Jm!f���00��6�6r��G%���2�o�T�O�i��Vb!E`�q^��&#f�����:|>낋:0!�6���A��?K�ǔӉ �$�_㎯�"��W&Vp�m��c��A�(���ڭ}� 8��__;�b,����:�l��&��aI4-�܈��n��x��T;_m����W�������˕1���G�Rx�<J�Kp���J���y��ԥ8L%t������J~�[���L��֎#!�;��R 7��mT0�R��n�G����-<�Iϴ����^]�%�)�����;u��D>a�^�a���nX�H6��y}��et�U`h?�V�f�|��o~ԡ1�c�=k�m�l�����p���������Q�E%��"| M�
RU���ݓ��[my(�/����5eSC��^���	q힔�ƫ݀������c�EFz���!`K��/�d���7 �r���#k*&*:�
ݗ�I~��8�H	h��<�G���c\��M�y"�oѣ ���˭z���ge�������@"�tk�wb7�~<���(L���ݾ��E����b����f�Su]��k���JG�ɜ�,̋31BLS˖z������sV�v�A�"�/�)C�!�A����ܠy���hvsLo��kZx�;g�Վ�B�/�M�����dCY�
Aܿ��A��.�$Y����5~�l��7���N����A�+m�_�	�!3 <�F��D����oç>*����2�/���Xʃ�#��F��3����-Ĥ�z��S׬/�����|F?�hq>�Y�KJ��AGŶ�A%��ŏ�X����TM]��?�M�>l_�ׄ	;�pZP���O/eՇ�F��2npٞ���L~�b��?]O�"�19��q��P��4��9�b�\��LP�*Q'�V3p��]RQ�k�a�ځ�ߍF��?&���\��&�����^�N�+�"굁:\������pV��&~_+����2ȼq$�.΂B�Z8#z�/I�ҟ%�=�ar�M� agJm?�h�Cf��	C0R��F�b�����w��
;;®Q�x�v�Q ��6nC��� 3\<1��F����b��3�H�k�U�oV���L�5 	���Wˈ,�������7&�yK�n�h�^	�A�i���K��V0Ջ��P�`��y�h
�߅A�5-�ڰ׽�!�U�b�Yg��p�(�Hwh������-���b���Iu���=`�*�q����� T���+şC�oN=���-<~Q�����e�l㏭�F�O9`j���e K�<�qu�+&��Q;3O��5��)�x��S�$J���j�'$L���:��{��`�~o���c�X8��5������	�C�����ZXx�CI�^aa���Y�N�S�v���$:W���@�D�݌[�mH��ޛ5@N�7���|��:���:�\ow�T�6Q �)��R�j�/Jy��}��sb�}D��NF}���ա�g�O��fqN�
�ry������&�Z��ƕ�4����J��� ;�EF[m>BJi���\���x�LM6�8L~	��@?�^�(��v��v��u�;ڪA�˟�!�`}�;U��=�\c����,T�N��n%��t���������j�&[/��6�)���Y@�vȂ*�8=m�&HE�P�,W�l��s]?o�q�,=ރ7�kqM�!S����dV>@+�]y��EuNu�c s�	�c>[/h&S^��
�u�@���H��\ض��P����T�L����	�sWd?m�;�$?�M��6U��|/�����R
q��2�\���4Sb���o�#�5j��r��V�??V6�,Js=	�͂Rw�jD��烉m�5��N�[�����J�6�gI�q݉s�2`�'޷D���x��؄Ԑ�s���2=�eȨޘm��螿F�'���Z�� ��za�F� y���8B��=<�N[���i�4$�A�}���![atz� ���S�a??N����`�(��Z����mJ��:����w�����|�'գ����l_H�젷F��}����ܺlx�\&��K�|���a쐗�G&�)��V6�av������>QO����6����o,b���$r�\%�l�r/Sm�xM�����WC��O�������"��,�w�	"�H�;� ��,���I��!S�HW,��bA����=�}�����T��L�$z"���G��*���9{gO�q��X$�u�tE>=�0L�_�����p�se]�s�~E5�`�=OB�F@TW��~V��9��5�r]YQ%�5��Ot1�7r�T�"�8��Nv7�z�D/f� 4�y:Hh$���Ǆ+�pp��M<-3������N���Tm�nw1����1�a�h��xlqK�밟R��s ת&�e{�@�I�<��C*)�q[�_�63�}���}�}���ݏB>
yƎC�MBp	P�(�eo6h$z|��د�hl�|#b���U	���3���,Nܾ^�L��ģ���W<���[k��Y
�v[�G�m�勰	CK��X؍1ڭK[љ�3��_���o��Ǽ���Gp�gVჂ,Ԯq~�Y>p3���ɱ���Dbc�@��˹������gPīS}1ÿk��'-�P���y>�c}_����\�/�o�}�޵�
��f�/��C��� �t"��\�$�|��"΅�p�����Ш2�:��+8�y����f=>�p^�+RS�
E2g�P㻈솺I_���\���#�}����4�f��w�V�h\���8������"��~ST^�fY��˝�KH�V��qA�hVF�~b���M-x��F�4u\$�*���2�A|�b	���L��h��i�2����w��pLAz�[#����j4�tn��F�����b��nj��[�ZB�������&x�qQ�,���'�]�+(ίK�����ؖY� �(��,�I�j�l8xσ?�Zr���k�Z�P��!�エxK~A��L��#o��r�a�G�FC��°N�Z!�}�:�'X����W_�w�������M�}i��{Vlcb&�l�i<��vv���)Ǔ�D�H��T��[��w�m��'�M�dT ���̏�����'��8�F�~Q�J�'����:�Sup�"�nT�&VI�����ۘ��Q��V=��V~ފ<�h�	bqz��t.���(c��La�Xع+��6o2=�l�W��j6(���"k2C�K'Ny!�)���=�ͪ���S�y78&ga������qk��l���(��o�{�'#��>q�Tf��U�OTܞ�F_�	����~^P�oǾX���h�V�֕#�oi��E��p�lȻ�~iI�\�FK����Q&�c���]�&���?�ܛ֗ŰvŜ����q�����@F]���ڳ/rn�z��?�x��	x��{�Z^NG�1�QmD�>4�PwI8 ���|�걥x�ݜqd��*��T��Z@���:kʩ���K=��a�YK1R��4�C��r�͛bl�ɑk�����B�W��'��ѩ'Es���'��|{�b��=]l�0L�WKP.A�CU�֎�U����C�����g����fjzjW`�X��b�;e/�\�S�j��&h,H1y���O��Sl�tRpR/qx���Q"��O��hTF��=f'���{�3��ˬ�(��-����9������g��qZ.%qJ�DO�6��[�1��(�����WQK.Z���nP�������o�Ř=�b��Fˆ�����M>��hŰ,�������?Ua��V[�o�N����5)�b�İiw�-�r�-�N2�LZ������i��l�/cڗ�@���?|�|kxxL���rA.h�?� &���Ne.W��!Pz<��K��9���n�����N�~_�ԅl`�6�L#�},ȵ�k.sc�S�d;:47b+��۩���QPS�OT��Bm��Q��yP���V�J^����h�C�}W�H%���Ӽ���4)�.��=����QY�u ����Dm^�wA�{���%��YRq��x�_�y;r������?��kp�M�`�~1A�� �فD
��?�WǉN! �X�؍w�dBlv%�ב����I<���a��Ϳb��tĬ�7ZϻkY駀=(�(�\�����hk��e�|��;��2���j9B����/���=��QH��jU��t�@ ����b�I��vd���L`�z�;e����^9��J���q�
p���LE�)CJ�%
�T9D��5=�0��U�A�&Lv�`���6*Y�]*P��y�Di��w�]b���v9/l��C_t�Ӭ
'�����Hql���7iwu8��B����zźYm���B�!Z��޷��Ф"_�a�"K2��#��"b���X�����XM��Ta�T��$6��X�1OPG-��2����1�����Y䩆9�D9�
&�]�^R��j��-���ǥ����:���ؽ�3M��F��.�ej�V����w�}3�Tl6e�ߘ�n;�ͤ���kXإz�N�����[�Z�^�"�P���Yh��q��BP���'�i��!���soV��?6����G]`�ݪ���q�螚{�*
�N�]p�x�,��ł�t2����	�n��/����`!D�c��qԖ��բ�Xʴl�%�-�|J�9&�Vfc�tI���a�v�~���,`��-t(S	��I���˻���E�Gdi��5˗gzE�J)�_�f�Q��ON�L������-�i�0�l'�Pa��Kn�v���n�\ӂ�Td("U�WRG����T�Ua�i�aA�f�%Bt ��>U�lVѫ���Ď{��>JV�D��o�PU� \��.Ki�o��5�\�ݏ��_�����"��wtP<�5_c�Y��AD#�H#{�=�����>g�P��S8�4�����q��	ꈬu� ��6;�n�?��Ӻ4��3�(џ�p�bd�{��<���s]bc]CҤd:�t2��B�+�Z�w,�Н/&۟�^V;�$�%�D���t�����]�~(�0���CN���56�$�7;��6�c��>�\	G�/������	�D�gR+�}>��@k
ϟ��_�[�@BDaLP.Y8�<]���^MO"UR%pc_�����,�'I;HǢ]"�Q&@_,?��)(O��\��>�`��Gj0��R��iŅ��N\w�C�B��"�$�-�6�l�W��u�V�����y��pY
���ˍ��xB�+	��#~��Y��2WŚ������L���}EM���h]���E��*}9�JH_����f�������m�k�7��	�S�@�*�h���;�9�����P���n&f����Na�I���]Q��*�F`<�c_��r��{u�~�.���f���������f:,������s_�K�7��3r�9��c�}�+�a}3Tu�^��t�6��_@T��]FeS+�Cu�pVY�+��A`!,6
�pQ��TC��4W�s�
�Z!�F3a��´���.d��{�t5C�r�n+�SJ��f�ʤ8|��\2��eyD��:iA��[H�I+ƭl��&аԅZY��|�3��� ٺ��
�#�ի׀��ۡ�z&�Z�j�l�-��H,č�BF�+S;_y���e�����L�D( ��j�l����Ʌ���;e��?X��{����Y��GL�m$�5��"��2��ʒ�,E���2~r��B@�Bd�Bo����3�ro̊+��[��zF�
����!����y��
;�4jV��Y6/�rh�U-�7�Ji P~v�D���G�%q$�h�H�%;c��6�vk�@k��qH���#H��U�mV��'bKxf�'���?E�44�6	^�}��`��>��;N��~CK�o�%��t��Lvu�^!�4�Q��&�Uʟr��[�}�.5���3�����I�?+�X��G�`(���eQ�%�����m�4�/1z8oj�H�2�AX=E�SG�7:�)��yݦ&w�ҴiB�`�S�v&g0;�t�T��/���Ûa����E�#+��\�p���<���6b�g�o�R�=�����\>����A�7z�aO��en�7�$+$�<�W^�c3�������?0�Ht���9�W�%��`B�N�n��{;��IN�,q�-v�F�	�uH�N%�h�G`b�i4	]�aNqzӼ�摹��(ӡ<
��"-�ڑ�3���MsoYO�#�~ҽW��k�tU��81����|����Tb�E��p{�S���||
�:9�����B}s<�l�ty��%Z��ZҚ��"E�����7^�F�~���n��ӳ�և��Rϑ
3>S��ɘ2}9�s8�O�i;5_&^��^X��o������1	�EMR��
T�l���a�w�5�F�Y��ʥ��R~���)�ibY䵙�!�r}1�i�j]��&��[*��ܶ�_Hef�t^�øSrQ��ۖ6%Z X�J&�	_َz��t� ��,�l.(s ���b(�9�)��kѽ���|�,.�؍��t������j}��p�|��4��,p.�h[�=�Y�3I��d�!NX����5V0��ĸ�c�J��h&��Z~��=|�-���2�C��^� �f&��`��B�I	�g!��u��nf|�e㻾e�lȟ�'ɹ��&�cֺX����<����3�qk���;�"�]�C�<nOu:*�H�%��l{����6)����CnK�G?$j�I`�{�ޔXi9��I�>���K��Χ��T)��������fl���zZeq\)y������V�:|J��X���L���JImY;�����N��'��q�0$�f��m�s���`LB��I��`�T��tt"@xs���Y�职�[h�$3M��Bje�܀q{�k��n@J|N�\9�9]��I3�^����"�+�י/�Z.{Y�q�`�J��l񸁼����F�*h"�#�:�%w�L�U�%b��o�v^�t�~"��,L����7�vo�q�5�֭�����~"�?f"%�zˋ��]��'���eil�����)�5��ż��8k��+G1}�T���L�wx�tx����Z!�BZB�c�u[$��&zq���]�AOD�wz�57��z��Z�
��g�n�(���T��}���$3���SO@B�Df=uz	Bi��`\���d/�"�8����XP�5V���m����?i+ˮ�P�|Y}�?Z{zS&��7����Ƥ�VXu@��:E͟v�����W[�dJ�3�D��dp*��/vV�?�l!g�u�|����!��'L�En��ljcB���@��iF���B�ȳ�r��n9�]�E_xJ �`�V�,�IJI~1 �>T B�3��h"7�VP�x�G�"�	����U�%�hV�ZCP"!�jmҕF�/�|�u%��J�"}T��)(�;�zA��	�؝�=�ө�����fUҴ����$nRusn��29~'Y��%��5���/��?�6ЯEW��GB���U����1����Qz>��	� ��9���Z��'�)(��0�� �?�����o@���� �͸i��$`�#���*�H��~ ����CU
/p��0nr�D�>ۗ�3Vb�N4���I��d�p��z�$ޘ�,�oss���j��2�~ �������R��{�t4ig�f�
~�E���Av��/]3)O��_�����Ҝ[�Q�f�@ �N����z�?�]��;)g��M�Z���pP(�:۵��S�V$K�C�L���Z�~��	�Q`�%�j�U�� 	���|dڑ>j��:fQ8į��+<q�`w��Ur����n�|~Ŭ�����4�@܈e��>�^��} uԣ
�8v	?,ס+��D��M��>[������)�lSoI��cV�HyT��[�P揌E����qg*e��[!�&����z���r��-oŹ]x(䖙�PǍ$�s��������&(e�De�X�5l���!M��Y�V�}����O��I�eXza��������%�7���AK?=��f L,Nm7��V;�
:��;V(EV%ݰ!~P1~�&M�}ZB^n��D���OrJ$$K��h�\`�̲<c���6|J��̙ؒ6�%��ms`��lv��h���v
�!�8��g�kݤqt�9����'��.���7��e<�*�P��H�[\�i&��a$������7
�;��Ź�����@��5:�T0DTڒ:A���7��X*
6	{���CW-Aǩ��^�����Oޗ\��@���_z�$��5H&ӜF9W�_^��w��$鰊���/����	�ۘ�+�.��;�r�N�-s2a����������eM#�Ή��a���u��x��+�"��Dt~�إ��&��
��'zC�qtzuX�AB)ܑc�n�~5ϟ-�ƑX<�(�j2��DV�̟�o�����9ʍ��bį���-A�o$��T�Ч�Ǆ���k%<����TV�A��Z�{6�)~�,�̞�"����7n:�ʾ��[�_���xD���v{.�h�e�xݘ�闬�=!c�#�R2]��0x�����IuEIP{�|�G�&�A���+-9�>�3;gr��M�x�%�!¿��O�u��E6k ZE���Y�o �z}W��g,��;�7����䏢�~0U&g3�p��-�`�
~�D�i�H$�HҬ�֠d­���7�M�_�w�KH%k������4�E�^N;�=�x �Q�A!���l��G{2��ۇ�\p���DdmUL�Yc� {\���[Բ1Ԓ�"x����������wR��k�*��te%����:'��J��AL�9�h�>��pk�:zn�w��ۮوr��ao�h��Pd�7�Y�sE�XFQ`��a�!;d�.�=ﻘ�Q�ɧz��3�w��M��WD�,U�a�xq�% {�_��O�4�S�3s��6`CЃRi��i΄��$R�Qh���4u��i�ݓ��������
Q��W����B��Q4� �	�Z�SR+�w��!��d��l�?���$p��`��<*J��IWd�s 0�g^�]~`2B�rS���<9P�_lg���"�g��7N���HF���1�,�;�^�eg�X锔���sY^�껬`O����,s�2y���~�HH�	єk��|��(?�G�+�3�]�o2g���x�ύ�� |eLu*T"�x�
�Hm�dj��yk�V�pu���n��7Jz����v��<v١)�ۺ��Q�l,`s�>�u� a�1;v��BY�W]�vD�Ɵ�N�u3>(s���;G�,L��ڍB+jhe��4��v��-�<�LL��T}�KNys�}�=���S��;�c�y�mΑ��[
m����aԞ��R2����>�A���b�9z��W���Ŀ���
��S��Q�M:Ho��J�Y��E�V�	���I�n�K�����p�z�d��H�hH"�wA�����:��eB*�|���	5&�Uކ�%�xE"�P<�V����\ Ɣ�NV��zqRl�L�U6�	�= ����/0ѻ�>���ZIU`=�����=���̯Sd�����0X�J�
E�d��k=Yf j矵Q;Q���R�T�=����$SLf�X�Z�o/LӨL��.fF2��^�7Q2��⣯c�B��@�@��s�K J3��~�PQl�����!�2��[��dM��,
�/��5DK��^*�-���^5�˃
9��x�y�X��[���Jj�~t�(�7	�ro^��9���	iz�s�Y�+Ѻ�h��ǹe�������F,���:�C@��u-lf�Dҗ���QoKc��'�U���Wi�pռi�V9n܄?c�V�'������%�N��@�tF��q��!�6�BǢ���rx����A��'�����KAY0��	���׏ݾ8���	p�Ӿr�N�~M�P`�t\�?�2HK:}������ w�&wa�8@����K�+ڲ,RT!����4І��e�|���:�	v�8|��wm5қ�~Fo
��%���_��&�1�$�#���k"�Lr����Kn}Hu��3�Gd�{��V)���b���GbQp�g �ɓ�����P������l"27-�QI2���#�S������~��X�� ґ���k^Tf���J�&m�W��@�?%�wSZ�e`m$�"/��_�ݜ�(�^T�[�|���o�k��F;�:��V\ (�zX���.�2�������
aB�u]g�Ky� ���i#��:���#�M����R&��͞�5lBk2o�p������~u��To�Ņd��߄9َ���T�=ڨ�/V.�O
������g�2ŉ�Zv�냧/�M�tI�13_ (�����U'2栵��}��k\m�Bk������m>�a8`U�R���5�*�}9��ObIE��<�;�(�0�!�\ұ�.���m��H?��kw��:K=#�8$:��x߉�z�S*�>�d�5�΍��<�3�QF�.:���4��$	Sq�QN@��C:f&�_#�D�H�l��d] ��]�L:0��`��s;�E���F�F����d&��SB�h��޼j�+3����_�܋AX,7$�+t�x�4�?\\��� #Q ������AbC`DNN��Ԗ��؏uO��7GM�I�bq'�N�Zr�3�Q?AD|� b��V��0؜�yŠ���0-�ep�3����։��<UTs�Ep�"�I:��Ϭ��Ա]�`���?�Ff�g��m�Gθ�5=���9s.�����+��p"���0���!fT	�Q`ušvF���t
����'��w����+�H�����M����-
�T�K¤���B��"F�\�����@f>,��?s��ղ�r��yP�:}m�i�7�Բ�#5>�Ȭ�̑��'D���L���dSlj���)c'�I�r��ZP�[�T�5�KP��V���z~���6�:��T����jݖ�h�=��^V���W���d}���Fdg˚h��b�K��<�MW���Uaa��n�Ne�L�J�%�-����c���9��{��KL
'���`Ϳ��)i���ȕ�p�*��XI�87�.�J/�l�E������9�_��u�I��v��K��|M�VN���j�F�q{IZ��I�G0}��L����p[�:^�=�y�V�P �8Jqo�������&����˕fDh̼��t�͟%2��ϛ&�
�IP2p�F����gkIX���Є�z31��kL���?jw�9�Fڕ����=�����	�m��܂]� J�JZѮ�K܁�ֈG��v]rPq��/S�Xi.�}�������߮�!�P�����xs;_�3n))S��z!�}2�:�!Br����aPԚ.�ϐ�TQI��EY�3T��߉S'ۢ���RYݲvw2���:��fd�-���>8��Z0t#y5���2����|t�G��>�;P������Ab��,���_�	�̆q6�������h<��]p���5��_�?�{�CgX�߱{��a���^��oN���e`�9ȝ��6K_%m�,���F�F+0�Y%i���JqhᛲL�c7����GC�Uox�lE�)	�v�H�i�uLg��!���}��@��nX"�*˼WX�k0��^�M��]ސ��jN,��~�D�gC8���`��H	��A�0����6���g�tI߉�a��:�Q�?��t@>��,������D|�|3Y__
ñ5��؜�q[̸��ܔ�����Ä�q�`�vC�[w��#K?��5�v�����	��/!Ul�x(�%��Ӷc&jo����|R.!8m,ԩ�o������<�{�(�Իznд�t�+"�t�����??0��jfI��	1�ɟf&q0�@x5�ၙ�a�"AP%�n�Ma�6(�G#�!�֌�ꃴ��I�a0�7{o��aؼA{��kGC��7<l7�jWȨmF$3��!�t~$�&&o�ÙNjJ����oS��"���=�F�@QUF-���
��@rcc��O�v��@O��Ua��n�=�,�o�Ґ��.��$�8F�����
���ҴS�Y@`�
`H�: |l=m�vw ��P1I�N�F9�෉~&�&8��EL��f��+9o��(Bs�f��6GC��p�ܗ�b�y��;��lT�D�����Rh��wT<���b�>`B=X��*�8f���I���l.�jO�� �����UQ��>Ǟ�2��`N&_e_� A�7�$�N�G/�e4aKJ���VO��t�	��Q�i���)Ďq(D���1���wJ�:����u��kh޽s6+bt�Ww&��d���'����N@o�*Uv�f2	��Ϭ]#q6"$g���Y�:g������鸇�w�P�;��h*6��K����zr�"U, �[�R|G�+]s䰸�ɫ5>Rpf.�%��f�[I�m�����D���#�B���7;��h��^؝�_~Іd얿�?���>��wB_�2�p ��,QG�0:����HJ Y�����D����D�����5�`Iy���ZI�x��� 9h�氖�F
���L�/��՝Nls�ۥ`QXVؕ��t�R�]Dq$�l��5���@�p�iG3y�Qk#<��C16�r����2��Ǡ���j�`0�Ǣ#.�<�
��Z�=%��}���^�㱱;����o�mS�p��Ft�J�c���DWk��fN��Ý��˗��rKH\�M.DU��Xւ�������������!��_�啊.'���,���<�\!�����<8g\�&$�]
��J��#�f�B1e���i8�I}�M��Qi�3�m�rM�,'��vt�*�m&��>��]g���AP������	R:\ik^?T|�͐T]�T�Ȍ���Q
�%.ig/
 ?D��N�%>>��$x�}�]���p�]g}�8���u^!/W�3d���UP+�)�Yl���t)��6�.t!%Q�M�
6S�0��x#�+�������CC�1�k����b2%O��ggF���]yٲC��	t��Y�fb;�hH˝QW�Hr���y6���VSa��$~��A��jk��p�����J��"[Rs���_;�w�ُ�iH=�?�q̎J�"gD�.�P8>�0�`��:�U|+z������X)LW�5���A�&���:���&�YF���fv��J+V�)��0x�'1�JNҟ�	�f<���][���(��Eܯ��4��@;g5nQԼ;�g�k#/U(C�ނ��5�� Y��S#�����^dd�d�Ϸ�K#;���=0=�����E6�[0 ` �O��]��ÄD�E`Nd�w�����qQ�o��Goݩ����t�����"��
���Bt����.��M�W����kٛN�.���M8���t�@uP�S؉:���fy1���ȁw~M�Ē� #2"��)PH�
�V��,D�y��-5\�El��N �mޟVA�M*�WIw ���?�9z;�[���tJ���U�_g���CB#u0N��0�ki�x��4B��B�"E2����ubW�~u	��l�y��8X�p �@9g3��/�=����,�)��-��P�ǃ3���F�b$��/����l��i��NX`��,�b������D绞��C4�E$����a�I������X��^�?�1H���)PB���|�xY �V�Қ�y���PD�1�VY9��y3~v� s\"�CX�0*al�[���Fw�p7v^Ž1h)��
���P�e��T.͕����>ۤK�H�M�Ε���К�͇�h��3���>f��Ց�DѽL5�-mn��8�^�IGS�y�W��t�pz�J�]�5��k�̓{P�t5c=�i����v?7��:
��p���u�p�:4�<�ӤP.w��H8��q&@����S�q *��e�Q���Š�hU�\�R �w��F�&T���{�Ɂ���(�Vz>�ai1aR���.'0;yO?5.14#��S��#?��2W��J֐�i΁/%������,"��Cɮ���£�fwE��ztSC!����mr�qwƏ������$�wiP�>ġVJ�B+E�;0�������酂9�ױ
���f��<r�C���}VT�1C�H��U������J��[��O�O�"�UӸͮ�M�o� �]� �˰8�$��S�Ჾ�i!D�(u�(\V�N$�1�m����$���)d��10��	<C�!ol%Ff��n�~Tq��P�ZU)�R��l��\�Y��Z>�%�o�R����чV���[˃��!�F�\��⾭�}}Z)(d��P�cp�.� 5���ɫ7ט�mQ���Ns�%�2'0,�M�Ї=�U���	�%ou���c���a��YE����H'҂�_3��o�Nˬ��VI�;���K��j���"d�N���؏�O��$��P�6׆;Ź�r�y����'�#�N�iZ�Dٹ�KW*������)��RCBk��(��	Z��zМ�7R�2r��S����5?JZ���s��Z�SٔX��tv��"���g�0���Xc��a��u/˽aS����UB��q �E,�;(�{8,���\"�����"��et��{٘��$���^}��vY|�,[ &�l�%�Qor�$LX��G�[�)�!eҮ�U��`�k�<G��)i�#l�ڛ�Pt~f�Z�>k��]����.���QQvV���gX:�s��N]�8�AH�N��*�̆Fy^)�r��El���s�sVp+�������������vOM1bA-��E(k�jٖ�dpI�ߎ>'���1��{[��f]�� U�D���#x;u�l�X�x�le�a~#n`ї:�ؚܽkL׌3�3���p�	e���∼$��!_`d�`����<�,�D��Pg��Gv�P����[�
iB�4tT8���#��O,�e����2�m���WT3�%@����٨��M������~>��� �	���u�R�i�4�.I#E�>�U�Jm�j���(�6i���L��z����j�1�Hn�o떧7|� UK��Ғ��mW@��{.�!�ؗf���a��Π��~axV3�Q�Ik8WkM�O��滿��*M@frqŻ��89zD���,0�5(�N��2PҦ�d�A�j�|�[M����d_��^_%ߗ���ٛϯGhR���o	ש����*X,	}WӋ��'I.�_�r���.��	^�FXwOy� ^�T�5�4;������s�r�X3l1���˅����³P]ц-fmC6���&���Z#���	#A��A��ֺ�|�L��)��^�nP��?�����fW03:X9��VT�q��V8)��~L�hG�sB�;r(���¼�2#�ǽ�P=��g�Wa�/}B��)-�r�U�1k���Ċ!;�9+ejV�V���Z�xQ!Lf�9%5J?�"i�j' �dZ�y~���9�`�c�k�2����0^JH��t8���e����\S: 1r�Ox���t�AB#W�!{F�T���Ї���Sҽ]����' �,S,)w4=2��:궿���IЊb�ٔ�:�-9�O�$`Y̷|̭�bV���&�L��+e`�|b4��Js���`�Y�/ ���d4����� ��H������OS�}]y�~�kn���ҚC��
����y�f���M����&�����/ݶ�&j}�F���qs���'1�7��Ʌ�A�k l�[8�H+��f>���|iV?�T����M�w���L~ީKU��[��؃㊴�������_P���S��"���V��z·��ˉE���Q}���f�Bu����q�ƮF3Nt ��� %1�	T��T���}#�7�k��@��2t�li��z̳_>φd�˃I9k�:�E ����./O)���ټ;�#��������5�(�č���T0|,�A�	W�3���U���L3���-�����ƒ(��P ͵��L�2����y�,�^�!����
��(��.�h�d�ѐ<�zS�c�'�7��#���SA���v��A��b���B�K6����k���ۻ
�?��TT��:\`������,+Q��yq.�]���W�_7�w��6b#Z]T�����{�e��m����9��>k"���U<o��k}@���8 ��.E�7q\*�Q���n�z���{��F�1��[%G<�@�mf�M؁��=~F䲴��fB�Gr���&�����(�iY}��s�?����Cض�����s�6����ps�'�p��f0O&7/2����ɗ0t���u4�D����Wm���"��T#���!����6�>�%DhA���a�B���l�1 �8`j_�r���/�A�RK������/:u���2�i0���o3�!����
���0~��'���(����]Oy>e���[֢!����Փ��EwtAr�Mu݉Lax��{vU��E�0ĸ������!BzA\�m��{��9ђ�W
�Y�S'�5k�53Ҽ~Fɩ� r����ϸn,u��]�v8+��=_D F�f��~��,KI������fi2�J{��9C߲��-AZ�&AJ���=Zl�3�؂��.�A���^B��
�C�k{]M�L���-hiXf�.f���,����vlB�L8���ͩe�tk*��f�$i�[�/��a��#�S��}���ZA������W�o��=@�����2�e#��Vg����y��:"���rls^	Q�M邳u=.(����-@RZ��?e�ѝ��]m��Ԋ
u��x"�?�Cq��vB�y8l�����`�����I��=2@�;��Fv�=�#*�+�m��B�E=li�,�$n�o�n��g�0����`���[���0{�ze��A���W���@�ۢ�D��!��n�{�$v���ԧ�;dʁ9sx)�o�G���0�V�x8؎k�"��S���R�-�{f�pv��fmwx}�A�
��E<+:���#HE��w{�|5d͡H�� L7J�����W�ׄ�M��ڔI�mZ�!����],߈7��>�����jE�8�`��x����#@��jT�g��4ZN)HK�{Z?tɀ���T��f���OnM0�J+	�#Y�.R%�
w����wn"!���+,
8=g�(��lSU��l</���ܬ r�q��?T���Q[]�ͰA�(Pa�K?c��a���h��f�G��n�9:Ԯ_+T���1���wt\Ft %1�4� <m���w�(]�{-_�<ϡH���Q���� �GX��Z킈���Tc�6�a����"�xqM�g?��Xm
�T�8�;���
��HA��;�:ϮGH��u�*�B�k�ˋ�W[�SYIt��k�K��q|�A,�*�~�����n�)�Kov�ZR�y�R�0�͘�Q�D͎����a�mŮJ�*�����'D\��j:I�z�0ow� 7��ۥ�+�&$�i���&��K)UI�=W�+�dx�5���%@�nXo�7#o��"�����+<g(U��:�qYzC�:���/�k^��cq�$1�q@*�(���=�/o8�ޓ�T���^��^/��f!H��D�UZ�vۨy�؛TU!5��>�)7w��қ��gp�-2Iu?c�����Ҩ.�s���(�N��˭.d��: H��	<HZ�&H��c�Uh$��ࣧR��L�q,X*9S
=�X\:�n���]�3���'�<9>ګH�|�r���,�}�*	�0es}2h�����D��6�~���[J���*��h���-�խKk��M�Ia{�N�=�;�y�j&fQ��x^���q�=�"S#�U��0�	�Y8�g�[I�::�QO3nZ��s^�~.��v3��:ƕ���p �M�k5).-~x��|�_d��ׂM[̍2)
@��:����y�g��X��R�Z�L����S3X���Kj�	H�Lᖆ����R�i�QKhͭS2佟1�c-�g�J�+��F�ݚ�`����z�h�-�>\�����������,��`\0��M	�!�8���jN�ӓ�8�D-qP�_���7�5�Ŀ�F�H��k�����$��~K�}	3/x6D'�����d�T��W[�S�Q��E�'mS�.i�6K�}�~"�A{��X6��e���(�Z�{��(���;6�X��� c�Χ��� ����-�*�I�32�xB"���2^�4��`�q��m�-�b�mqw�f�i����>�*Z���1�v<�����,<����-L���0}^�hŒ^�eG�]>Q#�V1���;��$�N������<j���MW����Gp��wp� DT��m�	h���JO�����8����>�Ғ�),Ups���Yً�˰m�2��׸x8��ӽFmuZ���ѱ�������Z�6��ƹ�w�!�5E�c��U<�=�.t�Iva�uwb�h^6uJ,`Lg}���>�����
k�%$�ٸd\@Ѻߥ�j���W��8,�j<˧�+H_����ۡ�E6��1�h��.��
����_7��%���g7c9�I6�fQ��n���l�m��,е�A�x�~��/]{��eE����m�ݙ�6,׊���L�m@ㄬ�Ir�1ᑑΣ�XU�0���F���X�uVyS}�3��*	���6h��7�b"C��vLN!�8�3b��(���q�c�ʅƤy�������LGti��bٳ�\�'�-�(�s��ǯ�#c�?5�t(��6*���US?�5����{���7�H�1Q�eش� .����9�&ЮiT�ǵ�q;0`[���U�r�����`���p���"���w6R����Z��+k�4�|��
#0{��}���-�DLW���w7��݇GfD���a#6}(�Q0�0	 ԍ:��DQ��C}�9�F�#���<'��������/�h��-^%8.+���6ZRޱ��k���9�!·ܦ�Fo���Ϊ �)8�#��{I��m��`�������<�gR<��iE+G�$#�8�2x
�*�Hb"`H{�Ej/+�ډ����X��܋u��ѭ��b^]�1iW�7�1��;h̓{u��s�������|:�ݘ󌐯GT�f��J����W��ck>I��Vu�D4;@8\#SiZ�P���+8&R�=�*1�_c�X)����Sf��n�D!�A�&2��Ա�{
{! �=�{e�X�Z��wK<]C&݊�2ׅ�UUy��l{�hIؾ�ǵ鄥��v3�+�E�?��k�2�J�&��������ȕ�Ѯ!��t-�d�jWDyη�Ӿ����U�i]��ϵ�k��a5��z묶��GT��ks��La�TZ��Uel��ځ����#s?3f\��5i�,0�Տ�͹}�H�h�����KckpRP�a:D{�����z�p�4m:Iq�#�kMe�?`�V�W���@�Z��㛃9�$k-�y�Q�d�D�p.ce0��	Ą���
��Ӻ�Ѡ1���lœ���Yoc�P[��VE!_��b�<_�fn6տ�K��nj~�X�*��̹T��}�߱m\�uaj��S;zP��n����p�k��T[�2�LF*^;�X�oE��,�Z�Y�.��3j�[�/�4S�&oLh�L`�Y�p�~���!ү�`�k�̽9q.��BCv��F�ͺ>Є����kk�l�12�1����Bo��P�ǀ��SPP��$e��}�:��j�����w�P�re����7=�H�r)�X��~:2[�Tۅ����_L�_ICbr�i=����%�Ί#*���}ϥkR_�J�÷�;ɏ�5.���"���Y��o�r��%��~�.�);(	N�J*�"[�O�Xc�����H(!G0�����#n��w���J�%
�M�=�&2��������Y���]Rp瓼���Zw�8�c�̆9c$�C�D��5SP�J�Ƽ'>�rʤ�xwy�H��u}��o�����H��	ꁸ�w�%Xe��nۋ�
����ϒ�	�O��S�Ŋ��kL��8�HL0E����{Q���sK7�V�Z�^�U9r����5!�Z��f�����#�ls�*���1�^a�Yi��yb��N�GWwW�v�`�^��S�#��G}��E
lW A;?�*G�տ�q��`� �0����u?��]�8�T�y�-CYӉ�~�p�n�:���H�D��~�6�ٜM����Ů�$�9����4�#Q.�<+�4M�D���ͩ��$(8����eO�CЭve8kQ�i�}5���&��^�H#���O��*1�$�N��J,F}�	������n�@�R}&z�&�����`�T���;�e�l��ai�Z��'�تq�0G�b��u?�2/?f��ך'xf_xo��6(QhX��|Zϲ���<����D�d��8v�n�tDT�e05"?C��a�[I栘�V�E (�0�3	��QB�2X��m�@��Eg�"PĬ�b���E�nY���k{T�y+ME�u����L�%���L]\������vsj��C���CR�~Ny<�W�m=T�ty=%��T��5m�1/� ����¯��7Ҩ�۲�� :h]��H
:�>�SR!��s+��=���A�@��~�g���g��K�6����I�uTڡ�kR���\�d�{˹��}+�h��{�(AQF�A���I��S:Κ�i��ODC�lݪ}� ��6�G�-� Ϭ��P�i1s�"���s���4�s�W�''M7%�l���Z�����{�� gF���L]��`��Jq�-a۳��)�:(~��L�`W�Ry�c�݀s�A�{%]W(�C�����F��ا�O5Lo������1�~?����4��s��!�Q܈I�ml���	��g4ً�G@�b�M�_y�h��Yͧw�����׎����=^
";� t�Mm�Q�/�̍�ôs�h.̄�W��+���g�-<bԼ��"yZ����yW�u���dr����E�ρ�� �Y�|�XOs�{]�9y|ܔ1ee�� �5��V#�J��	��*5��Y�9�4��6�D2�,H�:�������k����O���7�(�v(��B��V��a|��#�
.f�o���( I���ı��bV���M�(��yg��EA�T\E�r=U�7�^0Sz��JU��;�<���|�N�U襽�Qk|��c��#�$����ʟ��S���1���ǰ�f-�A��[�X�_���Js����g��H_����c���j|�����Vt[���{�����f��Q�~W���ƂY"��Ō�HS���M
���)ؠ�{jP�KF����PT�r��\���E�Jת'�Ԑ>L�EH	tFfƨ�yl�U��I4๘h�8G��*zp�ϲ�n4�o�46�Nlk}C��й��[F����a�"�Q��08lS�#(t�_*��E��Ѧ�����Wbi�\yD:R��h1�U�hT�i�x�r$9�4�ED�������)��GX�l�M:�]��� �E�&ș��u�!�����5�������X�Oy���|�����]o��q��룧���R�K�6��Ar�h����&	/p�^U�̮6^����܎5�N�'�E(�h'n�{y���x���E�����D����Q<���b�!����S�%�]L��E�[9�"�fV,�6�6�"� 4P��$lX�{J�M�V��{�xg>�)�~G�V+:T�S/H�pU�d�hR��$�6|�L�5��x�#�(F.*νV���Z�;?�mg�@3G���a�3�C�#�Q�ȫ�Am����_�W����R%;�"�{�\��#A/�#|��j��l�%J�2>u���t mm�BsfK��5E�-,Z
�J�������9\�b$q+g�sgSJz�l(&�∌�p�J�Wa��t^e/ �9a�3Q�6�����$.�1�P����럶��ԥ=��5�S����1�j>��<��n�}KZ��7(�TߴP�ʠz�\�a�I?j�݀}wʁKc@T��zu%�n�V�;�D�L�������$���`h)3%��T.��vy�t����P����~�'�]���f�mV��/ � S�-���H'=�S���R���q�6��0�)�>�A��<<\~1Q�d�)�4ٍە8��.�5�n�4��|�rp5Y��Щ���_Rˢ�]O�i�[���"����`�<�P	�=�����v�8��2��By��j�V����c�TaJ�2��pZ<��ޚ�9{%�WJ#�:�$��t�'��,�o����Se�,��y�O���ot%�����L��B%�V\�/���X�����S�L
`/|�&���0��ŰI$"ߕ�x�p�o��ROG�B��AA㐾Y^��.=k`��?����)��>����j��Rz���8��sr��m�$��=��#��c{R̙n�>+{.�+Q�v�F�a�Ō��`u�HAޠ��˷�y�1WAv~&��\�Y�
 �x��݇�6�v�,NՁN��{a&�E�5E@�6B0����f��4�}
�k�3^�����=;��K\��kտg�{���ȿ�1��Ɍ_i7��&Q���c-�F�^���ʐ����8�Ͷx�_��c�ܟ��@t���K!��+�i&�b�X�S���=˥�=N�)P����($w��ƌx�������
-�9^���& j�IU���&�a0/L��%�$����S��Ӽ�Xö���B3�ofΕ\f�3,��&��g{8@���>��o�:�*uɊd�:�H�<,/'À��["���}���� �!�����k){��/�"��"T,�s��=�|��~���'�f}!Tf���&��#��Ƚ���I	�c�aY���#x2��ٌ�=�g���B�T�ˢL9�2�w���9M�>A�͟3aZ·�;�����5x_Tk;���n6�m�o��舫��ʀ�|/����$S��
�z�gc����5��,�DJkw	�J�6e����t�=!����Y�"�ΰ/@�_E���t�	"UG!׹s�2?�v����5y_�'>���J�cIXn���y��&�v�x�m#�H�%��<���H2�:pӌnYp��4��Ai�l�Ư\%݂�8�_�l@� �M���1ut<)��x�I��F�;�=*a҉|˷��&!����d'��;�l��K���3�!���Ii��tb�>]�	G�9t�x�@9l��WXT׍x�]GQ% m��ԀMg������g7E]���בj�Z�o�h����e�H�s�l�u�����\N�YE�S�j�OW���g�-/���«��^���?v&g���T`�-�b����	�xzk���b �/4P�.��=iH�PϕN�k�NZ[�e9�*Ը+�k����DJ;��� ]@o�me%�W�x� �uX� ��S�̪c��\
��I���=L
�[��X�=��P�/��sH�pv-|E���p�U��XP�^?�7^YM�k;�����zgXy���4�U��L̌I\`cNNa��k��^�h�.OqUg�I<_� evۈ���憥���ӺW���Ɉ���
��/^�_ʀyz�I�/g����:����9 ]%xqB#�9�pN�[=�h�)��I��.�Շ,X�ý�63����Q���/F�$kDEY8a3JE=����jpA�$A��w-�	�A����4����: e="(�Ж6��iqw�w2*��گ5���z(6��[1S9p��Y�|�GG��0Yŧ���P>�{��[^�"N>*���8,G�L��v��mjN@�������1*�3\��t��{!G��\�m�G�Z�aa��'Ϻ	�yp����f�&a���D�&_&��eۙ���|o�x�O�����y����p��޷;��"?�u�}�f	o�_��VNP����kS~�P7��$2����* ��j��lb&�Wb���Oڨ��d���A�Y�/�ok�q	�!S�*�mPu��B�<���+R� ��7��A�'��I�ʱN�6�U�˚�Jh� \�Q�m`&툜�wC����=��Ũ�}H�X-�q��#i��g��@=Ã�M��d��3��SW&��C�A��n��������h����܏��
i�]�:kR9@�[�%:���a��"���-�Yd�<��s�=��2��&�S�TK5�d�Nmۃ"���:�N]�.6�a��7#���*���nh9{�E�3�s�N��f�K�
�Ы�F��o�_�����B�En��
��np֔{��������K1W�x�( sK7�Bp�~g���Ht�#kB�%���RT��[�!�/�^��C�a��^}���Ap�/���v *w�q�׶��f���SJA֌�}w�;l�F�a�'A,������{�VМ$���o�������G�	��F	�>X�%G��})�`U��7�x�N�*�C*��j�_/�2��0�YOJ�!��y	��6�fޑP�z8��\NE7z4�ڏ�MB-�n{K4oX�����#a������������W�^4����_w��q)z�X�<˙|n]��&���!'�
k&��%��s$�,��2��<�(!0xpK��C��E9tu�j��<D �4�Ơ���g�fT�k��6J?c˚�0�S���ַ��`	�杽��G`vlWxkC�qt*Fͣ����]�Z[5u�!�#�t��f� ���ځc�QQ&�����+z� ˫PW��m�7Q$��l�0���0z�h@+n���+Xd͑(.�Kl�y�,Q=���\�#����`�L鉄��{�:Q�3'GF���e�������ݐO�*��|b�ڸY��iS�����d��q�b��(���yV~�d涆�qe����L�e�7e�r`��F2=��#�|ڷ��锦�����5Eꄯ��`�d�G�,�Ƥ� g���?�L�:\���{���T��­y��_���s�f��%��F�y��N�߄�b�8�7���<��`�ч5�h�����¡��όMd�Ҭ�ty�~��/E�`���Ɖe@���r_��K+n,!�ú�:��Y����Zd��	�z�@�	��>�_�;(�V�إ�6x�Z6��=��^�tW���������i����qcK�43�VX����&�ti��C"���AAi�j;/��K�hAa��o�>���gDQ�k bN`5��7�܆��1S�{�m�=�l��UpYPB�5θ�xCqu2<>���l�'�&����ǲ �}X�gLX ����[����yhoM�4 z�>��a�-I��R�%|���4�P��	�{�����e�	$��uJ���I��Of�׼��z2��$`Vs6��q���j���:1(\�N�N���ԅL SI@j�d0@�حLJT�պ�7��M">���?b������it��������O%�	�M�A���CJu ��u��x��"Έ�A��a}�/�G-MAIv����O#zr�Y�"�u���Hհ{�� �ZdG��`v�Y/P���4�2��Mؽm{	L/no�v�]�������U,3m�B*!6�N�"�Ս��ŋ<�q� �V�2��.�^P�b<rR?�[��9u*�#��~q�u%�0��<�<�G�P�ǵH�����إ�m�ʀ�[���*xܴ4VW�t!�G;���O�dP�;���(�Z*�m����E�(���Ac;�m
<o��RF���M�9����U;��IU,�<�<�rDt���� �Ǩ�����w����HO����_w.��t��oy��3JI
�m�A�g�o�P�k?�0��LF ���ڤ9X�-~�39ĐZ?���ߠliTȪ���q� n��A��翿��[<#=����`ZrEl��=�#2�"�X0��@8����:ʞ�Rr��H�s�Q��FDS3s~��Qs�y�l,7���XFFes����v���M���r�]ӻz���
w$�2���Cd����BWjbmn�� ��(/s�e�Qx҈t4ġ	��ZF'��j3�"�+��6�dߩqX˖���� ��~��l�=���V�wq�H��2�k#]���!�b@�MM���x	��	3����=��K(c=xPJ(�@g��d���~Y�/&�M�>�`�ՠ�Ut���Zb`�vT�����Îb��lxP��z%J6���3�ӕ��|���|`�e%��:����D���*�&�q݄���-V�;�P�֕��)f���V�hL�%k)���`�YZ��fU�C/�o�]Nз�v:�/�y8�m���i��Yl䏗�ؐr� >���C ��������_F+�Y������#��Dy�>+�;@��E!2l9Vu���,;�-ņ����-c��F$a� F��Y�J0�V��gb�qp[�Xot�}��ґ���ϧz�\�Q �tw2I�J ��.���fo�`*���t��݇�-��z�!ڈ.Ų�VM����)�թJ�;��%�$�=�矖�g��羖�s���j=BĂ�U�&�n��H�F�@���Y����\xf�c@��rA/	�Ŭ�L4�Q�q�*v3���h��(��������,��v����� �VRhk��M���8�B������2�Q*+������ӯ�T�|W�05��FN��z����U�&;��xo%[��s�#[�!3k��,��а]���+��+�n���;^�	C��g�(dI3�ڟ�a5��$��r��']��)g�Xk�dA}ډ-V�P�Ql�~bP���-X��3A˖�D9���v0�z?PX��b*c�9�ɟ�9�%��H�����R[����}�k+�c�ԕ	ȯ���C]� ㆖�ï��R,<z6������5�e���6�-5���~*�P7�<���>��e�h�X�$6>���9td��mUGe�.��'T�Ö@h�֩
�o�W��Q�����O�+���0.d"�t�fm]εV��誇^d�p3�K��V����3���?7��+���U���X�j<���f��p���+o� 1V{`h��2�pX�w���L��%EX�j��(c�g����a,'�XIuӰ	_	7�m��%�_�Q�ո�_�L�ߋ�/矃�񥁄�e���A�yl��8��y4�9����Z����-���ݾ�z~,B���
��ż����"���`�c�-0�ղtNѤ�R|:��U@�)�o�������G�Pi� .�5��U��}Lեz��2Y��]$�r�����
qh�H$Z3��q��`��q5�u���G�}���-�Jk'F����a��P���n�t�~n2KX-�c�_�z�'v<�M��s�-���{t��,������$�p��{��`�H�&�2�yn������+�ԫ�p�?+�d�;�'��
��_����d*6�t�8x{���^c��?Nt*(V�t;a�2��\����H�Xh��h�Ƞ���;^������'�3Z��l���LDhܨ�x%����1�Gs�f�-˄'�ɐ�#��m2�����[�����	�� 
6������~ңs_ڶ<�u�z���ނ*򭱧�raj<��JY0�"`������ ��~vj8v��O�/�m[�H[c��R*�6˵Yv��a �l2�3��L3=��%�o�.��DZ3���J��-eN����ַB)ʛ�S&�vͬ���X±}�C�(I�1f۷����JN��3@���z�+����b!n����Ot��3Q�����r�Xd�<�a�E-A-�ԛr�Ou��A8��L+����X�������k�C���b
���H��K�6�i)���ҁ��eī��n����e���G��x&P��w��4s��j�2��!⚩S��z@Ҫѓ4p��tT��M��RƼ18��<��pv��K��u���5� 0_���lN�l�9.�0nδd%�n`��f��J|��h*����r�A�%G����n��v�xj�ʱֽ�"�`/�6�:�|�bc?ȸ_	��߆�������vps!S��p�Z�O�F���"8Mo4�K��/+MQ�����@;ܔ6[(�RT�\���ю9B@ �"��f�Ӆ*�Ur;"<f�U)�vQ�K������N�a*�,���+f��uP8.9aBԴ8�7^{��Ո��9�tOT�[�mղ>lm*�NEB����<��rzK=qL7�rLJ���o=��W߲�ޒ��	X�}��@�Q�Ը�l�X2����[oy������
t4����uMw�0תp����+��%5Z{]'Jvx��2r}�DS��~��h����L����ak�g�4�����-s����0vV�H�;��|�d��HL�)|�u��Lq�0���s6s�8�&�Ern���[�+�>�?Ӊ)ؒ���ƻ�u3���{�������� �RW���dŶ:��ַ1'o7�?(R�mVx�CX��t�{ӈ͵�C%������o��D�7��0�Z�17���{�m�C�٥W��s����ry)Vz�	��`s�"���p�i����LY1���{���l���I�&Xo��[��.��ƹB%�,8[�L53⺵^�Q�Q��ɛ_��xTbF��$�+C�\{s8��~�=CU}O�^X�Gفf��ƣ�7]r�����Q+Hp=����O5�VG9\b��q.�z�~b�{x���9{�'7\8W����%�� 	��R���W3z������Y�ЭP�!m�O�9z�x��KSA�cD��#L��v��1���ڼ�z��K���x�t�s֤|F��G)��o�P)�>=�&V"K�k��w@��M܋�g<E}*���0��Р5�Mޥ�A^O�Uuo���2������w]�#9�+q�tz2¸��X�-e>�ϼC�6��n�]�;�n�tL�ǝ1E��p��()$���+�r&�����ak����t������tnB�d"���ѹ��;�����T)�غ�Q�j~{�$��0���Nb�@�Qk|�=
{Hb���a���>`&:`��Ұ�2���W�׹t��K��lͫ<̜�����;�����i�cE��jI٨�ūX/���?��Q�V���na�?��cL��Aҡ��-�9����#QEL���5C��>�A��Q|�PͦB}�}�{d��wRU~���ᆁ�F�Z�~�˫I�JJ4d7��g��Gܹ��Y�L�Dp}�+�@9��uz��>M_��Qi��`!~vŁ�0�C�d�1G��`�(��������v�����ύˌ=�d�Tt���fW� ���C���l����ʺ���B�TUA��	s�����/2H�]- Նl�Gʁ�U�	���m����W*�Og�����O��!��Ers����*m��P�*�=��G�{�ߒ�4&�C�Ç��&�;z�<mj���q)/~�CRHavlO�AxxQ�����+�ǁ�}�.D��RkCQtK�C�Qh��	�k¨fN.���Y���!��1�0Z<-�2��Y#[e%,o�˽�gdM]��)�9]�	��E�&�JQ�*|�8�� �L�v�6�5��}����"J�wN�_Y�cW��>�/�3�QS��GO
 �8;���hl��ѱ��&��U��Rˈ��W��3��T��z�~������#?�ҩ�+�6���q�,m��{���J�s>�
i�����T���U�c�1h$)�o0J����m�����z�W�N���g3�X���S]��/	��7���Í���'����P�".9��\`b���W���L�U��Cw������i���.�8H�U���>�R�㍦�I2���S��$A��"�J!ݵ�2rj�;��Hz�9�,fx��e1B%f�z���Z�^l@|���#ew�gR�(�sD�q;(��H���Ny��^��LH�>QG���Z�_4��HE�������}��Xb�@0��@�`e���0D�����n��L��	3�{bJ�%vit�#�6,�?��f[xxTy(�[pP���?�`V<��9P�����N#E�wo�֕�ZO��6!_�#�E���~]*�IV�헠�ߨ����Q終.Y���s��HW``��Պ�|��p�U�R2�g��l�r�0��iU�jCL?��@�$F��F�AS8˭q>��4{�f
<�6��H�f킭=�D�'���U��=��b,����+��H���u�����L��aڥ�������{%i(xAuK�Z^�L_:����
H�b�G�v���SB���Z�O��H��|�>y�?�� ��jR�#�)����J�O_=#z2-.� �*ۥ����P���M��Ǥ�f����L�Pl���SǼ̏��R�#�W~<;?7%���q5)^ɪQJ�Z$�����ˆ-�R< *<�~�rA#S�H�[��@����U�*��UQ�x_�evI��_��5QY_�zb���xąSo5+J-f��FJ��J��d߅�k���0C���"�T��X�3��+qP�h�Y�V&`�i�����j° d]��-�|�)_P)}(���Zqk�������#��0|��!Jw�ݐsj�Vy�f��I�]h>��*)�����ۻ�"Re����}�nĿ�n�����3�6����~�f�#����F�R)kry�ų!�s	;Z�7��/�j��=�L%��v!m�[�9]7�c�K��66��T��\�����}O���n�4���d�h��a�Jkb`��6a�
|4{�wh�F���n�aIxW`�����SBCA��t|�b;���-:Q�5���6*�7����c$�F�"�)�qn%�����R@=3$ԭ���i�t޶�·e4gd��+:$�4�P���1���8p:���ވx/�͜��L04�?p�ؕ3A�~����E�VsU���RA���'=j�8���a�\�o��A�M���Rc�w��#��P�KcwT�{����aH�ΒΠ�̊�cWV��ۤa&�'��V�d����s�~��OS�_�2}o�
R	�p-�k4�_/��έ�\P"�Z}�^h&�=Is�@��r��>X|7���陬�}��U;��`u�W���,Cm�T-�Z�U}Uo��?�p��&=�d?ӡ�jr�?R�&��P1�$b�v�7�����=pDN���;��^��e���m÷����Jz�TC�z��.Y�����4�9<
D�����M�>����#|H�k1#���蠸lĢO���9�U��)���LV�6�S�P"�hL�5��A���%��6qKEG�C����z	5���mafO�5d���2���
S^�~�H�M����E�<�@B���W�f��ȣo�x?'�f �T��<��B�K�C�X^#.�,h
l��e�?Y�:|�w����Ǉ�R�.��0���;\�1��Q(c�>��,�T k�����d)�@��s[��Y�]�p3�sd��壙�m�����xzW��oΚn�F4����a~�է�-�����ts�˙�vG�!qC��kBQ����B���P��&D&���?��Q�?����V@j0>��X4�ّZ5)�]�[�x,.j/5���/��+ʼAG�z!7U����m��c,Z��;��ݍo���K����C�������Pο�pTܯ�n�/U����m���<C*E�=��(�Bq#�y�$F �w����5�y��?��O��K�B�t�PO=6|*�-.��n��(��+JG�e�q AV��r�� iF�U3%#w
=7�lZ��z9���A���u�F1,������t�p�QVk�˸hZ�̷�۰�� j3�r���BDy�ou>��ġ)Z,����m+T�M�>1V��� �m�J:�+B��{P���p���E��I7�-k8)�ƾ���2�?��S�wG~������2kt
��_���2}p.0��qz�?*��F�KU��{.�m]��S�X��w�<����`}L�*����lP����$�cV�I��.��,�n��&�a���@k���V4�F���b�%XwWsu
и�� Ѝ�ӋS�d��������ƢC�Q���6duoP��t�>w���D�
�R��嗄�;?�omU��V�/�	BS�ݭ��~�m�򼭘��v~�m>o��S _��-�I�4,�p��UQ� ���ǿlXZ�"l��]�z��E1���M�����
2a?ߡw��?�rT]#���W̥lu'���x���$���pg�&�]$Ҙ>)�� ��e7nd���F3_x��6�>7��m�{i�������C���O�Xx�/n$bw�F�<)N� ��S�~��L�)��6GB<�/|._��O ��q�|���xz5��6|�_qlû���"p���A��4MkG��N�\qt��(��x��z�??~ٶ�����qj`"�Z<�I(��o�en^j]D>,���JB\��1���e��
."ٴCv�5s��y�:;�,��%h�z5��]A*����& �j1�����w.,͍�6�B�3�����~D�M�U���I��8�#Ru`��'Eµg6M�����}�j�X��H�ۈ/	+f��-�R���v$�l@BO�횬ʜH�cu�t�}d��d�Q�ѹ�Y�ز=nC�������QM=p,��(��#���� �K��X��E�����9^�Zq�$��hZ{�}��-U���~o<����/gr�^�p��{�	��2�b�u܏�[��&X_�0a-F�<�ٖ�Ao�iУ�N�Ez��P��H6l�Y~�a��J`J*��%mIt��%v
��^~:A*����4�3=��s�}y
���L��VVn.$�O`l�9�5�5� N���鿡D8q�a���x�}q������k��&�`���I}cDCMIӮz/=�l}祈@I��&���)7�?G�d� �¤%��ڕ[٩^���.5UD;P����v�d����N����̢%���)��y��p5k��?c��u�y0U�8�N弴n���1f���H3�������y�8�2��s�A*��H�˵�4�0�)�ٮ�+��Zˍ���_�&\�	1�qѥ�_ .�G9����uJ&P�d�h��]ֽ�$(���zZ=��jd�}�O��p�l=;���r^fV���+MB�V�C�`;���i$;#ғ��KWk<�TΪ��Gz�~,�MwH+V����?�6�6��ԫ�!�| ��զ��l��^�Q��}nQ$�.��@��C��*�k�����e6{mt1��\��k�����fH[)��^ʾ��D�އ��uz�eHs����j
��'����[��~I��	/�h�~�/ն�!hqYr���ȓ�օ�ɴ�ps2nz����ʁN�3�'��/��=���:"a��z9��:���$]R���`�D�YL*��d ^�YdA;������xi,��xu���!Ӯ�]*T����qm̓��봯�Rh��C9戀$�� �~�� *�����횞=h�V��#R.}��H�n������S3c�|�Ī�EO◸���E��� �d�2���K��;�V	�^�_p	{r��z��@"y[VV���t�:���8�����U+���zq1ж�����R`�>�D���长WD�/Q��꟏��ȷUt�m(;��f�fo�>�S�Q���t1Q�U'df�||� ,��D:�l$ᓿQ���_�� @)4f��m ��7�ĵ-�M�p��Yu��H���ĂrYl��d���p�S,@w^����'��*��l����'r�$��M���� gѥaK�I2���*��UJ(^�[nԹ�+�olY����w)�C&�����4���vE�A4LY�����"N�功ah>�s��>֭�{��FԌ�+��A��r��yr��f�ҭ��"��o�~����:�-�a�dc��-cf0o|n��2��d1�h#����6���vP��(���W�CvqO'&�~φ��yp�p*ͅa���}���7���Z�J̅Yp1w�-�*G%�9n��铄Y"s�[�U���Y��siZ�)dv��g�S]��/`�u���t@!ý[�7�����AnF
�5R�/~��r��<�\����P�+��7CZK�G���'�o/X�!��N!��XQQdB:������`S�Y�Ӑ�7�:ϯK�t�ԯ�c�`�a��H�\�
���,��������`�|����p�z�{Q<t��8K����z�:�U˝�=��Z�_���0T�a�I�t}����$%��g���ܿ^(3��ؼ����I�38J�՛�T�~3�O��r.6{J�:z��(3�A�m��nU�V^#�G�z�}=<��V}���^����Cc��G����U��2�$����E�]��fh��BET���Ea�Xx�?�g�`Bt�,�¯���x�ShW���e��֘m�ݰ�Uf��Qv�Y����e��6Fղs�#�Z%�Z���(�!�@���>���R�Y0z�e�C��^��}��a:V��~���@��<(�^c��.F��ý�x�2��8�~H��y�MWw�%�Lsvc��Y$�{6�'�n�m���|G����7�U���piǋ'�MtZF�1�j�Y-#��ě�Z:ϓeZ���};%��'n�Lq$�R�z��[� jt:�:AͿQ�a���
CxYrw����E���v 0�U�ݺ�>C�����4`"ٹ�\�'s��D��EF)4�\�L
�U��2n�@���XD�
B���W6D���ԡ[,eQ�����j��	�n�<rW�����0�cM��(o݈�m�ua����mЛ�7[�Z�E��-�QOk�9��%v��?5�%�~-�oO�GY�X�j�F�'7�j;�r��y�a5�\[���SwF�$6Fy��������]�Nu8tM]6ڷv5���{��d��%�s.#�F��Qo0�u�§�o�3]�Dn��c=�i$~��J�N��z�r��i���.�\:�����қ;�����0�u^��I\�3� I$_�?d�Ϗ`>�,���H4�3�g�״�^�T׭��Q�|H+�;^��bo���-���+�S�p[q��fPK��=q�#|'Y�:������%B����_-�"��IgYƫ*��Z�~b<�O����	d$5��S�Ci�~{���c9ll?#�=��ԧ~�8��#�m���E
�2�-�Ƹ斻Җ��K}-����I`(׊u	���dZ�1��@�$�XA+٤fW}�<�)��m��%s��Ŋ(�`B�=�k��RU	>����Eh�]������8��Z]�5�[�����@���qN��o���Z�e'�tL7t`		5=e-�ko�:�\`�y��S�X̾�^hvv�(���i�}�,"�;cgt��v�����7Gl���im�e�i�k:�B�5�pz����3M���C�y��)|te�^�j���*�:,��`��B>�;h0�	*��;U*3����}�w��ĺ�#�
C�^Lʴ���E�(�E��]�x�� ��,^��+�6��z�'z �(��GE؀�����׹�q��~f@���i~�ry��g���	�B�ʡ���1.`������j��H�(�4_�J;�3c�\q�nG��@+�y�f<��aiC\evM�E`}[	��b,�t�83�\`�%϶̠��4F����Ҟ����?:9��ѭ�OD{IH9�%sr>S�)���
�GS��ʗ��Tr@<�4Eru���sL�})�:\h�L҈�����8i�3AZ%���r5�%���9b�'�_�:���L�qۻǠlKϸ�ک����)�;\�g�
3�2(����1J?er�0e�߆�Q�#:U�h@�ɜ=�\�>�����L�|NR \������7^����m�^p-��	���w3TE���#�SJ�|D� 0|�j��n��@	@�S�}�s���t�A:Cu�H�c�苑R��G�q��q�k�yy�f�Л��x�XU?K1��:<7yM#el>�D�Ju�X�Ws!^�%�`񃏨(Τ�h��X��Ov�>�,l!�1�+àJ��O*�B��aBw�o�i�*�{����8d՝����zT��A �����S����y'Zm;��KiL�VK�9�?X�x�]�^�,��A/en[���k�΁ڋ-�5�3]�f�
P���b8D���,/��e�VC&���U��7��t�,�m�ڪGl��E��Nf�+G}�N���?	�5�еd�^˖�N�����2O�I�۸k��?����\O��;Ŋ�-��r%	-��.c���/ˎ��S@�>�(��}�w���y@�l�Q��C��$v��|�ZT6i:[�fS��T�r��AX+��`��k�%��3]gg,�n��*�/b��}�do��	kБ2��8��E���G4[���)�~�M�b�I�4�z �L�n�Ъ���o�?�~�el֕i�����:�܎/R��V�9$Ny���S�R�3�� C��+�M�OY��?,5߲'u7%��C5�����t$F]*e�#@��Pj��P�(K����������4��ӹ�����$�ʈ��U�sy��ȡ�C�X5MQv̗g	���S��mJʇ�"e���
|�����C�`<x>_>�n7�w��DK���6Z��qV487P�aFT��,�Ƙ"m9��U�6�_U��O^�L2���J&��ٴ9�F�Pt�)_�	a��P�/�)���dIL2��������j��+]�i�K���+��o��l��VV�������缡���O:gz0�fhl[H���킧2�V��~�����-v����$I֗X�s�Z���(2__�H��k����m߳2�B흈�����P%���c���Y��,�~�no�L����X�I_����v9f�9�6��v�d,��J��5XY6๟Rk|��_�;�\ާ����%�?��<�-+3��S3;�>jO8�x�E3���D0lm�r�=[U+��~,(�nz����{��x���e��LJ��T�v��+�_�"�C���Y��QJ�
�7�y��=�_6��Q��γ�;飥�4�lQ������
�����b���4����&�1*@)1�l��?�p{�o gy7�>;�`�ۃ�ti�`.�,ȃ��A[��H�N9�t�[%�hm����F�P}ZPNǅW��{|�e�6|�T��/�7E�]�S��e4�,})s��[��p6����_�����M�5��#�7�4E�Gc����ڀ�q{J��lGɒX�o#�ݣuB���v B\��]��RnL�Ś�?�f<B"�bA��Ǆ��A���*;���j:��F�L�H7���:�&՟��Z�X����ƕ��3���)-/��zX�،�}3B�
�ʬ����׽:��0��d藨��σ�r��oļ��A�hq}	ÿ��ya����| ���U��� tj��}\#Q�:�#������Ѭ��f����aZy$�mF�e&���D�Hx��k��= g��KKo��k6��eY�M�'�\��y&�X�x�⁘����g|�u1V����:z[��ުC�: 4�?��T�sQ{,b S����>[ܲP�[ey���1�|ڽÖ�M�f{�3ZF{�Tݝ1�z���V�Y�^�ha$R[J��)6*9�bR��ނ~iJ�J5��z>�-�V���*�s��U��v��0e�@/{��+��[�$2W��$������Li!_t��o�S�^Kʦ0%j%z��58"fr�rO��$^'������	��#���i�P�Z�{�Fp�|��[�T6d�L�l_�G��/}�'�����W�F���<��!3��^N��>��i�{c=�~�:�U[ESQ���x���h�2$�$n?�"��t��u!b�\_����2�����^��yH��e��|J�WWi��K�FX��,i��&@�?GZ���#�>�/+7LY�;6s����D�Pj��*�6�;���@�/��D��}�	��(�\������Nk��P?�Zؘ��Y1a�a��F��40M�}eO�Q)(v����,�ůW������X`��N�u��5�b$����$f��������h�'@e� �t<e�x�=m�Q/U1c�T��+��^J����;~�M���A�0�/Z($Vl��ւ�7]������І��?{��9�"?���+§PY�V�����r��lT����3�!_���g�L���E
~z�b�x���z���{|�ߐ�";�B�f��쇹�T���3�f��\j������/�//�P�a@�+�}�0X������}B�k�"X��<��
���^Y�S�t�V�Yw��FNA�������2�U����*�Ч�1[��|��Ҋ��|;,��<���u1!'RKk��;ݙ�1?k�<�mk��	ӱ����֗�y)�ˤ�G��6�B?�����	_P.��
�:�x�����q��0e�5:3�O<��W��$�[��v�o<��)��0�V��(?���`�g�&)�?w�x�H�(�3�]��p�ʠY�<��'h�x�co�����-��Dz
_�[�Y�1	ھ�0)���1�@ܸ���������ir�[��J�	�G
�v�!�����M/���&3LG�8�ZTJ�����䏾�=��Z�Җ����]ɜS�#r/�/x�3����G���z���,F�Ŷ	ή�m���h�Ƹ#nSڶjB�T
6��\�Ȯ]�^���&M\w��� >;}E�W�>-�(Ҕg��wÚ�]���Փ�Q�l�sn:K���)yj�)��np��k�o>������r=;�譼巑��2�'v�ɂ9�V���~@����X2Ue���v��B6)d����0^����Q���~���G�V���%I���e1���r��,��i�e���UMP�ۊ�����
��=�R�#�ßy�j���$O&
֧������}~np���&#�����0�� �Z�z4���;�8��57D\J���,�<�FW�� �)κ'����+gE��Y��}ϒ�{��D&��BL�R���}��������:ۄ�ۙ#(��Rt=�Q��H��I���OH�&I���	T<o�ֆȇ�@5ܡX�����������ጚ��jw7���z�q�{<��� ����^kQAMI#���, -␠���}V�5��o��E/��5�B�f��@30N��z����An��VyY��9�[>\���WI^QdNs�N��
�"���X��x�[�l�S-�b�b��~Q�S?@��&|�j	�?���������$Ė"��/���́�`d$�e����#N�����7�������֊ʕ��L�	��?���H��lzj��S-��bӒ(��]����¶�,�Oܠ��7+��t�᭫,T]�\6�7� ݌^��^�^I���-X"n{t�w��2�P�I���{"����Č+<�T�Ա��JΟ�qr���*D���� ]�;uJ��(����|��Mw�����M�<H~V6=����3S畍(b:3\z�X��<�Ͷ
��	Ho>e���T���$�H����	(c�
�m!Sf��{�]�O�h`a���M�J�ڂ��X��4d�X<�K����d�h3t�:��Q�#U�Ȏ�%V�5�l���yr1l��4�fb��}iSr{�&1N\����>n������B���M�멖��li�N��?x��B�lz�gv����4{S`R<�	�P;N�v77�|��*��wn�dGC,~�>&4;�T� �����u�&�.'|y>�y��$�G��O�;�`�N#}���Y8�ek\���R�y����������L��a�$�1�P�|��"�m�1+HR��=�ߞ�BvT�����U�C_�V �����I��ʺ��(`Vz�:��\�����/Ѳ�Դ���6��هz�HQ�aP�! �D;M��-Js[C��ʌ�n1U��,��t�bk��
:�aӳ,^�x��F
��ά_qg^҇NpBKA�M�)�J�z�m���;�)�qΊ��#/�S���u�������@bZ�\�8��&+��x/:շ_�5�cYu����EƱ�B���R����O{n6E����!�(b����`@��'A��ʿ�/l��	 ��Ū���,����MӂTP��դ��_���-$�|m�Gd�Z(�[�a�[ \I���C��ɟlg�\^x�i,�Ė�`!��J��������dڳ�O4��r��#"�����qy~��ټ�9����f��a�D(����AW~:��s��1b�t�iX�g��
ۥ��5���jw��6_0[.��<���G��/����>�n�3nu��b��ś��'�V;(���}��{IE^��(��S��Z������gx-�"a���pV�<s�C���]�NkC4���Q��B�����,<��vf�[a3I�h��sx�~�b�@Xg�^���� ���<����+*�4ݫ<��?IEp&K���}�w�(��f�i _����u��"�@_lhZ�}�(���X7���)��hm�^��6���&7,�g���
���U�a��r]!v��%�EIK��cW�x��"hz�ɑ��Zo�G�;i�χ�	���y�KV�9_��9����(���;��p�
���"x����k������$cL{R��?/E�w �M�:^"d�N������	r$&�1E;�������d��8����B��_�FMԻ����wЫjc#�s�_�G&~҇��u�8��62w��p(��b�[�3L����dmn0��^���|}i��H*"+��y폃*�6��'����F{\Z���قV����WıN�����C�,	�l�s>*_����g�1<�o��9z��v즻~�*h_~?x���GS�&�b��>�g^s6��A^:
j�=�	=;�^�"Iw���!cq�H�3��8;���B�>Ǳ��Sc��8�?��y���z�9���W~��Q���T�#-_��搼�[��}ѕ�1t����4E�Ӎ��b��9�Uq��cq����L�pܢ�k��r�z�O P��'�˝�i�?T^cZ�eʿc����1g~�v՝���?�$x4jL&ڒA�I�c��"�}pf�4�e�=F|$z����θ�ik�Ǣ�|Qw��f�1�.E���(��|S볲���䃋Fuc�z��2��,E䜡!�����0��C������K()ԕ��YY���1�9cءoL��EI�x[k�u�c����P.���a^A`��C<�C���'��ߌ=m�U.O�b�FS�4��=�Yk���n�ae�t�v;lta�a	�ґ�D�~�XG������uX�8V��x���#~ZH�9�85����
�k��-����8��ྫ´i5i�������V�\�����D��׫@��Y(=����8QTi��<��3a����6i�)���9��5�t،��}����M���%U�qι���P����yw��QQt�K$(����h���U�}�ZZ��&'���-�9�7E�Y)�p����.J�9���Z����.z�D��h����j��llt*J�Je
��] O��B!�O�!L]�#FJ�N��鿺�J���o��_�f��b�����(S��8�����3���+����ySy"9ܛ�bM}�@�j���p����n��VYa"��w���ϵ��
�\V�uQ%�ol#���(m�8]Zs���̴����Q���o����`�Oة��;�u:hLN��us��!����A���Sq�Oc��n˛r��s@]�$��/�9�O�Y 3��
d0�����s�,����H�2�����Łs�Uhƪcv�v#�Bl�L[�dX6
n6�)�T�f�����&H���C�s�����7�^��s[.U��Tw��Ds'9��������b�>_@�**��9��-�95�΃����g���h�C<_����a���I���d
l�<L��1%�SL+;�& 
=&L��D�*���5��R�J��"f݊�'J��ϖ� �d(��,5j�h'�E�E!ӂ�N�+�*`���l��ό2 ���,��=�/(�v�y�GY�vqἮN�������=۶w�H��4	�;!{��Dq����Iă+k!��:�#���a ����=
�he6r��EZ�p��
������L0+�T����ePn;"���ߞ�G(r�H��?�� [�5������V�zP4e������s<���[2��y�cU�f���܍|�z6�~HE\�~D�m�s����*�����d���.��qz��y�=0=p�Q�j�h�5T	p�M�])�:4��ӻ����r��ǽ��	&v�!#���Wt��eDk�WAit3`�l|�C���53��A��S��C��R��~b�S�b�����n�3�)�I�����-��a>��a�S���P�φ����d��i��R����d���V>���|?-`�LЩ"�W��]
�C#'������ޒV���Uwy�a��X�v���ˊQ��M\$e�~�0}#�O|��*Bd����Ha��+�Io)C$?N�����CKH�"��4+@�l����_?Q
Wa�b�*L��E� T�
�/���cSk�Ia���HT-c7(�����M�"o�nN���y/�&��_4S����j�Փq�ந��x�̀�/g)�.��U��'���S��(RQ�u��y�9(^Z\h�����R�_+D�I;J���� ڰn���D���s�Nvд�C��{G�"8��\�{}Π�Kr��W��/����*M~5��gӜPh&|-�/�^j�)q���w	���1��_sF�2��A�|?L<HT�"��y-$��,��-��-�
@�X��/�@�l��̿g�ڝ�(6�}�g��.X�b�x��_�6t�Y��:�����=�qb�P����Y�S�h۾;�K��:_��Q6C�l R<��aK���B@��9�m��u��hnS���-� i	�ְ�wD�o�؋d�U���n ʏ]ǜ'δZIQ`Jt��7M>ı
d�5t� B��a�׻ט=QM,�h�l���5�r�|���?�vҊ��&	�9����3�4Q�G)c��趉���n�UҠ�R8*t���˾^�x3��h��#��7�haSJL1�>Jn|/����F*�+R��Z��*����K���
��(:'
3@�fB�$��v��Y�ɣ}߹���K��p7�޴�U��maMy�bw�:2�']��U��̜b)��B3��㫸�O����˹��W%�s氷�P�C'F�ܗ ������G2�����0�*~�u��[Zy?�g�����K��ֳ�-�(�y���J	5�?�})eF��v��h%'�7bs��|	�i���֕;/���@�����:�D��=T8S�]��|%�
f\$Y�Dn ԛ��[��|A�6�X�����4	�ps5��X��)A7�\�9���ZES`y�LU����iP7)˦#��* �E^m>j�m�s�3�k���=���̀����|��P]'&�N�vEd�N�s�3��O9PG�8�����a<��o~ܨ4�ր�`�&x,�Rĸ�u30(�,C�
w���e)��ٛ��:��w���7}��#��kňg*���5QB���Aƿ3{�}EGI���~��	i����(�r�����].gP��|3� ������7��"�T[ER%��ˆ������8�K��mJ}�z�+�j���{�,��������M��Ï�'��qz�f���yE����_π8p�I8~T!_7PJ�V*��Z����\��qޟ�)U��8��nQXH
����>�7��-��f�hA�����*��ɚiYuA��.�w>���bBU�����Cx����=��|9�O
auG�ƻ���ےl���*��}������H8��;��j�T���	�Jr���$-��?��0�.@�F#|2��K�+�A�bM��N]S�"R�$�`~Y�tY$��7	����&��]6��{��O$�3�����8&���5��\c�q�j����P��i9��Q��$�`3D�y�XD�g������!���AN�/h��8L����Q��g�����g��U��[��L1�J��`��Xߊ�TA�` h��e�����s����Y�}�v��9}H�ލ�$%r>i�+4�%R��+�L�Q����I8�K��[}2���E-w�ו�dv]����$D�?�� H�6����G{.$4ol�g��U�-�i����l��� @x#Y�� I��ƾY�zf�߅X�ui~�{7��g��5>�����u,uN� ��&���]�Z�����h ��^9���O�"���zF^F��7W�ǻ����`Z���=
��ㅌ�4#�'S0T�;��$��2�\emB���q-�y� }X��D�ca���UΡ�1z��*�-�<�Du��l\#�ΚIs���t�n{�I�s���5�a�*!����~��y'�JY��lm*M��ZѬfJ�~ �H��
dV�U5�ջt�S��'dh��ŕ]f_Ĉ�s�>�ԙb�̸�>�T�bB�_�)�T1)��ܾ6i�H8���T0�v�$x�\�"$�.��2����𹋇�/٘YZB5���h�b�u.�~^����ث��{1�u}��  �\C�6�ֺ��í$ �<糖��(�9�lr�7��D3��+�����K�:��k��#{S�s^?�c�².)�*���P���m�q]��v}���&Y]c�B�=H�e���5���!&����1���,��N�蔩�^�r�c&P3��%�'PC�V���Li��������g4/K?��D����\�1�m�k�h)<Fʫi��\�3�c\���@�O�l���kb����aanG�50W�0�0�����sט�Q9��$J��S���u���z4d�yi6��$NX)���\im�2(�?�����s�d��/h*9uy:���4�>�t.�6TS�-�kd{��*���)�-�%�dgib�rg�s���	�d��<���^&�A�H��2@3c��T�5�����t�U�h��;)�C}�@�!0�~`�xN��v6�		�("�U)�$����6_ްƺ����AY�L�K;�k�S�z}B��ˑ,�J.�jKj-��p̄�4ݕ�08�1�Z�!/�Gԫ&(ۊ%slqy���y��{��m^L6�����V�����m�<VƬ=��d���u
.A�fm�J�}�+��1�B��Le$�P�LQ��>ڐb�Cxl�ª��I=��	�,R�М@��z��Y�ji����}	G��%]��2�/�m����}�x��ad����_޿���QN�)~�j
4����xEv�q�y��)p�$��U���
�]{��4���!m��'��s�Y��s�r�O<.��9��}��$�m{�2x����>~hS�ۭ�L�N6��V=�_H��D��q.���] ���y�jɠ��3< �ƹ����Y�Hq�ў?���+���,�����mɫ�~���U-���!t���.�B	~K��+�	�xc����!�oz
d_J��n#�}��#&ӛ=�v5���4V�끢ڔ�z���S:��р�n�7�pP�]��*�	;�ġ{g$�����b�`���.iq�����B��[,��0�TKr��)�-/������� όC����܄�l)��K�Ũ�uLS&���D>��dU2�����;N�C40+FaH���F��m-��g��o)��ٚ�m�ob, ���Rj�@�A���!'8m?�L(q��G�l���0��Ὁ��\���E�7��\�����$�������B�W�'&Is�0[������=W�m)��ae�%���/P�l��a�*�i�z!S��n��{9�[I2.&Va����~�/Q��I������%����e%��?%0 �N���%�8��,�L�:z_mO���[J��A��)�����C��PU]�Z���K����,e�z08A�-�e�6�&r	��Bb�j���6��� &��������ZUl�h�<0EV��ܪ'U��B�y�Br�pB�;f���4S�D�_��zP&�o>)&V��-q�s��>��Rg���Z�*w`���E �����#�hCƭ��P~�*��1��'�3H
=��M��x���������JS���Y#���?��o�����ըK�7�E#�� ��kJ�<H%I��dbN��;��^>�	��:F��HO�9eA�)E=g��Vɏs�q��/��%�ӈ�EJ�����BG��	@��yu�_^.�Q6���;|����H8�`YP)�M_,"���a]_;w�`��2)b�,y�m� �ͭ�t���.�����\��Ҩ�Q8��[@����7�ȏA�'n�Z�a���aE�@���6��sW$;�55��ur�߫�2�S+�/�߷��3��N�)lpFFn�l�^����3��9��PDX�¬$�Lx5AD���Ā��?���Ԉ���є�����&iRƧ��ӆi�'�i4�I�C�c�R�5��Z���8��*���^
��EV�Q�z�>ܥ�g�/O�I��\�u��e/m�!p�DP$��w>~Mڪ۬/PW��Q)�E�������6��e�C��^��X�i�ߓ�j�,u���E�l�)�v��wrŗ]��妖�4�s͒ryI�a�����f��h+{�.�\�(������'V섒�
�2����z�t�c����C�/8&�MUQ�Z��^�W!KvYj� D���-F�D��0���F*"	D����ii���1?�:��BA�%�ݘ����9y�+>�GI]����!7��r�%t�̳Tv�|��ۓ�>ֿ��]c����m]��7���<tǋt�{{	h�n��Ek�����l~�"�ZB��K�)�u���z2*5՗~�P-���V7R-��<���[1Ф��TҭM�u!g���͐���Q[i�����*ƅ�Vd�>a�F��/�=�r:��m�K�|l��M�t�9��g��ȑ_g��I�Z�g�T��OsE���*59�&��q4����ոV��R��/�>L�8�@	��J*����
}����z�BJZhA�2��Γذj��t��/�7#�+���U��r��CeF�����wͮ�� |��>�Z2~��GĿ7�֙U�6���fM�RF1�����?� �+%m�|�d�+�X|]�����ӖC��?�7��S�%����OI�z�C�7D�N���e�KI���43���1�<����%D^V9�'�=�a0�c��2���bäm���D�K钕�inV�4�4a�K.��0�Y^��#�x�����Z���v�'��d|��h���z��!�8�q�Z��&x���ӿ��Z�KKt�����TؽL������4G��4��Μ�`�,�0/���U:�9�%q�R��Ύ�h�L�+�Bh�w�����A�T����ߺغ���U���G�Eh�,,��F�N�8�,��8!�g��gcz���#�8�M�m��q#�>B��ܠ}��Cy���8JmA��rs� v�\1�%�5�qO0ֳ���@�'|,�$�dK�\� l̨'���U`�M:�H��C9�:�S2ำm�t�1f���$`v�:dtqޕ?�(=�"��;ޑ������8��v�98�=�,|���Vevͪ������e�2AP9�Ϙ"y�w/���*4�L����[����Q.o�+�_B�� 'yд�L�#�����{kЭ8a~4�mC |��~�*�~��R��8#wQ�H��V��8�*#$�?͘��\z)4<�Ca�f�C�RZ�Ӕa�K}Es�%��u��~peЁ�&~�*��7��!�@�,�p$:5+�`_�G`W��R������tE�2lLR�>U0M�l�|�K@���y��8:T�a*�:�暵�ɘ�E�8"eZ:��?QcB��!ҥ�ؔ�B��w��G�,Y�?q��T	K�'Qʹ�{x�u$X[kyA���֤;������z_� �.��`	�l�����L,��$��d jr:p�ϭf�{�q�>�H5���<��f��۟\� ��7S�C�O�����P�0�-�H����qT������q~!��~���5�n���q��E���qI��0,�rb{������Ru*�D/���Fg��JTs������:a��:*���7��v!����C�t�$�ԡƃ��k��L����f���%�t�A
��`�H���;�O\�4��c��9e�:�����N^�w�#
"J��L�gq	:h&S��%8�ˇ1o8)s1�v�N�r����Oߩ�d�ܘ)l�`s����5�,2=�j��jQhɊ�ح�5�Ƒ��<r\����*��T�"jo��	�.��t�L�ڐ=y��'��^���!�?� �U�AJ �)��k����e��hxKG�Q������p��ipP�UE|6����I�e|	�M�������Y*w%�U�X�(/V�u��p\�\6��ߦg�u�X$�C%���:�����cRٓ>���!�=��6ͪ�i��4�Ɣ*�s+�B�{~b�y7��n�&2��#6�������fToS���ʎe�Pa����uAF�fU \��9�Dj�=�;�+{��R�}\�|�z6�m�:FR"3��w�����[C8�
^��?"����a��۸�C��pZa5��/~4�s�r�,*���|��QUu�Y&���p\�#UJ�f�V�@���2�d�_ǥ�y)o?����|�Ʈ�v�pz�g����Q��V%W2M��,1<9T*V0Oc�̓�_$�h�w�Bc�ҿ���Ƞ��_+����4P����t5/�F��G0�6����b�v��^�5w�����레;C�˲��� K�n�F�g_����Mir$򀯐�[��+��ys�g�Z�-)�>� �
V�g������A��2��*(N�"�A��o�t��|��/��T��k ���|�z�R2u��#�c+��9q���͊U���тqxZb���O'�<'���Ӥ��"�YhVH��tS_�GF���T��;� L���A��~�41q�7�
�����\�����;�Z��5		еX�&������*DAn����a4�A9��t��es�8M?�_�aGu��X��Vt�۝����ڡ�
!%��C�ң�yנ�{ �3U͹��i�.2��UE���@s�e�~~2�z������Za��B>		�I��$�j��	�v����e���f-"�X͚�aHZ�{i��36�a:Q�r�یw�g9��W0ӷ�F%<Sڷ�Db�u�F;@D�*��[�� ��7�w{��%�~вC�:�>I�9۱tw��u�@WA0��LL ��Q1�N����Tܞ8��[׷k�ÞY�=�r�Ota�#y�Jyg%�I�~�rCy�>9\��o�YJɷ���>>w����6�;�t�!�pʯyo��\fF z2�tj(Z>ka�s��иT\w�����lqd9[30����;2��e�V�{�V�qL�}�c���n]�h���{E#�+�/\�s�rS?�A�&�aV�^3[�O����|��"��3�i�F���u�:N���BN(rd�$�҆�p?��y��.����n��������x�x����Y�A�s��%�<�.;v�i
>���X#��=��A�����7.Q��kL"���|��Ln���[^O�����HxX�!t�����u1�L=�%�JdX��,��}�_�j�?O.�#�Z�a���:��+sȬ_tp)���ߦ���)[#���?�>�ă]�&��J�f�Yg�%���i^�W�(씸 �x��
�uP�9�4�ż���fI��$���5��bk%�<iq�Ԥ�"|QXz��..�e�[����f(KE:'���4�_�Tъ|U�W��?*l
h)�C��gݎPbJصWc��u%Y�÷�Ec��;����E�(� &f