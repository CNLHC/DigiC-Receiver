��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���8}6l�����"-�Ɓ��i3���T4$L��[�	ݤ1ד��v)����5�K m{8��u_[cQPL{��8�� 5�+���K @-��,wc�E�k�ι���3�ju�kg�;��[*�3e� ��9��J�5PG����T"��)�f+2]V��E��z%����7�6�H+%�!���e�F� n��(��cC�+8P��Vɗ�ଡ�L���udL7RR&TĚ���� ��������>s�$jD;�ܓ�1��:�Ա��@\YHD�#ɧ���h���M��)�F��@�:����ӒJzv��kbe��(̖�;�����v��tE~��ɺ>k��@í�`���;��&e��-�iď��B�s�@&�Ƈ���v�a�{�qL��:����G�>���������jD��P�Z��h���!�o޼&Sټ�c\O�w�k2�8B@��0��w�2a ((�8��E&V:����2$B�@���&q�<��b៳��򌇡�Abq��.;6��Q�����lCF��	�F�w��
-�	WC�<Ҙ��������'B��~p�=�4k�Z� X�P~@�6���������mA����W�҃�����[j�B��l��$,]�E`T�
�����c���N������{d�e����{7ݶI@[>��.��2B�q�>��W�z�.��A��򞧂�����'�`�߯�4�=T�bƻ;mQ�0T`;�����1�?�;���)��G��7�kv�?<���ެF~��TA��{^6��(�݈l��WϦ9uJ��vy����+�]�''������"pDc h%w��;���H��:2�o�Z�_Q�.%��X��z喯����S����sb����!�g�[["����C)��Dd�n��ET'9 �X�<�5�taܚ�*D�z>)ٰ_�2���k6�����$�#*Wbؘ��l;K��7�_ϰ:�R��l��p�}
����)NwC1fNfÖ]*����#�Nm���3}y� F���T����+�8�&)��_�����N� 47J{��[0:��Ck�O�;�ºF�`�����<�����6���	��H>^�am?C�vk⑾hF̅���O����X�{�U �4��d�."?mw�S�z��&0��\�Ɣ�0�O���V�W/����|�Sj��|B�;��[�B�7�ݓ��FS��@4v ���}�}��q�w����Q��[c�A���f�|�_���<u����,�Ո!{��)=� �QQ�HT��;U� o����g��Qyo~�B%(�9�\�B��})���IC����a�m;���k��������~���5�� 0�hJ�T@)v�\R�Z����f�O�ҭu�K���.5T�I�-���ex�Bm$�#\���m�Հ�K~�j6~@�� ��lRm�b4�q��|�a%�M2щ��L���fl���ǵ<@z��F4 }��f��w�E�]M*�=_�aUh��� ����P�҉�nf�
�̺����|> �6CD�0l����{C�V�2���Q���D��~*f�#ٰ��[�F�ل����}c0�A�r�U��6�c_v<���ro�T�(��J��E�M����8'�2��ˢu;y����+�U������u��>����?���x�H(��?#��-��F������C7��*�ľjɐ_]�?�����C������[/P�8 �l`��p�R�-|�"1Ik���n�Te������2�V6�{;�^f&��s�uЄ�{U�{O��ż��V8�ҋ�a����RY��o�������io��IǛQ79V��#�5:7��_��)&Z��֛���*�9����DQ'Gx�X��t%����D��Q),�����C���ϐ��?�E/S6ߏ���ី�n��<$0H��m��9�����z~{;�4辡�F�����Fz�R-G��������΂&\����/`u�GB�c2�	��Jp��?�������B��':G| t&.?��g)/xEOPQ�rڧ+f�a�i��M��A�������a��3E0^R�=����mZ*�m�C�t�|-G�"/P7~��J�X�[lZ���_Y�|�6�h����+�#�z�. cV2�烘�ݾ^���\�x�:Ӑ����^ĳ�+;��%��嵮��
����K�����Tٶˀn��길�G-ӿW!�zHtb�q�И<0e���B�`ꇐ ��%�T���3<�۰:-���/㝈�4�DT���=�7�}�~�ϑ�����نT:5tI5F�~�2�\hf�X�c� wq��>ɗ�,"��;�E� �(?o[�Q/Y���������v
sC��.qz%`�{����(����p�K#����X���o���.\���_��	�	���~ݕ���bF�T��dDZ��W)GT�'�vgY+�)��%m��v�t[ :��Y�o��B�=ZD�0��e��q�T�os2�aT�i��R3�~�o�߆�%��cڲ�yM?sD|4Nx3wO�[�<.7?<^ɓ�@0Rm^�?VvB�F���j�9��
�a���,����]"���c=y�v�&I���i��-�4/�݃ި/PL22?�~^ϰ����(��iI�FX�W������4��T��w���*�@_ܺ�䤡��|,ZKkh$�����l����5m�|�G��6�a�+~ew*iv��s\��I���ù ��S>��٫��l��t���Ґ��?|����{�QEE5����m�n��L����Ge{4Y�����d��s�(b�Pm��ja��d�>�
w������JϾž4���_Ƅ�"U;�H���HJ`{yS��ʳ�C)>���(�`����˸U������9��d�d&.��Zq�����X��;,U�Ps����.���[%�E��*���m2�a����*��҆	�͓:��4�_�j#!FX���0\�)Q�S^�TRu�1x���xHH89x3��x�e�����7���;��vN�}2�2�y����,��B\��^��pW4��,�.��U-�a�o�Qx� kI��Y�K��U�0C���
��T|�6eo����Ɉ�*&�rw�6k{U�j[Ɏg�x��bƁ�CU�tpͺw�f�?i�3,��*�j�����z81�5�퐇�����6�`< U���N:�6�E}=��`(W4I�^��w����+�+<ſ�����m2���$�/	d�]���k��g�>��Hc^XbA���/�ysٹ�-J�(�?�)�����H�"�����)z7��S�o������xC�-'E���WC�H8j����.��Q9�yT��@�uL�����CJY��r��c��R\�6���Z��[�`W�#+�c��o��+��rq� ���)�:�𽙷��쬻D6Ue�}H6�8H�S��bA�1?RΫa�%c��[�m��4��fI;#����<E=TY���`�G���u���6)���م7-�Rk\K�i�m�Ba�p%�N} &\Nbz�u��Y�N}Ny�n��a
r��%��������ݠ9���]�/0&���:r�Jެ���7S'_N�'<�ټ?������pN6<�"iZ^��Q����/�����KyWQ�N�$Ə��a`�>Y͝R��ˡ@hM��=�aM���d�� ��oʵ�A��J��7k\�;��~j�)��F�K�Y�C�����0*o�[���n7��`J�݉���h����SI\،�H�hUZE��7��:�X�Y/�����m�Q���S��t��xpq�"�*3�@��M�Q
�ۇ�zD�)���Wl&
��#}DI\��Uk�Lf����I2S�����J�@|�}ڛ�I���7�y r����H~<;L�"�M��M(
�kC@P>���iU}�k���탺zn���˃����t�۸]�g�x�B�����d�*��(t:�!Ob�G+���Z'o�sh��c��t�p�i�gǽ��r.�����H�@��)4�U�!�U�,SRd����?&�k\�����?����G_LERR<���^��Ʈ� �Y�@���;���P�_�>�"y/6đ�LN�t3���f%tL�)��]G��j�n����0)f�x���Y!�r��]�.��x��Ԗ���*`�m�9१s�}L�5zzО�U�a��/̴)/�AEO�l�ʯ��R^����}�+��'n�rC�����Մ���1)8�Y��:��['>Y�$�����i8����А�9ת$,�R�D2K���Y�=2Ҙ��S5�5�A�q�����4��GۓAR�2�����n%;l����P�KjD�ӷ}r�`��$	N[�v��A���������@�}��b\gA�ڋC�yɮ?q}�V���0~P�`]�)�G�]2���B��FlD����$�W�$/}%�\Xk�q�����]:��FD���:\r��#ǆ���[�N��D���r��5�;��F�TC�mes44Z�{߮��h�r����i�
��1ǡa���˸[�F��������WTx�_.��4R���>_>��C-�:Q��Q�_��F�6�<1�!���G<o2\S���S������[:j� ���-Z�qd������1$$���<@^����l�ݟ��?9԰E��<8nD�<}�t�(a4�Z'},��\�i�R��s�}�:m�b3�~��Ce�]����+#�d�٩�Pۥ���.�ķ/4H��<V�Z�ϧ�&"frs����#6��\��I���gxJ���L�Ux��s���ām�=�r?��x�Y�� ھ�ˇ��UA���f�޳�����:Щ�0�����iE]m�mz�Ħ�J����z��ijV"��0.�kb��
���;���{�7�˂�b��� >���b�%&��\��lp����E3d��;�:p����	)�<�O#��m ?;]<x�/$�ԙv����"�*j��X}~U����R��J�.�`���R�t?��h�B�@�1�%����;_�MBd�W|�Ϟ�A�io��A��|������L �UԾm27�j6��W�E��I��X�r-������=�*��J��A���0Z	V���'�w<�GI�d��T�k/����x�� �k�z���	*&%K����������iq<
]g�)�H�V6?�}���'��?����� �FV�k�, �㕟(�:�Hk.-Žw��{+m���0�9����BAHs ��K�d�$��l�$��8�Kh���|:�=Q!�;b�^���τ>jQ�%�a .�[
�3f#��[�:Ֆ�^É>�/-Os.3�������X��qnB�e	���1�خ;}����M��5��@��"��Brd��86�=�/M	?t~;�����H����D7R��B�����s�� #�R��[ܢS�r�ܶmE��K��1ġ�]B�J�f%G;	w1>�u�G^*G�^fAU�X�*Z�ݬ�� �6�}�m������<'zIݖ�A��6� ���4Ӊ��NKh�<�8����^8:���ՆI��m�!����_���ۈ�����Ŕ�_?�cQ�=�o�7(p�M���O��'c�yFZ��S�"�e۠�Kߋ��阣k+c��%B-�E�p����tE�$�� k���k�lN}��G�v�fњ/��!̫?���<IK�����
�Q��i���Y���-�*���E��!�j���KQ��B�D��+U�e���)d�0�&S�m�s��X�-�ܷ�A$Kf�R���U�̵�x����V�\nٙ>Bx0,�t?\y7�����;ZF�,w��@�͋.�&p��Sg�H���!��>�dǬ���R�3�ʡC'�D�T���CI�;$اг5
�g]��A<�x���#��htT�T�P�V�lQ���c��q�峞(k���6��� ���`w+f%�Q�}�bQ|�u�{(#�QFj�b�ݱ(@��v�K�(��Di�b��l�		Ll^�^E�N��u���GK���$9��� ���u�Lñ�4�qe�
��X�7�{�L���y)e[u�{��@,�EM����CG�D��Υ<k2�վ����W�PEx���x���>V�Yũ{��x�p�������J��Ȁe��;aE�o�"c���1�E�y*�Bʶ���z��PfJ�Q�P�9Or�N��܅4�2'w�	�W�5��?̎�b[%�[*j�}>�k쎑�ͧ}0����zf$�n�	���Ho}o�e�WtvzB���AV4�W���IGM��S�H��O�V[�,� ��~7]�'��� �z��~D�v�Kp����R�@e�l9�:Ģ������YO�o�T�f���ݜC�'�GX-�1���mG�Q�>3s����8�;s?�0*ʹ�ۃ���q���/�y� �v���	pmN��#)��4��਋���1X	��2D��w�)M!���3KfhPȏ�oM�"[Ȟ�N* |~B��j��ZT����֦�E��Nj �W��
�s�I���2�����)����2˸bD��vա֜Udn��[(x�J�	��������5�y#;o�8h�]/��A�4��g���15AԨZ	LKV�!��4K�I��2�/"�;`%���ןn�gZ]��+1��qg�����}T�7zjD�\����eQ�Pzٕ�9㤀Lչ�pL~�D��c���դ���p��δ*����u�aV|_�74!P[>ŔO��x=��a-y@>śAj��Zuro�����p�0]"O������W.��l�muyg%T"x���:�
�!��#Nh^j7��Z$`�,����}����7Nu�r�4�[K{�l����	�=�+�ﭳ��
m��}�=�ж�R	�a4Ԥ�7����F)���$m������&XE�+�������1a�g$�u���G��F��i��8�@*�q�Z%���������Cل񔝝6���e��3��>T�$V�\ԷғA�Je�������b�,C��h0�� lz�g��掍����F����n�'$��ر�^sB��cwJ������A��u �'��W�`ݾ	y*j��V�
��qL �������Ju�_�������e�3[�u΃R}¦	�[�|�p�!릡?�����2g�{6ԞȈ��1�Gٲk;w���N�gOc���}�E2.}��d��ח��G��2 �$7�8t�V��AǬ(�>�վ�3�8'�3�2����.�I-}����]�U9X?��,k-�P����G�sM�H��D
]UE�06��G`j/M�����,ߒp1{QUn&W_��&"b�xhm��rWg?D�g�p�#���>	�)������j�+�2V�r��B�_�+V����n;Fo��U
բ-�k��X��*0��{��~ɋe��~�0w����RA ��Jc����Y,'��rto��ciyѓU]ۘ�A'����H$p��R����;r\�e>����Z8��� D�9�GZ&�r�r�:�ߟ=^�<�t�_�Q��*�q	�Fa��W#��IJ<ɉ��p��[�NjFG��{�XfI݆
���W����Ux`(�I[�W?��Gi�8�lTt<o�����O2�T6�=���q�����͗��[��U��Ʀ�gw%܋�����(�T^fR�����X_�~���	EO��΄���$+t�t����^�R�Aݨv5�	�I����� �l�ʛ��U٫wu���ZE�����VH�p�.�4�A�N$ʝ��!Jv��P�+�Xb�)4K���8������-��O�qy&-�������G�=��W^M