��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���8}6l������w˝���q��"*aCQ{Q:8Ts��E�<�~�"�}��4 b�A�����zU$׏��6�5������F��~�qƣ�7��^�ۍ�
c��E����h:W͕�>(�D��g�)�u�ڮBs:�<U�<�?L�_RF�������C�+N�~��Y�r�"�nWP�y� )�[�Y�aa��-�=-趻��s�c{�7*�x�3���e������m����ժW������`Ugs[��cf�������ncηQ�������(�ҺV@3C�ğ�fK���/��oX0�f�.��AN>R������N� gg��u�������d2U�OD6K�}�F9p���ͩf-Ϟ�Nb��Wb�nR��E����Z��IIpt�;+y'���C݇�Nj׽�=v,�x����ŎNռn�m� /�X@�et�("7��3��Ճ�n���M��	��L�(Uk���$ �$�.����;ᱹ��Jw��`������Č�-���R����T#~��.�p^Ѽ@7���_Z����'���s�fqRQ��&֎�~+s5辿׳l�F��&�J)O�!J�!1��B�pI-|��Kq�:Z�P���|��k��?�Z����n���~��=1���fR�y�H��`�G�J�>9K�e��	�t�PTE.lw��emZ>��B3Mu��5��%q�ޛl���W[�˄�c'W�k�v�4e��ڏ��E�Y��xu~�E}�C�T��/����=-��`�Z�$���z �iYV��y���U2�y
�l�̔�CX�^��n&��Pz�7�]B-uU䅵�����R����#}�dV-���g�D9r5���i"|9,<r�������������Ι n` �
��Q� 6���xC��q�E,C8{��h-f,��VVkM��V蕻e�d�3�L����)m�G��d:�pޟ򋒇+���d��@�5 ��诎iuHs�R+�����x<��d�j�T[���{"&�@�;}9m�F��D)���JZJR�6}�(��=�h�6��Mǫ熒�����~$�]��o�y9������CV ͙80�X���k낀!)���љ��ޛ�T:��?�6�,�t-�L6�un�hI�>ŭ�7���D��eƻ���"V�"G�q�#�4"��"*x���;�(-7������)�ڔ�̻��5](�s 0����J����w��s��*��_��(�4� �fʮ�C��ߣ:�E�u��t�3���qL+^�m�������`xqv�A�_f?��s@d�tx�ZƼ��D-S���?ۻ8���|e�O�$�Z������Jsnd��p��#$�8��h�+M�V=�	)Ƽ����w��L婛G0j�/>/3�p$,I��0�������;���F��v���b\��ߤ���Τd�������_��0X`*E[X�mQ�-S@��d�������s�r���qeV;��_�H_�Cm%0_J+ve�Ej�т#�P��S��i v,h�I#��泗9�(A���3{(��Ų|;�(�dM��>Nrz;��l0��O\:�Y+L�Uݺ��^�y~��'�KH+Y����)�?c<&�f�̌7ci��ʂ�}�3X�����mz���ܟ�B�3�u�	3V��e��g�њu&�-���w��2��aD/ǘ�GO�{�Am��tr����,�ҡw�[�d=�y�����e�݁���W�!q�����Z�Ѧ� c{�1b���k�����R�|���@����ݹ�*��@�e �������wq5Z�'=�qx�L|m���
��֕06K(uW4�د����Cȥ�#܁_�g�,�Y,���=��.�%5Y"E|cv
�T�l��F!�Nnʕ�vn"A�T�V��M!�.B��C�o ��Z��7�`+}��ĚW�i�[v&!����X$�4�?*��B��*�%�;�x	�r�7�M0�ˇ��"��B��Ł8r4�pPn��`��C��Y<|2'/$���P��	&�N���`!�sT�����C.$�Z�lm�]�\;Mp������kC�vd����4އf��|�R��A���_Y�P13�зu�cm�[xŴ��%N^�u0٘w�x�n��*������6�9]T}TK݊�!��/�1Ł���(]k`�C0��Ӓ<S ���ۺ���^���.�o��W���[�"V簈��_w�1�^�I�m4JX2zt� a6��y��������P�e����b�X�W�=�z��2����gG�z��)a�%��2�hp��̯rց���D�WO dp�h|����4 ���s�T��Mt����3�PJG���H	·�P�}aq[qBP�����ܭ�y�6B2iU:��Db���׈]��w�>�����9&�ed��Y���$���OJ�HjS���O}VnT^Hmv���D��a,0�.%�⍰5Y�����b ��_'��-w�"��1*�)4�K����yzw5V4g-V<���&T3D초6��|y����*��=!�Q��8��Gbԏ��l0�����+x}<�,�������"]�z��,
 ��S�/d���i��ŊЛ%U��=�8�}�u���q��zQQ��kʽ$j�oY6(1���
kZ_�V[+n!�Ә\��g��$@�q#���KL=	�Z�6�T#ÓͅW:	d�"!p��펑V�8���FC4�#�_t�"�S{\i_�Mkk�����6��UaYڑ.G�I�@ 0�9p�K4�m�O;�Ĕ��z�Sw{�[x��������p�>Wm�鈴�$b�OY&" �3tX�
i�R%��p�r��%���} #�`?�(iu���G#���RG@������S��vf"��V��s��뺷/�O_��{��>����6C�U/g@��684����r5O��.�˽��/�J����+?i�1%.�J�8�d!_�B�.��[*W��ʢ�p�B�]��vIA��"��A�y����ei2$&��tL�W��Fz0k�wG��d�g�a�_���KE�� �}B嬣П|�sͻ]Re<���h �u��ܕNO0�@(���_MϚ�i�,uƨ�^&�%ώ6Y4�<6�(׈���E&3I�mx�~���ΐ^�<c���@�H�8�ѐ�����LF7ۖ)�w�����Jk���� �պ�8yꋍ_���H� 0d�����f��.��5�u�{ϑ4G?a���GAQ�����y��W��K0DNd|��O\�Z��d�$^O4�̵��O3��jY̲�����4�a�?���~0�-�z�e���s�\;�ļ0�0��T����������s��!g��j�A���pG�r ������ �b��+�	�&p$�t#�(�#%fzp�^� /^�JfoF��4\�	,���b-�D�"�;cBB�Z0S�.�P�>љF6=�y�b�KfީޥoL���$�o�1oU*Βeq�]P����0���
��(@��'��y����/ N��L�j�Z�B=��\ʧ�+9�<�f���ц��Ә鬫VWߍ�d��B�dQ��]��d-(��|������3m���:�~�wЧ
�:+<����H�L�ʛ��2�RZk��2ى���0&Uxe�e���\�[U����J�Y�=��,�@I�F��>ja��\�,YB�z�ݔ�+O��/;�u�WA�ƪE�o&���1}�f/o���AL�b��;�n�l_�����Թ~��U����f0Mb�������;*[w�wFNP�gH�����'MZ��3�WkQ�u��r�͛N��4쓈2o��d�j���lN��	�������I�Q7f)a�����jԷ��g���G_���3Z��R��d}�v�Z���U���0Щ�D'E)��m д����~H���W��y$�/����/4���B�6xt��2fi�/>M+Vj7�WB�����
\�Q�H���exF����ڑ�S^�o�5��2��%Q�PK)�l�+��8�9�F�:����ְ���������ۛ
N�L�����u����B��3�֮��J����(V�2oƈQNk�e����qJ4�A࢘�>;��-��e4���˰�	�c�~�r�[��3�.xd �	��!@�.F�J����	k�Na��*� S2B�!�<[�T�~<�f�.�<焾�g�Ƃo��O#�����}H@S��͆���1,AU�(��� ` �b�KT�NB$�:o��g�������ğ�L'�/Dg��B�
܆a���h��7Ň��lA�)�g���߄�y���n��1�2���h2���̾�(�5�Z뙬�L/z*��.��#\oK'Oo�ץ��0>I�I�����G��-��t����J��+>�0șM�q-��K]AY#��'��ҡ`�	(
���lˁ"jpD�x��% ��[��>�<bϠi;�����l6��\��r����Ѩ�p/A"�m�b��;�B��~�L!IkT�_v�e$�Я }b`9��l�A�����[�6z�(�K$�zuVQm0�"����|9�,hS��Mtm�v!��.KK���KJ��(q�����U1�U���X[�0W}.��=vW�g	
�S=��A�t͍_Ӻ|?�}�f`z�&/��Uŀ�&fxڈ#Pβ� jڤw���a��3�'��ܼ� Js���>�q�0Z$���ϟ�|%qI����3u=�^d+~kʪ����H�TJ�keW�r[���G�AE�	}r&��3R]������I�x�&g���,��:<aN��+F�]F�C�U����E��ݺ��=�kFK�D�1sN8�����Ԛ��B��|���M�W)��<?RBmL%�m��ra�ْÆ��%YD�)a�B��Z+�������xw�/��@)�CȠ�BX�p��:+i�5k
#�n�&��]��'���؜G>!����0��~a���4q8+@��-��Er\=�m|J,��KN$�Mx�*p�Z덯7�[o"��.��V�u'��Gǥ���go�'Gp� ���a��U��.gż�9R��ݷ�鄕�Eű�w��)�+���2��S��"E>�9��d)Z�r?z��j�<�����M��@���`�w/<��G�cBp���wHF����%
&��8
j���BǘW�(T-��&�0�V�=���@�[�]��i�aCd�A9�c@�ͺ�^s|d���)l)8�3���<7��^�%2~殀p�K�?�Z��KA��l�I�4��@aa+������$��q�F�H� ��_	�,o��C�*D�i��� �&��S��t��b",��׻�\�W����@� 'r8��>U�W{m�oسW;�-���L=u�QP�.˯m�4�X�[�� "Yc�
����.*w�<1�g��k�8L}X�?�"�G*���?���G���h���H�p�d�X�ǉxR�d��	,ǺVx�1��@"_X���6��ݱ9�h�l��x|ZD0.3U�#-32���_΄�]i⧤��&y�rgp2��z���Vՠw$A}34��d� ��Ѹ�V6I���Z�x�F�pY�)2����jƨ�>�R5��f!&;�5t"��|]m��p�1LƦ�zx<H� �H�:T��jm��+�ji	.r���}Y�e%�2h7�퓢��M���Jz]�Q�o����%�����5J�f�?��v��rP��|��C.�������JPY�i��#7<T���s�F������	L,��1�D1 /�p���:7��&y{��/����q��*g T�3����b�D����a���Q��SQ/C�^�2�v� ����&Z3�ť}H"%�^J�Q�2;A��z�9Y����Kψ[򗷅q�Ԛ��Vڲ���\��������O]�e���+9����ҟ�#g����2:��i����w;�8=Q���s�Ư��
/3��۵�\��D��^FQ�#���U�L����hE?1�/]E�1���]��q� ��r��x9��*>�8�3�qF�ʁ�Y���k>V�!�L��D���p' ��Z�����`f)�F���^3'��g�h�x�cg��U���?�UmN����ؤS:�c��>`#jF�����^o��?"���E�����>9�Bo Z�8��u�k�V2�eg��nRMZ �r�3/�]���;��-��O�����gC}=��-�#�0?2k�k�;�HX��-(|�3�x�l{����	�y�$����(1��vѣ63�J,� ���6�����.��;hWEkT���/J⹬}�?j�a�;Z�ǯ~dH�jk�Q߄��ؿ����u�ꘓë���}Hꞩ��6��7���x*BN�݄�����|o0NC�̨�ӓg�,���^@�<KnJ���~�Kz�r�B�e�>~��_�`B �0'�&�NEo�C 	bGk9�囡�wMEl�Rri6����Ĥ-��A��t��/4�j���9����҉�p3����'#��%�nX�V�-}(c����٩5��@��`�P)<���ԙC �#׶�<x�"7��Z�zX�4UG�[+�ŗ�|�z�Z	��$*"�r@�LJ���Pm<�ySO/�;�3 �ė<��/D����ՌO���0���P_��ې$=������760����De[��P2���=P;��^�d	��
#8�.7�o�Փ�W��".v���.c�䣬�u�S	U(�=�F�,�#�\�ל2���5�Xw�,1NzvH��X���%�@Pg���_X�|��,t���-g���V� sԯ�C�%��P>����?!�O)N�;KM����փ�e���E?��4���Wx�s�f"���vh�T�ߢ���`�g��Q� JjM�*���J8FZMi'z�=��?W�V��`�`VBR��aX�UA���A���k��k4��g���mu��lR�@�J{m���.<��BO�$V'�*�2�	���i�T���.��!O �v��v�ۥ3ˤ�adZ�n�̅͝�&V�cK�;��YcBS�5��/���Kb������X���[&��ˑ�s8���a?E�BR|H&��U�7���Q0Ye��.�ա�<~A�5��cı�kCu���.<ÜF:��Y5wS�se��yr�W��y^��Zu��:����rcv �4m,��DQ4_�[��݁�%�F�����o��"�u�2hY[�S��s8��˶�j
��Uz�=:�^�i!�����o����d��;�g��MFQi:  ��Ԃ#�WH D�2AS�����!}ζ/�a�-fL��5b��汋�:h�{7�z����ߡMܔ�m��	����Y����Bl�.An����C�&���bn��Fv��-�)�RE��N������{��l,B�!a�[�+n�Q�jp	����ͫL0��՝�$~N�i� ��@��ƹ�L���	u�c���D���fI#h�?+��>�_���Þ��/2-�yX���ϊ]�{�A�۱��(v��i����}=�5�lH�[�s�e�o��_ ��
�T�b��zѢBx==��+#K8�ر�~g�w��;��V����~�L�:
[~kr�%��Iv6�;JvED�����
_@��	�ps�K/��rz��p�_ߪ?˧哺��d9Wp��u�g�el�+�q�i\ �O��S�YrgY��6{�b�E�7���n��x k�_JS��D�s�A���j��Bb�4��R��������
�l��|��a��������gq�|v�wر��%�_�M�jRa�,mir\�W��υ����up�ݞ�:�*9�����BjF�5YH�>��,x���f\M��v��,0�m�/	FJ�ǃ.k
(�v�rq+���G��(�td�K��O-��*e�����\����\i�L�{��N<�^�O���s�Z��$׺|�Dy�m�T��eOs��n�>���?4M8�q^�/���}W�^p�Z|��֟�ԇ�.�����g�.�a��EJ��GT3F����q`-��S�g�R{�L�;h��PGh���_X�2x�qD1��"~7h]aM*i��r���|�n�Xt���7?��º@ux���t��CC��c8�K�M ��ӸY�T�.C.玛��V������~���@��u�OmwF@��;朡pml�wtT-�(��uS��-��Y�Vǚ������۴�K�`St��{.��C$%>"}=o�,:ј�0�� �!�����{�\�rMy�]
��t<��n �1�Nf�>�8,V��FA� ^�qw�閣�����^< [aV��\����j��<�����5���T��6�?��W��,nd_h�U�-Ɛm�:>D�pX���9w�6���d�d�KJE[*o������
�Ȫ�tʓ���=��k��j���+�TCy�>��Q�c9�M�Z�ϭ�a�a)pI}���3:-�G�<�'��W�z1�r��o�O��+Gis�S�0�bd�d�B��Pba Q���*<0}f���ֈ���(�ac!��mT�K�.�3�=_�\>���q���?�.���~;z����+O1��|M� ,���/u����hIf�)�Z@t�EhjhԦMR�4��-�﻽�/��
�:w���-]��-�#٬�J�q̯jw��rz�����y�~�IR�p���Ư s�f�`��6r:l�f��x�w���A]�� r'���\��yY�x��v]�'[9�Y�:S/SR���gJ����dX� %�goa!u���S(����±9��R{��	Y�0�&��ɾ�í1�F��K�4���,5�������.��yC͢F�'඘��BڒNM%-�#%.�bd��5K�:���.���`J��Go��TyK�$��s	�,�W�ݒ�CT�C#�I��oIS��!��11���*0ԻU����d���᧨`|�_ʠ���������v��!�˜��*��NUD�~�g�M�-��-m�ʯ��3�9_���g�Y��?�'���)�ԽE�b��Q����m� 3y�GKq�����i�� -���cM�}hw��
BYo�a�u�8�ޱ�[^3�Yg�RݒǕ�h��@�U�R�����x�`\W �@yS��Y�����K;���� h�[.	45\�+7���FL_�������w���|�ch7�_̣Ȍ��,��^��
�2
L������[-:�x�����l��yyyJ�(o�����V�x9�Up����7���?��i�44��6���2k�P]��:� �E�~w���0��#	���@I�Cud������`����ÿ��L��i#'^@����S���&���n�`�k����&Qp��-�ľ�vb�w�EQX��M\�-m ������S��M�B���C�e�#�߃�O�1BJ�y4� �+��ٺ#� ��_�d���3������}7NH�y#(h�W�+N=
`��a�V\%��!v���Wч�2��G]��[y�B� �rּ�ӘЊ�8��@��O��0��浦�Jj%�������\1@a��9�?�Ԉ��2�����ڍ��&����'�!=��O��JC��,�I:O�0�MgN�ෝ=aֻz�!�rE�p�p|���W�RS.��"��fR&������;"7g��^ ��G��^�yȭ�j�-2.j8񶔸K0��%�6>������g"�5]�a;e��ͅ�3u��ԡ� 		Lj��B�V��f[+�:ǡ�Q+�^����o/�}x�<h�>������"���f���֫0鱎8TIbL�O�v�/~ <T�v�h)�W���SI�9�nR��}ǋ��׈Y5҇޽�.3.]�}Z3���b�p�I�)[���G�f���x����=���~��ߣ�dj�}v�L��hf�X�ϋ�+S�R� JP�I��^sB�,�1�ˢ����@���g�윶@!�Z��V�Z�	
�E�R�V�bb[�-�<�M�y�w��c&#6��X*�\�r|��w��J����zBܳFÕ�z�<9M��hv̠�QB������!��4�
�82u�)�T�75U���`�����ڀ�m,1$���>�KÍ$��MR�La&�HIlIGXN�W���[���',���
Ix(�ػAgG�����\�=2�� l7��t�6f����v��0y�.w)�/*��C�"��#w�����W��9��Ҁ@Ɨ�2���JU�o̸���]�n�t���fAv��Ͻ�՟���J��>Fcu >rJ�	�c��� q�l��'>#��� ���݁�K�ڹ�iF�:�1'afW�юE�zJ���9�	뚯���V�X��C�Tޣ�.�v�f�DE�~��_C�����)5S}���w�ޯ�b��������5ty;RZט���\}��eN��cP�JV�&w�u�)���L>����v��Ĝo9B����ac�o����(�{7��G�D:4�%�������G
�D9���1��{+wP�PDK�s|���7!�X�Lr�sn{�iи6A�W�o�w�!S���n�~�����Y�T��T�13 4�����/R��䛍~�?�&��V,��/��[n�z�3/N�1�o1������m�uI�Ao%���kf��+�^��T�Mg��,j�B]��ɭbZ����.�OA���Y�ؐ1��9{z��}����L��Q�[T9z��kF��uXK���di�cq#�T)�3�8M\���Pk�G�礉ИS�4�H�.�,�Xb�Q�`7�~?���E)MX�/X��p���R��(�e\Q��ˮG���k��xs�q��ѵ~+�SGVM�Ksl�Xp+��%
�_��% ��K����g��`|MC�������ԣ��U��Z+�۔�,�������5r���J�;����u*��B�Z��N�B��e ���h6ゖ��w����ؤH�7ɾ�K%�eǊ�����-��J���r�\=���e;����U�*쵀C uܡ$�Vψ��W4���.�����9 �~Z����~D�I�i,s�"�7^�9n��bz՘��5wэ�����6m	ȇ����b�M��ދ�ף�k�<B�����L��,�񧇵^�
ҵ>�%��N@i�4�JM�-j�iB�����p���n�'d")Ib��^�vQl���j����M&�'멩p�3�!���~1�Gj�H�k���c׻R�u��+�z������F��	��+:hOT�ujՙf�yT2t�)��&��m8R}���������9�յL��"�	9�}7�X�2J}�:��-I����J~"A��{74$f��\E� �^E/0�:��Aھ���ڟ.��0�a��0���6���a�����k�yA�bU���7�b��w��>_��헫���$����PC��>�0���в����EZ���ȸ��Ś6gMu.51\�,� 6�ڻL�
o�E����0Siy '9�ٓo����{�&���h�X�c{�f�`UX�,_hGJD�AH�߯�[\�~\(I~�G�5�ۚ�:��͇�Ʌ\Mi��]0���c��s�(`^���GЉ@co$00��খ��"��w�k���M�#�F�ݠ`	���[�y���w/ᶊ)���;�6���,���>޴ɰ�u���D�e�3����m�mp����3���k�Y�0p���	>;r�p����{��GjAq�����>�o���!�c���~qݤڷ����Ȁ�<Cy���mz��	[GvK+%�Þ{�)��������xy��oi
AsD�HA=2�=��������4ZX:7�B:Yp�6&��!BpQ�k�!,
:������ng�:+�*���Y9\� ؆Z�LMB7B�߬��r�q��n˜^���)��#[���c�+E�
�Ů����h�p��8�H?�u���KY����e��ѝ~��F+�kcs�aSs�RX�p[����;갑W�T��V�d�8XO�~�U��B��Y��H�#�[$����z�~:"�Z�Z�p�n<mq%[8bi짳���NS��H�2����:�����A���r�|̊5�j!��6t�Z(��y8�,�$�~6���Jk���kN�O-�S����>+C�H����a`��M}l}|�Ӄ�J�D���K[����s�^?�˽z0n�Aމ���G'�"h3�=
-{}!NA�*iw6������@;R�U�/��ֳ��i���eJ��.��ͬ�%@�M~p���X�-]���<2��d/�}��Y�����֏���a�4Ծ~��W��)��( ݤ�07C�Zf�����}���&��D�ؐӊlcZ��;?���������'����{���eg�,W9:�傄>�$�e7vE�q>	q ���#��VM/�Ra��^*KR���q���"np1|�t�ޅ�X���_����T���PB0��~�dm��t�X(�k��;w�O��CT�]�PKV�~*�0�g��b��R*ֽ4���'����������&Y|{�s��!�v�ȿ�R=K��۰e�PSa��
�2��q�����?��=����Q�) jA��y �iy/F!�a�^h�e�c��Ōe�U�P-����hS$�φ(@&���J�W��zN�i@���P��pݽ	��4���vI��Iʪ��>\��;
�
�������h�\�uIH?�J��tup�p
)HLPg;Mg�@!Ѐ�n���~���Z^����BfG�|S�	ě,�q��ψ�f.*.d'�� 6nCo�@��#C��d�HS��Z�"���P�J�:�J��&8�qq��t���"bٻ:ͽ��! ��w�b�N9��f9��Xq�/<7-�#ۙ�,��h ˝}���5[σ������6<�W�6�����W�u]�E&g�!��N���VG���0:Y��gGf�u�@��T
�F���#�I�}�j̲��^-�^c�9��­����FF�4.��~n�p�$%e�@�^20���H�l������ա�i�B���NIb*�Vi�\�陫��%C�K@�5^�Zo����<��������ۉ+̂��Z��!���Ib>���R��V��"�Gm��
�1�if�D��c��2�T'��.�Rr�q�O�ⱎmb++\!@k+���Y�49��(�����J��a/����Y�"*�
ϱ�;�;��n3��oJ���#���y���C����t�}�G�q7n�;=&��k�ɸW����8z��9�&�@��v�s0 D�_2�� �ck�|��B!2$pej�33`�o�ÿ�	��u��+[^�\�h�F��(��6E�s�԰�,���sgnu	P����G%L>Ѿ1]�3gM��:U�5ʌ*�� ���7�5�D��vg/�I6��"5^��	W�||E�dvc'rI~�I�I�A���!�
�T�鏼�gc�������K��4������l��_,�u�<�+�5�3EQ�%w ��S/^�#j7u����;�K�P���{�m]�|��!��X��5�:3[�;�3[��-i!�}D��^�'�-�}�&�P's������Fs��ړqM���*�=���~��0�&�z�`4����
���2i���i�r�ӵ��Y�d@n��}͞��7`q�O����&O԰�'�i���Ugc��6�&�ݶ����ӡ��SS�- �*�ۂ'<w충	A� � �'b�>,�Sx���5�	��+�LN���>��oP��ɭ�e�wI�5��Əi�H:���h�@���k�����s���#�S4 ?O�G��������,�}F>ڨ�%V�7M�&U@���N}K�c���������?�qr��N:��]�D�?_�������a�k����L����0��wT{�H��� �!� �6F�h.6:Ե������T�����u�!�#'I�;gf ��zm��V8#��2�e��s)wU ��@f�
N���]�L+]��͡��A��o�Иc�}�ꊟ9�B0v���A~v�)8�����M�:��f�n�7E��6%��)p�A��G�|?��D��zw���Tb_t넶��w��|���Cp5�,�_���^�����r�MLJ�>9"O������g �[���B�0V�`�4�;���`��1*y��2�՟q�P��C�7y��f��kt��T�Jb2�w_���h���4��9��0S���H�>���z1�1-j�ƶ|�}M��>�A��x�M���yyu �r��뎢cxF��v��̑#?�`t�ƨ1��6Az	��Fe���h"5&_J�:��xӞ����wW$��@�1�Q�L�y�Bt {pk�w��n~E�m����3���A�;R��=����x��S�ؑϼ ���V8����aR���%hݎ\��p�ڃ"�*���S`�UYs���V5�GZp�G�.r�Nv�'_0�8�A#��%I)�J^3hq4Z��Q�%���S�qf�L���-J��%��m�Wa=r?i�^��A!���a5˱o9 yC���.���Ӭ�8���sJ0�65�uH|��u��ڍ{۶����&1�	��?ޏ��R�U�Y��>h�G
,�t�KP������x=^�Y7&u9K?�7�rJFk���Y'����)܆~�n�6-�Ů��||��U�|�'
����)(\|�[�S���Վ+@�\R�����y�bua2oݍ:d!Y��{�A�ݫJ�@>�� ��[������5���*�K�������O�e�t��kCw�}���P��}���m�A�mB�S�=D�|g�p�C�>��/<]M���~0�fA`��L��M��cs�v>Q;qKA�_��f@.#�L)W�hիW���q�~Eo?b���:���d��	�n㼖�^i�����/�����z�����_��Dr�8�"��nB�on�9�����ʗ��s\^r	��^��j�'���6N>�5�-[o�@���,b�fx����C���gs"�g��֦^�D�(Y����,=Ua)�P]ӧ�t�<�%�sѡ��J��$�W���[��'8b�$0��Į���/xAs��I�W����^��ŵ��e�<��\pt���g6�;�����*M$a����� ����8q�q*�W�L���\:@&��Z�i��MK0�A�l�7l�uE�����i�#џ��%^�5�*P@{��n��0�fm����R������#0���s^�i�@v�QRs^�U��B2�}\@��#�L	_�wp�Zp&��kn1;*԰��a�;�IM�B�T��jX��N?]ן��W)˷��%V�����!{J#��ɻ��>zzaii��x�:S���E��5���^�����Qg��H�ȴ��aX	;%�j���g�FU������bt�������~�(��j];��R��	�{��4٥��~s�_(�w#u��1tv���4�d��C���Ob�^��������y��6^�y�W�*�(7�����B����5����W���*��KXǪ⽫��e�o��X��M��?1w��HB}?M0V\b�$�*^���=b��p}M"�=�q%(�N.�`Ŋ���^tI�nGj�Fi�Г��JL�* >��^��5��~���R-CȒr|X �d�����G@��-�A�;v��ًLk������ج�fKKy6^=A��3��3B�d�Gn�.�7��Ul�_��h�K*��μR!
�*:�:�x!«��)�Sk��ߖ�T�~���5�1�G�"��#7����kD�����żO"�*I�� -�V�Whx�{- M��ȉU�Vn��#G�/�et�:R�M]��ĘᰧO<�<#�d=q+��Q�_)�و�!�w��b���n���oF8\j+"M*.�5��1�-�B�o�f��~&4�	&��N�DZF#�������`T�G�ې��ï�0�e��Ex��J�����JV���0�*�Ѭ�(�ɼ���$���t7i}~H�U���\.<��7����`�D6�
y�X7&=N���������K��>��v�sp�f?�:���x�����yIPRPo����8�"�7��5��(«���0	��Т[s�j��x`b�p%�����<0ę�F��������9��-dr3μs�J� �ij[e\���v��5����lkVy��������ģ�pTx>�k�e*�[����&�Vg/5���x�48��p�BbQp6�i6�o�S�U\�)��5��ۇ1ԟ�Q�"E�;7#Pc����ɭ��O��~#k밸~���uRār�3���( �F$}�A�;W_�H�d�lS��-�/h#�kp(���5^F�$;@�z��;Q�p#4ZuB�%�r�C�ݓ�X��0���Y9�U�*;_uD}B)Y�XIk@^����>��)� ���F�ͣP����r��n}r��6T��̟r��Tr�q����k�b" ,��Ҟ��ʓP[��g��,�>S;'�����mns)�����w ?~h���ψ_�������0��]����v� �]�����"I���P�/]�)V�3]�S��/Oze#]�[l�o��8�Ԭ�~�"��u^q��G�	?e���yS���o�W� ��Dگ�[E�JڀŁ+�V�{�%�m�:>��������(�*�@3�o6�+sԍ������J�,Z{.�( a"��ET��%>������,�"�V����z?�T�c;q@��מ��q�5�C~���x��߅$�=x�oMQf��G[Y�2�ʳ
\��~p��������8Ñ��kE����n����:Ф!��+�h�6L�B�.��->E;((��ffp#���@����(�J��.MԃTJ����TT.��
��?d�i<�a�0���k�i�)�t��qw��`Sl��LP%]4R���9���$�sX�.������gp�)lQ�5�!r�7�
w!C���t��^�^�E�%wڝ�jW�ϋ��Q���
�
@����_�rFi�]ǽ�|���4���i��˗�r��a���ߏ�cLWmoƆ��~Z{JP�)�f?0*�P���&�Q4��b4:H��!B����H��%GNn�Q.y�������8R5l�hx1�e��sI^�(�HZ9x\d�K$gf�2~>㥖K��>X���n���f��V;�=���;4U]q]+����S��ꜽ��v΋��J+y�O�[
�q�O3�$��6�H� 7r
��\�pH��(����U����zo��o~KJ��A,��`9��"���6�H����;7Ot���miI�Y`���а(U�B�3�j1��Q��@�3�?v�ü�N���i$��c�:��V���fx�a<���UL�5�.O(������&���BG<���f����Z�u#�]wżm]�������"��=�s�ag���-�j���d\��:ݣ��Ի6Zi�HZ��dI�l���Ҽ�&��X�ɷ:&ϸ)�2Z%��"{/}2%�J�xm�
@�)ӫ�S�u;F����g�����n��8���7���e0Ǎ2����2I�x�_��Y/���w���h��x=�#�;���Pw�UVE5��&42�w5��6U.�Ij��GQ1�(֩1�E�:[��Ky���z��՘%�H�{��P���dֺ��9eT&%�������UEA;�C��yh��A9=�9��;�H/6���/�Ib �Q0��yb�����z�E�YS�)t?)9��a�_��;o�!��i*%,m����)&3����>�L*���i���0��uGB�� VB�ڥ!D�--����x{)]��;69R^1OZ=b]�_��'O��^���30!���I� �d��[�[Ȯ�=*�Mrqg\��CV�QKa虂{Q%�th��wS�׈�y[|~��� h����xg)��j���C��gm�U�vA���O�~�"(����zJ##�1 �ݿ�~�]��j��P�mPTp��E�QBcEӅ��~.�S��q;I�{����6�uJW9/3�TQ��%d�����S�"0�*"6YE�'}J�<_ d�V*h�2o����g�܏Iܞ�ӣ�W3�B�)s=$'N]KM��R�`�3P���u�]�'��dKh؁]HOc���,�4�'�67�sY�*�ƛ���!E|˯�>3��7�p��Q-�����T:����a[e{�\�!�	�W�Zw9�S�%M�g':@3x�?P1�~&���x�hJuڶ��gu��	~iLy �p� ���<ѕ��Sc���eo��R����$�8N(æ��0Cc��h"QD��H9$�#��o����=k�]?��]�Nè�J��K�`�+:��a���"�3-��o�d}SW��+<в2�����©/c;��i��*��Z;u	$w]o���
�Վ�M�\�k��6=�!��J.��w��m�f顅'h,b�i��5jB����թ��ޡ��v�-��ֽ��<[��s��`nJ@j﮴@��K���w���$z�A,N�$xT�����9K�A��F�T�_��`��j8M����?n[Rlﮖ� �Ū|�zɨ2H^�>iK��B��NK�O������P|hc]���r"���s��}��5�n�>�٣ݻ]z����Fn�$k=8��n��3S�|�:�ʹ�	m~R2_ �/��)��b��zW���p6�
�oI�Z��Ų'���*I�1Y�V�p�m��rGQw��A1�4��`>�.����00��tr�zE��{�x�%���d������g.Gt�jP!�u����:�ͧ� ��+kd�?�>��L�d�5DF.Ӿ��Mp"�Rrk��5O����[�b.A�<~��G��"g�\lHQޣ�Mc�V�W��&Q��3	�\�?e��7a���W8����m�j�
]��x�a�>����%P�Y/Ҁ�.�)X1�5�ȑ��>Q��V��R������vDs���U���.K�͐����r����G\-.���/���~�Y�Pf<K��1��c�ͻ����#x���ꡦ�}@@�'����s4'�a?
lV�H�mZj���K�xOЫC�o�&��L�֛^�\`š=|�C�$��Ą���F����1��7o7�.'?���� ����1d�p��#XZ��zKX;��
����8T3Y*������U��`���
�>D^�m��ɚV�G��3q���b�z�I�R��ç�B���I���u�\�k��4��Ȟ��y��i�ɺx����Bc-2�6���js&	�<�gaO(-���
�	��OH��*f�~�$[�~��}�CG�tX�պ�.4%��?�F�.1Ŕcq�t�z|$`�"�H&َ���N��Lv����=B��O�~�7b�Pr�N/������:dM�xP��X��寮L���wM�� ��o�NO�����7KE���/o��o���V8-}��@(H�?<(9���4�.`�4������;��p�t9a3+a�<[�T�w���ڰ�G�a?��f��F����'� �t�'v����>��}���nr������Ř�������T<TI��ev�`�|�!��G9�{4�O�mOYW�20ꝧ�?��-�rwj���H�6�x�Nɳ0�����д��{��� ��s�fk�.��Ra�+E`���$�w%W�4�uD�L���06����A}��:����Ə�u��r1���s8����"�/ƪ���7�ʼ��a6�j]�&��s�$��~li�~��PB8VE�k� D�K6��,�ї�'W��,[�&�É�8DwIm�������b�64�:�Ѱ�G.�wq���O��-����4I!<?,O��fm)7~Q8�ϯ����=�T-,�YXǕ{���E���������{P!�a�#M�~��v͙�{�Ή�t�,���'�����󿾧����7�G�Б�u�>�����A?�d��R�O���S��T�ز�1%��/7���J1�U;T1w!=]��,M���� �=	!FL�K� K�K����d!�������FN�����K��Pg��4�v���2V?�,��8AX�? ���A�M0�T�L������k�7$�
o�%p��O�u%�i>��珬�V6_�JX��k���*Wy�A������pXS�8�����*"t �G��-�L��.5c�B,3��"q��s�T�_g��˜�T]&��HM����ϊ�R#�kf�/}I�$l����k�W�ڧq������ެ]�.F���q��F��[q��SO*�ńN�'��`��Þ�}"��惦�ӓ9���<�Nj]�b�Kg���V�㹩#�kL��cZ�A����YiUSX�����׎��<Ry��L�N�:��-\�f6�K��ybYui�C�jLf(�=���1R�A��^�E�����e/^DL �]��V�
yOI88�[���0�˘U ��(*��������ї��dN��3�(���@���jJ �.�)m�-#����E>��2���6�w���z��p��B��6Z�e��RUF�~��4Zl��z�9�V��`ar>6�kT�m��\�SHXdX�CsHR"�>�H��%�1���J�����S!�;�벂t�����N��n�V%+�je5W߫&�c�<��_#��(+3��V�~i_�F�ٖ��� ��?�/�9P!|�<{����X?F;:�_[O�P��<��^�iA�
i=�u�ve�vu�峓�3/X�T~"��p���ŏ)^�L��=�����demR���mD��~�q�5�B�>��Je�pi勠z�%�ݞ��y4G�=�Al�i#��t�Z]���mD���j��x�NP��'7+����]�N&aa@GLV(V��Rb�"�����)�6�W���\-��G]ʡ1f�i̦����Iw__x �.&���ts7T7}ov)<nl�P�ӡ[9R�N�/h�]��T6��0q�C�����j�Zm)t��i;%�_x�8f����N������j���Rw�"w�����DQ��(���=�ۡ/Z���`��c.>��}���/b��ᠵ��fܜÆ�#B}u ��%+䆏����;Moӗs��ޣܒ����dv��}]w	��-�S���` 9�:!]E!\/BS���m�m<2���if*���JA����d�K��2�͚�z�3z�!��*j�N��2�壘�$��Ӓ���Ih˼���J
Q5'4�A�����{�2xE�i�Z�����Ku�a$��V�o�+t 	'�q�!�47y���|�Cr�oL�d�d�/~;pm;�p'�'���'՜Y~�����<�X�'��҉�
�� �H��W�d��ȥi��F�~/�ic*��s�h|Cg�Sz�J:"Ң�>agn<�z_=���%SO�L!Q��W����T��HW�R9�&S2*�7O�V�-ٲs*��*偬�|���\�����)&ٻOMќ2D%@��nɧ�3�ٜ��F��̿��4�[��Axn㶋qM�~<�CX͈>���8�g�[(��
�<�A�	��T���i%�:yb�"Jq��UD�h�ەy�tD{�'�1�S�|Ǐib�K� ���;B��l��_�"5�E��e]����.�y�\�{�k��P�s�m��1lK��%8{8��{��d�xח���#�N
����ϙ!�4i��bh�.��R���I���_1b/]2H~���x`����cp�����|K+҇��a����!-���,	_�FggH-¼�
�ܜ�PE%s�'~a�u�W��U!ei����2!_4R���C:�YL���؛Qn���������4��IR|����sot�T�tnC:����1�b(��qcO�J���}.o����r,���u5�\-Ӂ})�F�.��?�-�	%i�j~C2���V�'�+��N[��F�H#q�lKN��p�sK����!7�55&��ѷ<�L[�p�^ՙH�*rt�����5A���(@�p�l���@��h�}J�M��[����.1����R�_f��U8T��pet^|X̘?wBN���%*�B���l�W�Œ�<���\jo�0C�"�τBG'�.*�Ys'_��	������*SnE{k	0q� ��3!9%Ѥ�A��<��7���E���@��{�@7Os�H *�[㔎@�d�U��G�2$�\~(��\qv����x���M��Ҹ-���J�{�:��h���E\#3Ƥ��̭���}Ͷ�Ip������w�A,7�����	��J��+�Q���WM;���-��?���#+���>#K�-	Q�kV�{���{��Q9�y��^�0~cҬ�Օlu�-��ǁ��Ƿ�c��Iy�����ocg����i����3i��"@Q��������wkU?X�fL�,� �+��V2��x�T˶!H��LT�w�h�\G=�O7�g+I'��"n��P�$�&�B�f�~X�I6��H�1��H�?
w+��S0ԔF��1�M4|>Z}ql'.Rk)c��@*m�<.�[>���60o�s�M��1U,X�w�:  Or7Öf�_֙�^�ӑ�{\'�;+Ee���W³��R�B�U ������H���$���CQ&ܽ��$���"3g�+�=RVut�ņ����C�'�D�>���̥�X
]��kR���"=C�p�8����G�[��>afK.�+ڙsLtWd�xF���@�IJ� Ȕ���h
Nׅ.,9e�u�Dv��Ei��e���_���=Ri\[�Cr���lY�w�*3�^E�oGB?�lR�+�'[��x��M�͋3����W�t����yy�(j���qkԚ=-;��Uck-�2Q�yG��>�U�c��읜K𜱇ƺ�D��*�����6畾b�ע2�Z�ԍh���6X� A(�Y��R!�q9���y1S�u�9@Ǖ5^d����<Nb��UW�0�䠳V�������'�n�i��W.� ���`\9�� N��b*�4�0wP���7y��r��^&����~X)������T��);����T���E����R*zq4DU�"@.�_aZh�1pq�bE*U�[/��>#�C.��r�&	�\7\ޝ_�ك�M"�����*�D] �a:-b���p�P�r���`ޡ���xf���^1��8iZ���<R�t;�6��v��v7Ҁ�~�[Ӱl�����c.B�D�@�r�1����Hd�U��f�����<Z��M]���U��"DJ���!�kp��#-$M
!�#����a�łA��غ����}X<:�>��&��F֤ɥ�:zٰ+�&>��EHux�I���U�n:����e�]�םɾ&� ��'V�F���8b�s����)�~߰1H���v.KB|��+�����Z��i��=�O�]�qrB��n�f"3���8��MX�F�5;eu�J����)��j,��=u^��í��I�e�N�LO2��(��#r ={it���LI��L�:�A�RC4�ϾN��V�2��#��?�2!A\Q�r��sG��D��>�}�饳y��M$@�侧2�z������U�Z)(8���|���/��K�{� +��񙢓XSU��G��}:���uVB�#]S{�cі�!���Q֜`�n�>$�ݧ��n�G� �c`�Z��s?�w-����oK�Ҭ�$��H+^t��(�G��Df�x���No�Q:��>8Cw+�h�!\uG��x�U1����{3͠pZ��ѻ[CL6}��O�
��CT��>�Ď�V�ÖP��m��b]e/A4ӿN�` Kg�/�	���q��x� `~�*��"�>�.g�3ɺ�TK�:��{��ih9���5p�*[��%��b��Ѕ�J��L��o5�)�=b���h�ʶ�u�e2�0ar�����J�%��T��򜥡ůE��k��}�b���нAP�w'b5`=2F��`�;����)J�X���O�Og�!��Y��Ƽy����	h����l�<��i#Q��Oo"n�t����S&˅k�J�#����e.�⍑P�/,'"*`�ͩB�����H�H;�����8�u�q�f�B(��Z�YCXI���zj�#/���>_�܎�'�<ɒVӓ��^N�@ TO�>7�ԇ���U�	���hً4|���������4�*R����%jl׫eI���@�W].�3� ��o:)[h� �/K'TU2�]i����j�
FR�17c:c�u[*��}ѩR':�ve�������[�q��\t�]g�&<4nc�pH�)��WNI��0����%U��R�O�wU������p���2�eo�������� �@5�?#v��H~���Q��(�(��.���mv�K/jĞ9��x��1����1�f+۷][��o��O(�쳞��׻"�	%��E�pi��U��揤\uy��ψ��������s�k}yP5��@���C�ҁ��6��f�eJcW�	�e���zk;�Pg�dG17�JM]0����I�L<i�g�^X��|'�G=�mg$%�ć!T~Rse�����QR���s�Jf\����.���Ğ?�����PpwߝT!f'?���7���w��R���PF*��/�z��V�1 �2�݊.I<���J(pЙ�L���>=�'��ȇ���tJ�C� &�%���JNΑ��t_?�}� �S�շ+���K�G�E�����}�0'_��WD�6Q[��x��A��H߹���LNbƚ�3�Q�>I��4:��YI��h��V"�N��pv'��n7Y�kUQ�+�g^%��	6����u��UՁ��������o���ǩ�)ud�'4��
�a�J�xQ�L�٪&q�Z-(�=�E2>����� |�w����wS��Y�����*�O@�h��/�#)M��m�
_��RqW���xw����d2�~Ybe�9���<+/�3����I���)1ݚc*�Н��A1ӘV�Wvn65>X���غ�h� �NK9�`0i�=KF�LR�~�L��V����d���'��V�L��$�.�d�z�J����(6)�2��1�. ;�5��m�v�ܗ~6_��R�l{���$U�)�V-��P�M��5��iH�]�,�ϒr��^�D���J��j��O�8+�H�����X%Mw�������.x�DRa�j8[�J��ښ_0x=�빦Ua�LD����a|O3)_���<�ׄK;�?kU���1�|��b�w>j��xo~�2g��(��KB�$�� ���8�|�(�eJ�Ӡzy�VE"�����o��l����L
��2w=��V]�v����Z-=�w�b@��TYTZ�_���"�%�ph�)&/�}^{����C*7��V
��
{!�W������ �g�ڈ�H/�U�����~���8�*m����\�?F�[p���7�ZĶ�k��}���;dǲ��0�ur��NtpvL%s�[����|�4��u�#���ǿ���!~��2��⊁��P?�SjY�ݑ��+s��g��&�.��B����� �$S�m�Ϡ�*]ԞmȽ�n���a>hהe��5�殅�U)���]�Ja
F0��NDu4@�.�CL��Ssl#����Tt���a�R�6���-�b�~�!(�o��H�B��GD�8�@�K��U��q��
!�',(�Ȍ�x�T+�R�"oѯk�FB���B��R�˔�q���/ꑶw�mINB
Ј���g9��d��'�,�o����Z�Y��c���_FE,��M��a���}��&� Z�^� ��CE��J?{���7���0ѫ�UX�MEH�Z�K >���%cP$-�@�)؝�;�!SpI�+[� ��E���|$(�=����9my�W�F��~�3��h�7������l�n�� ��\��U���:���P94(�,�i�5;�c;�τ� ��T���hK7�ϘƀØG�._b^�40�����7]<{k�4u"1�B�9+t�Mj4A�S�<��&+�Bֆz4�ϟ;Ac1i�L옍fX�jj`����1���Yuϩ�y묧Kk���{�oL
猭A�i��$�YÔRw��7���[��sE��9y��k�8m]N��G��ּ�cs݀+��\&?�3�Gmś��;k1���Ch&������MKiy�Ʊc�.t�~4g�6�ֽ��#yK�������{�~�(xf���I$QvXu��R���A�o>Ôej&��X�kǫ�T�4���6�l
O��_��=���/�e}9���=V��%�vX!�N�mG��,�`;L�&�w@Aw��,a��R�=���w,Ǆ��Dn4�H,.E��2�͉[Bg�BtM�?��0L�A��
��)9U�[��os��H��]�UU�:��1�;����K��X�Ϊ0���g��]#2y'��gb���,+	;�D
��݀�] f�<����e�޺V���T���u�����3��k�hw�yd���J��uuw� I+����Aq����&;���Њ�Z����)���I@,@+ >�X����l��U~U0��#Q��z�ց�&dW�uRg�8C�d
�M�3�YS,)yJ��,O)����+ٮ�u0hU�N�F}�0� )~9 �!	Z�n�:�_t�&Dk�q�q�z.~���-����x���]�(`�����)Q6!�]0����"�D[�������g	�LO%�M�d��\b.}!�4^�e�ꤓ�]�a�7VrP#�_U�ҩQ ���j�c��"���OF\Mw���W�����t;�I��V`���?��k��+g5�h���n"�������=�K*)���7!�
��w���`_!��y7P��#+�?!�O�?�����K�5d&��X�0n���º�]��'0�0,���<�be.M���I0�1֋�_H;[�2j��6�{��� z	�D��T����s�i������E5��7ڌ9"�(�a��s�_�ٶd	ve�E�أ�t��8���27���&Biz�Z�F�S�g�b^��c��[aUq�oD;�E��%	�I�5�R�9Ң�����I'Wl��q���m�ʬ��v��n���|M)�h�ze�.q7#C��2�X��B{�FB�3~�n+�rq���@�}�������t\>�����Fj�hnm��RK$j��8~���2��ׄ��%���)�FZ��2D�˿ɍ�{�w	�����$Ɖ�w�f@=��Կ��4\L��+bU]�_/	�j��>���Ez����Z��-�������p��`��?��M�B��s%�4FyY�*E�3�@�g�0N�<���B�ߩk�hh?"�k��&�������IM��aZ�Q���1EL�t,fp`>�D>���M���UXu�_��vgt���|�9��W�n�j@!�KP�-�"·�y)Èޑ�i���|�"�ݶ�ب�	���\V