��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���8}6l���މ����<W��	O=�"�Ҩ(�=ɊS�b�����㝥�5�^D�C�+]-k��i�=���IC���3�����<SO��	n�]��ؑ4g"�6x:��r945r�ҠNX��	������$y5S{�^Tj;+r&�2)to �kw��tt+��{��vO�}P�%Vz�E��˱�pkk��� Q-�8�s�
7yVO��V�!��L%֞�N�~��HK-:�=g.
�W(�2#�ߖZ0���G!�,X_Ɨ��KR��Kǫ�?��Qj�%�F�\)~P�m�)�AI{w��/i�'��!��<��35&m噭_��<�V��{<T)�9h�gљ��*F��0�n/��
��o��ɦq���LI��^��TS5'D$��>�g�d�����אvs*9��Yq�����m��dtF��'�ł�ZhX@!;[I1eX����W+kS����xʫ�C�/~��E(�j}x5�ί�	�#�S�����r9}ٔ��C@�(�~�+�$��&�ى���)u|��e ��r�-QV�.�*����̥��*����[���z���8���{�M���7�ݥՍ�~Ë	q[��r��s��󴻀5j`����aрk��/׿��F(��]�o��=t����k��� �
f�o$yL�Q���U@���?u�B�����ᑮ�?D�>pձC��ꑞ7�R�ȇ�.^82��\~X�9��E�������ݛ4s�"����ȩD<�r;?;HZ�%�툠�c�d�c\8Dn\)�	��Qh��Q���<����~%_�/�{�h=�ZH���Ԥ�Q�,�S����l.���l�g/yAwys̋7$�4�E	pQ�`����R�h��������YT�.�.�2%��ެA�=Ŧ��@!��EÉA�W:B����ؖI��Iй�;5*�i�cx�&j�D��X��ȸ��i�:�lKt�u�"Vԫ�w���7�z>�����F�L�<�161��3����XkjF">a]�4V,i`�W��n2�E����;��C,�ZaI��8�*[�=�����t�ٮD�W�u�+c�A��=.E1�
��~��i�y���a^��g�O��z�fuU��T��߮��Lz����pEZ�ѝ����(�������3�?/������Ԇxq��!�(�D��:d+�n�`
`2'�r|��ï�%٫��w�t-����,���0�F�L��{�����?�8
��9��������0pՔ0�cp2���CC ����IB\���e1�O�~+�pp�uel�!�#�G�}�Qי��Wo�ǫ���Ȕ����_jR`�i�f@n�+xʺ�.�1��+�[��B�[P�%���e�&��.�� �B�+'�^����}.~���Z{x��@�]!S�Н��i�o�^
E|��[�{9/j���`�E�G��������J�=䪦��`�[��������ꛜ�`Y- ���4ک.��ֽ�(�=��Vǈ`~@`;�%�������d�д
����1�
?۰��~�JlZ`~�����V$&�bTZ�|����Z�\���	�G����������i�t�q�~���Nʔى-�I[[�[�a�K�����3yrMy�Ԙz�	����(� ��Uq�-FE����o�f7h�m�z�rUb�B�T�и��h�Ӳ{�c^A3���g�>Vs�C�K��I�(�8b5���0���5��ת�ޤ���L��J�<�mE�U�ʸ�㞟E���휰�w*�w�87�'Řx���D�}d�@�q5d'1�v^j�Ѵt��;�����-8k�B"�*�i�e����@����a�es
�V&�^����cB@&��KW"d�z*Ǽ���� �2����8(}x�P1l�i�]�Qx4(���iB��� o�".l�)�h��p�0=�#'K b?ZkI	:��z��WkׄO*��e��3�"_�J��A{��x���7ټ�U���� �����K�H����m,"����%�e����)2z@�`��r��)~	���?�#�h���9�#�jihy���p^���?��.��*6�h�gY��b(E�_ste�}�� ��� ����ٵ��v6%�'gG�G�7tv\�h�^�NQ��u�a�ޘ�}�{�o�z����BR`� ��5>c������m�vcr������ۖ���<�9a�#qd@"��lDZ�e�稗2����X[�F�z���7�b(b���ɢ��5��)?�_�IՋ7�sJ2�����ؒW%�	���'�	���L��z� �H�c�"�+[�k�má}1E�	�	��[?l&����0-2���c'հh�CO�И����;����ٔQ�=j�tJ��کrg�>�Y0c��� S�o�;,|�r1%�=~M�����������	��p�e�[wV��Kmٙ����5�����-�@�;�}��A��<�y����^�=���tE\���џ�4x`U� k��u�ю��F;?�����%]<6�Fz��� �}*-��>%�5e��Q����i�Jcy�HR����ޗ���R�l0�ܔ��hS��XFmѱ�J��((dl�h<�1� ���8��D<h/�}ƿ;m�B"�Pa���T�e�ݭ��� ��_����iI4@{Y����+dQo	�0�a����tڵ��L����\��lN	�s&v�c�c\�N���|�7.4R��<���_L�K4们N��f��0��S��
��cpu�%����*rҹ,��j#��I�ii��ύl��Y�4S�?Q
��+s"���y5�n��G$$�%�F�U&L��ry�)�7�u����t{�*�~�ݷ+��Dv��.��J͡��i#,V��W���эb������l+���$ٻ�0�q�`.DP�[xg�)�y�{��hb�U]Mɬ�|�U�N8�g��Nʋ��(]V��ؽGf2R钰`[��e�ſ���$lO;��:����WR8�L#v�$U�a3lmtMU�O���γ��{fzL��o���g�xs5:A����ħ�� �kk��������z�X��"�� <�R�,ޒAS��|�)�2uJ�F��w�Z�3���k��'���f���#�#�.,�V��$�RX�WM]���qMWOh���u��9���4��W'e:Y��Ǟ0��6.|�C�]�w{�~��ҁ- S��Ku�p��0Ska&L���k%���2s�߆�8���Z�4c}�ɓM���{A��	��Z�� �-��_�:n�ؖ��aTRZ��my�d��v�CH<P�����
����ʝ+��
��M�J~��S"��u�Z ��%�j��ZUp��/�%�jbv̫A�Ϗ!!�aR�7�#'-i��dJe'��8����;]�B�$+G%'�>�5�Vm��Rু����m�`��lVg/�4#�p����p�t��������[�Y	���G��\$E�r�PH�g�q���A�����5氁�:���%/�h.�u���X���C���2�*���ƾ%B�J�چGi#ىc5x�Ԍ�1��(��i�̽s� !~����5��Vc�f�����p\��'E5�8�Ev�,ߣg��D^\Y�����\q�B��h(�{\&�ܕ����@џ�Ԧ?N����I�T���kXd	�n���[�`q�m�R��g�z?��NK�(�/���R)���;���\��F�,��!2�H�����º�9�����bT?N�\�0O�Y�Bj*�� '�d����-K�(k�7S�[�@�̺	2?�.3�g�h��
<�VUߔ̵�ȞF'��ʄ�f�E̺O�P��W�Ĳ������ֿk���G*y�!��K`A��~2i'���D�Ri�f]q�56�����UL��c���2�^�@d"�Ϳ��v�ǋC��\Oݿ'1t����uC���.L,E���m�6�e<ם�i��.�F�s5����u�7��	���{������Cs�s`��a��g%�5x~5rG���ۥ�=>��q8��5��PN������`Z���~5�L� La\C��zt���֬:[���o��us?�����jP���$al�v0�Tmc0U���JXf�@�ToG�����''���E���%FT�Vm�7���<�C�~W��<{��
$޵'����`zB0��&f�w�������	�7mQ��ٷ?$����^ޮ3�.�s�!["]ɽoa�F\�h��E�3�q�\k�BN&�|/����{�p���Uzb����;�8ɶꕕ�Do�0a�Φ-�D�����ʞ���u8a��4�
����>n���)�L���V���>�B��	�l�c�[�'V��v I`��L���V�燈���Y�ay|�Q��Lz�sd��s��?�E/TKT�N�8��M����r�Y̑eł��~�h�hL�U%��B��6
JZ�k� c���>�1��H�Q����ȩ�8	{4nu�r?���������{���i^���I��7�F2�x��P��xMCl�_��0Ђ�%�k�<6Ot�P�/2��S"2�Wn������=v��#�t�D{T{ۢ;�s(6�o�51k��[c�ؕ�chL�+\^i�C�{|mc�\k���q��<5=Ѵ�����lP�S����нcz���K�ù���|�F���c�X��]��f�b�;Su��&^�B��{B;��@~�vm5��RZ!�'8��b<�m@���k���xR�ܐ+:]CgǦ5�Bѭ�:����O�L�)�xG�(�Ӣ\��[&5M*�0��(bA2��i=�������zY�W5KD����Pr?	s��~��pY�xV�稳�i�5^4EO�q�|���lD˪q��~*>+�]�\LuB[zC�����uӭ��o���奎����,�,L��.:&/®�}�s؃A�A��-<�놟��h��f����x�XA*��FÑ�d�5`T� V'��!�a��I(e��scU$xn�QϷ��W����b���);��*d�ޑ?�o��Ѽ������ʽE���Q4�#ߴ=�la0oU���;�>�4Z
���W��bx=���Z\�/)���ӡ��6Q�[c�L��2�B�3H�z�PW藿�
�	60���݁Qj{5<�����[��\�`MaY��xM�!�V�c͙n<sʝe(:�aP�-�|ب��'��`4$sD�.�
����w�jMl�9�j��U�k�W�=���F����J/q�	:C9���̠�%G.��1���|��,�~v�2���E�Ԣ�!�����]C�Ֆ_�^] ��n^wT�R>d��8���g'"�5��ݒ������gQ�9ݝ6b#<�W\o����ㆈ�����L���'����^z�:'z�k7��*��,mګ�aE��u�q��R	�-���|U��r!�*>����s��c_�[��Ճ��S��L&�l�ߟ�Î6�Vǹ���ϵTY���D�M8j�O4Jd�G8��jn��ms@{�7�Q=��O��g�^���mp-�uĐ�-p���m!P�k�
x�a.k`����g���Kg�ðJ�}:Q��N�Qcjc��)A0�*Q�Z_���D��X�,�h�&k�Wg �������y�A������9�:�s�٫�377�x�оAIBl�H����2q�ӵiCW�W6F�L��B���[²��ߛ���o��܍�AB
��`��Vђ��L�)=b��Z��x1��1A��[4�.rt�4�9�x�0��� �_3�H�;��J�uv˿�`�C�$+�J�c�O8J�đ^�G�?F��c?oT�PNs��Ƹ����B&�L@E��٤g��#M�J̚�8]O��
�`����#d�~O_Pd
Ζ��Z����mRk�ޫ�Q�(��[Z��&��Bu� �� p��MfV�����^�:��
�殄~Lf�u��[���@�C�^r"e�������d����oyBn�~��1ʙ���{�r�ybR+���i��
ǟ�҂��Ҕ��E����=�/
��M�W�ӕ*jŹS_5�u=�X�o���,���)�ى����M����ɱT���~\�1�'�Do�*�8�%���4���R��<����f�zu�cwrq9���B��@� w�}�݉5����5pπ��"v�F�S���<��{���{�U���x�W�B�/+t��toɍ"ǻ��h����&,o3��������q�IHP�_|��s1�n��ꚙ���'�`%�����5��֩R|����`2�x��&�Zd��F�x���������9��K�� �^������:�A�m�I³(2^��&)<�籗��+km�)҈Ҋ~ɼ����PO�R�c`�{C!3��L!0�I���0�anMS�/��k��8��G��R���W��O�hP�lP�U ��H+Z�|�n�A�qd�����^�[�]>���;��[�O�Z�b<��CP�Zgj���/�F�!M(w��d偱��rqm����F'�UC=����Yv���(+Q"Q��-EzCRzlvF:���q4�f����uC�GԣL��v${C�']�nְF\���
^��3�Z����)��W,�Amww��Ua��Bs@���ܥa�����N�<��Aρ�FP���)��X��ɯ�r��P��T�̇�1l�I(��w)a>O��ȨY6�5����"`]. �3�3 .aΣ9>���z>�t?e'�5I��$o��*g���I���)�LF�!���`��]�=�F��g�_f���ǡ��Z^�)ܣ�&ƭͲS�T����`��B�Qrc�t������$�{�ɄR��f����ݧ��K�mҩ�?�a� ����h"�;���'�r����>�����7�f<O��C�C��~�_Y�>���L��訝E(n�M�P���o�z6H7j�8&ސZ6�`#��7���Ϩ�!{���
�s�����[ꋷ��y����L��߃����Xp�X��ᛆ��P�E��W��~�?�hᅝ�mIK�i����9����������ʥ������ �b('hϧS~���/UTX��^�ٝh����ԁ���8Q8E
�[Yn��_�`��\��ϯK�j��Mr���梽����]��h��#��Œ{Y���=�.%��JO�g�@�{�B�w�7{3;/,�Bے��a�[t�5�P	��������^2�����_�0��c���	L����:��v��&s��".F�F9li��n;lc`�/2KxY>�`�x=� �H=�c�GW���U�����������d�7�l�2o��ݔ1p6�%;�oLV��O!���Ő-d�9�!q�U+LW]q`���$�p&8�o�S�-��_��+$��4���xj�M��<��\���Y�3�X��kC3!iq��U�k�%I���,����t���F9���J��v���T8��/��HW������4�Po� ��Fz�%�'�CHW��+0\�ڎ���� ���N�Fӭ�IΝF����lA&��yu� "���a��(/!=��B��А��_�F:�`��Z�qO�B�A������y�X!_���8���ʇ�sh�*�鑽�c�<�棿� B,
Q7!'�g�Ҫ��,'�Z�\�Z#�.�QɊܐM��8�N���1^�����SI�H�&H,�o\����B�LL�0��t���cL�w\UH�"�D���p]Z��^?�R��a����+`����8g����w��^��:�J��e�x�����w:c2�?�bBƟ���r������힐_��Q��0;�C�MP����0��59�`��ӳB��� ���� r�8��xb�k�)$��٣��	��#�C��L�����1�n�R���Ł����yy��9��e*R�|N�4K���E��p��Q��M�+�ʤcs�J�H��$.5�h��k�)��qO��"r����ةE�������׋���x¸_���f�fLE�B:U�[s)^4�r2ƹ/���@\���J%��P-ͶO؞��(0��Hʕ�6-Q���n��p�[ܧe��� ���XQ� �z2�����H���☽ǩ�Ox?J����Kc�0��͝B��,3��w����������EKz��SJ�D�$n�x�6.=	��<������3���Ik>�&�vM� C�������� ��k�=�t��ш�`��hv��
T�z�K�E���Z���c/�@:���@z�F�R8�ws�¥�p����5�q^�V�Pb'�^\��y�� �cT9�P{�<�������z9�S�/� �  ���/�a���8���q�����>�ǅx`���C=��L&%~"��E.s����U�@��w�e40�ތ�ޝ�\���z-���@�����kh��ܸ��srĴk�����4�`nF��_7�c���ٜ���#�	[���� e4r���~��g��u�� ���n����EmnCEaN�_�+��mę�V��B��/ˆ���Œ��_�8�8F8�����:oe������xc8���Ick�m��n�A������l��HqS���bj�Y؀�$<���-���^�+0kYRǇ��pb�a[�Yb1���IƜ�"��m�XN��m���(����O��6��T���3�e
_��(&�3�aA�O�/�X���(�:_.f�c	�,8�۰�S}�����m�T�4��l�:ϴ������K>X�۲:��E��x�g���Hla��V�>��V1�V*���>1I6��}��C:�N�o>�-�+���DU}a�����e�5]W4o��Y{���r�1B�(�+�,��	b,�(Ki9bu=tyN��o�I�߾��@���-&R/nH�W
_G��U��
�q&d1R�r��W�b)�U�Z3�4���u��UN�~I�0��� �~ϰ�1]v"���i�����D�	�-�Ul�{�s��IM����J�ߓ�M��f�@n��إ��	E���n'�����Yʹ���ژ@#�I3����=�v�˽+�1,a>��,s�ƓW���-�yY�9E ��u0E:�'�na�����+eY>��&�2�����d� Of]hqEAyDp��aBx'4��d���o,9K�&qF��jV�]�&k�<S7*9:���p�㐷���9!D�i	<�&�8&�Aێ ��R���m.8u�������1��o[��@A9P
̆�w�t��s��{}��v��>4�T#�a�a��t�"k�����sE�|_y�TC�@Ui!P�6#�u'���	]��7ƨ�܍���^�Pv��ݒ��tϝ�S���Rh��Ql���e��B��4�u"���^��t.�J�`[�Ӭ�G�{�l�l�u}�`~ɺ��+�T<���X6��I��?�����.K�`�<����#��p��H$�%nxJ����ؐ ����T�y0�t�����Ppa�E�`�9��ڌX�z)�x%�Z#��W�9�h�?�d:.8e�bW�&� ���\Kc׶�ǝ��3O��I5o@#��k�7���5Rm,$_XlT~�g�&3�$�PY���H�J@6�ޝ�z��u�y����/��R�x"i�Tox�w��+�G���ف�6���:��H�t�i�V�&��;�;�5Aw�@��>�2����#c�	���PC!P�7ҁ%��Óe�4A �[le6"�v��(�i��aW^ M�����0���ش �M8������a�{���i����ω@�'��VD�g�+�D���l.���$��h��� B����9�!���C�Z�w���g��wwc
��XG�Hz)=�
���RC�.�zK��u�P.3�c��0�ZiՇ�\�ٖ�|,�X�Q��"w{:�:���@���+~q񕃈䝬�g�B�W>
����$���{hf�aU+)k��!r!v���������^���e�z0�g_��}���j\r�\���:��?QT�ӵzG՟J�?Ӆ���_YЁӔC�N��}�ȓ'n��9�E�����dE!9�8���e�c�1?���(G�,�R������)Q�7d�܆ǔ�ϩ"��N�,y3*;�0U)Եzs�B++ ���K�C1�h�'R۸�:�ə���w�������e8o��O��'��[��>�1��~��'��~P�;T%�0���P��rz��8-�R�h�T�*ă�B8��v�8�&6,�R�A�Qďjw�1� q���*���a�������N���c
���#�vJf�@�Cym
��
�q�0�����:���lW��;8�cxu��@8�e��a��c��F?#�g�z�k>.L�X].9mw}���r�����`��e4�.w�dql�ۦC���F�Z3���R$ ��)Τ��Sz����.~����Y6�R̖�S5�k�_�
�t��=!9�sZ�ޜ[3�4����$��B���������x��p����	�ݠ/C�H������,�����3sz�.��t�w{���|�)ʵ��,#<<0��m� �sI�l�{�p��|yWa� ^/��˭b�������#�9h��`�1��S��0�\�O�]=*�~������Gqer�|SW�	��1���;��~�	���yﾩ�_2�C��Oﲛ�z��~s�������$�-[�L��d�o�اq:X=��9a�ܕ��Z�	dU�`8(m��9�YF�@�y!�Pg��������jezϳ�[[;�9��? �7������>��u�$>_M�1�!d�}�Q)IW���oޮ��L,ړXNI��0nJr<̵֝�F���`�O2u@�ܰ7�#����Gq9��5?�Vx�'D��O�|@���u��������t2���O������-�=�E�%�e~i�;O%��	Z(�����&X]���J���{�R�>ĕ(�Y�+��Nh��QD�T��az:\�����ή�X� 1���f�9��Є�|�S���7GiG�9ö�� ��̰�V3�H
,&�gr�VD�b�A�ĚHNX����(��k��Z��>������{�F;bv�7��g�d�}c���Q��T��(��D˥�"���A�o�JE��f�|�RZJ��֫��4+be�[��� �=�<�hEk����Ɉ�/��{y�-*(�^�l�����
��6�^�iۓn'B���=�#�?[�ϼ��ǆ\��w�5z���"vJ���0��
��/~EK����	;b$*ge��n�j�ڏ�U�~�71V:�[m-� �������⩝�.���"��*�F����y\��`,��Ӻ��&"�/@�����c���S�+�MP+�����o���eޅXS����5Q7Q�V�쑛��T�5?���1柜7l�vű5�B=��mf�t�#s�@3�$�W6cvzwNc1���u��\mէ8C�"b��37Q�+@����.J"@N��*�pj?$~��R�I�;�'>���g�(J?"^D���)%`Ӂ�۪�v��$a|��5Ę[Ѷ���b�\n2���i$�t��I���	�'�o\��7�x
n�L�f��.YC�;�_���Z�"��_ ��+^��`�n�+�������_߷/��I���6�f��
��5�A��G�f b�ӱn�I�;�vgN�t�b�/�l�xX�o�oA#�����3�-���K�`"m7ZFq�)�[1 ���,v�Pa��5o�ށ���3j�n��|5�仁YS����I�b���z�`?&�Oٲ}���xАCJ�r�}��<���ǣwoq���)]�r��7kF�h�o��c��ё)��e���kM�Q
T'Y26�R	�@Į_%��v�f�Q�T����1�����5+^k`%���B#f�m`�Qm�m�8�`4*��\e>5�y��(��EgG���V��Q���3'H��:<����]("����8T���4�L��B��1a7���i��;�7>=W5Ӟ� ���J9sG?sZ�&��ʡX�4���.�XV�_���,�W�
@L�M?��A�����
3$Pwf�YB~;cڡ����Zg�����6G�I�~�!�=���&�?k��-�T��j+f�h1�8�7@>{��"��j#=�e���#ˍ��yU���1Kd
����;��ȵ���D�M��"W>�Ï���Xˏ�+��:�-R�O.O�a�<����r�٘�Y�$�����t9�/��_3��6�e@�~����Hc�MmW�!E�b�X%Ņ�6�{^<�~ۈq�qȌd�됊�v��z��< ���@�]�j���94�}i|���L,�dF�_�c$*�/_5W�}u�C��	e%M}�1!�-ȼQ��Mʐ�v��}"����W��<��V+��{��w�9MSt��AK�T�o��>�[*	S�pʍ7qM��lԁ�\��� ���I�+ޥ���[����xGȱ��4A����P�������Ҵ�����2!��%(�Ow�`��e8*~�������À��<�M|,�"�ٹu���3$/�9�DU��Ҷ)��n���-�j�����������6����rSy����m���?ᆸ�V��?9���-� ���Zm0� a3�i�qc�=�(����\�wT��C �����dY� MlK#A~B����n}���U��|
r�����V�o���+�pF7-�*�|Z"������ZM�]F��(9�g�kH���0@�BS��e1��2t8�����l���U����g]� (�%ݜ©��m�B/6���/��d�6�o��9�|^_�P�M&��\灁�"�*lʀ0��պ3�r�� ]r���ױ޵�^����"7u��=嗺�W��{T�o�j���� ��g8�o�o0X�N,���#�I�in��M����<5^��B�0��X���P���TZ�#�Z�v�m��`r�7ʇ��Pl��2(.W$�I!�	^(~	���b���)S៺v�L��咨�&w��"���QW�)fA�"*��˸搦��gTG���dܩw�.�`��d�C��Ly���N��L��x��铗^8SK�X
�m���J�X*��Zk�^l��b��~L�!�<m�w��X/e|Ol�>��'z5�-Y��.���r�e]�c�ԩ��
��s'�%����G�����1
[��c�v��5X�ifۻG�r�r't��rT����6�j-U�yI��M���A�~�8���D��F�-������u���B�~Uþ@��>�·V��/��ȸꪳ(���
`�I�d�d��eBǔ������d�wc)��޻���x�FaS]�SP5����`a�.�aW:�� �G�s �j!���q�[U�M)�?�W��B-Q��1(i�HuSC�~� ��?��v�w��[�頷W�߿g �\�yǥ��	�S�M-�	_����������=�P6⼁��]�Y�L�Iv�m�q�Y� ���\�PAj����:�s�[0ǍEb�����$MܔxMh��ʺ*������	!{���2����^��y?s)�V̨��V���8s�a�m6�{�o�*wΛ_zIS�����0��7gJ��Cd�O��*��w�;=:I=K\�;KR�D�������Ƴ��$��|��RO���[6�c's��b'!N!�~z���VS�</�OI����UZÛ-�'��r���h�{\]ޜ1z���2��v� $�ઍV�c��G� ��ａ5d��wY`���K�L�Of��Vg�$5H��&l`ivh �`�=fa��<��C�׸������CW5�N�c�c^3���Y��o��"��Ɗ���u���?H�X�C\O��h����0̜����~$��dAhe�"sMz��U_-��=���|��+4��̂�崿�ƾ��S�i�vÒO>�iZBϪ�kJ]��q/��oǘ�@��:\��^�8Q���Ǔ@��3�����T��ije�B���S�ٟH>��_�۳A�O��i]^����Q��2�VJ��=��S�S���x�|�X�������@O�|�JM:_fm� ~�1e]|��1�|��
X���]�&j�u��~DΥ�q6���m�{�6g����BQ�0;�N��	L�o���<�T��M���r�k���u�K�-�nrs�
��%b��E̯y+8b�$Q���+��!<w��eOQ��S����ݍԴ��:�+�����4\�{���P_s�-p~�=V�/��?�_��h���7�8��S^��P�d>R��'�*_Y��'�ܚ��-�ނd0lS]�j��Dr��W�Ɓ��q�L~�����1����N��#�V��dٓ|�`�+��8��u��T�c�V�����.f8���_��tH2�����O�����K U����Y�OH�.�>�1��xj�Y����
4E\}�n���?` �Z�D������g���Ϻz|�H)���a����YU<��*V;�)W U� P�H�a���^B��K��i����#à���	:�5�s��>���Zp��vG�;�T��.�.��z�.7Uy㲃��u�E��j���gP<}���(Z,j,~Ԭ�r�>�y��dF��kf���<�� '[N���k-hF7�6X�&�]F��A%��*���0�M�d�u�H@�g�M�ۿi��IC�W�6J����Ũs-���	|o��R��D^zm<�r��evĮ12�p����B��ʵ�u�����eH��Y�Q���k���>�(�/�&Zbt�V�O�+??#�)�Y�".�x��j�C��s�С��m�1�#�)�A�	�����Bb�M#{{v���1rq��U��{.�݇՝��	;�&l-���8s�T>�c��!��i��rf��r������:���5�~3�~�`y��3%C������#w��7��F^N[k��t�ųq������	`B2�Շ'K7��E�	�#����jϔ�q�>fP����U�=li����%)Ϊ�}t�u�G��F�Յk�N�^�QlM�c0P����?ޞ?d��}�w۹�!3E�'#p�we9h�q����k-���PC5���Q>��
ݩ��eq��˵��62rGZ�d�����G���b.	��)�_�Ή�1�t*�DS&�@�����oI��L%��":���QE��,��A��z�+��#	{������ ����h	����}&��?�C�䗷�O�w;����I7�/o���n�1B�/�qLv����y�� �0+��\�T����@�n[�}����zT�y�y�"�|�3� �
"�^x�������xP8��o���2K��\�@�l)�|H[i\�lP{@��js��}T�B+[�c9��Ȍ��GS�������,Ҷ��mZ�i��t\�#vA�8ނ<���6�N-h	�y�"�&��:��ӡ��ĕ��XqA�*�B�tT2q�us�x����Vd�����K�Ѿp`w������B�(�7�ld�J��������j)�`�ٳ��6��%��-*�i�e(�KX������.�j�� �a+�Qb�����\J�)v�����E���f�H��b�G�
�����G��^�I�J�z�m�c��������ϖhc�/���Aŗ��Ҝ�
(T��1��`��OC>H[z���9��C�.��w�M3��p����0~+	����� Ebt���>�L���*�閱��Ip�B�:�7Q����z�� WXi������u�̞��!騄��dIa)�HY�=�r}������,��'��:`�OP1���{ߺ��΍D(��m���{]wQ"��2N+gP��
���s�v�\��>]Կ�C�	f�R�IT�GkP�Y�`�ێ�#���C�]��r�WE����<�*��B@ 5B{ Y�������r(%�;V�;�hC��D��v�ޗ��)�s������j��#��G)���
_=�N�U�?�'�'a���o�uD��c�kў�:<���p������Wة�V���$���!}��Aj�q��K��h�a:G����lX�ٷY,*2Sf�<PF̌5�t�Ċ�υp&����� Pk���9L~�Àe���M�7�0�yRM�
ýDB.L#��9�$(K�������*�ª�P����B�M٥>{U��(8��NZ�����V�R$��@4��6���i�sy�ΖmY4�M0yU���<�S�z �(�L��ܦ7�U~�C�h7p>�W��B"�/����D��W���49�Z���d[�^GV\��7����h}8����t�&@��о�r��6����,l�r��F>kW��VI���J�ή�h�� S!�@:=�v$&)9�35�,��������+�B�P��M�̞H�p��U�.��iҿ|e�q*�۹$P�r�7D��p����.C�ߪ ߨٟ��44�Cd�7��^��q�2�UԺ5����tv9jp���m�K�#����/R,?�۹	�d��a�x/%�w�/�+i�P�=rY]��A�eu�uW�$#�$�7�4�M���4ĕЋ(t.�(�'�5�^��H�б�7M���/���-�zz��n7]u.��e*�
�?�V���:���	w���gTfRl9�BJ4�.G�*@*,�#������c���uЫ�ZA/���㽕�����6J�'k�ޕQ��t�РT����t�8]3>���¢��sT����M�〩�A݄X�C�x@rt�N-9\a?�I3�/A�FZ��%	KD��T	���zf�戭O�����#}��܋s���
���hS�Krj��߂�9l�5���@ũ�*D��fخ79�u���-�����)�Ʋl�L[�[�4n���~ue�j���4{�T�(���.}m�s�� ���l|E�!:��~)�0e�o+�����x1�fw�u�<���x��O٤��((�K����,������ٸ�<2$h��Kv��gћ�X���y_B���O�˧�l��.�����V���=7�����;�FD�D�P�<����z�e��h�ݑS�Y�r?+53�9sJ���G��{B�V�W�@{�IdŤ�?T�ٯZ�	o7_.��r�x�sl]�V�5u3MS.G_m���ʷt��X��n�h\��w�{qJ�j��Nc�x�;�f[���Ì���t��V`P�z����"vW��A��$L�T|El�W��9CfPBToI�Lx�܏�f���g{��=Q3�̫�q��[��<D����֮��3�G^�O���{��Ƕ��-L�n)�	ܐ��M�����O���ALJi��j6�D����.�˫�R&xp�0)��ģ1R4�FN5@�wn�a
�=6^�7:��:m��\Q�	2�(�.��}�����*Ԛo���_�@7E��i�k����ZZ��@dN��_pio�097J4���Z:��^QG&C��Г�1[��jO1�����]Dh�[٢��أD1�)0��ASѺK\lz}���;�*+���Gs<�����"�A�]aC��L�:�(F@�'0EX�qy�*�S1ɑI�����Az��8/`n�4d��,�f���8?\J:��͝�_����=h􆂏̗�kIp�P��61�
5������L\m���:g1�Z#$t"��^͹�}����s7	7d�F��t�e� z�C�72�$!#�9��H6�P��N�E��Z>�DS#N.o�c��pbGFt��B)���P�oQ��x|L�~!�q��kæb1�>S.���w���y�D�~+�M)1��(1 U녣�}��QF.�k�룩i�v�?�zv��Ѵ��;��Q�,� ���~E�:��k���i�7�Ӝ��P�����P�x�Z䱮�:�"g�b��jYvrLU��;N�?�x�V��H]���+d�=!����Y0LS�E��&���y�����P�uĦt�dW�rk.s�w	/ԫU{k�H��v��Q@ˈ�_>���Ř� J�޽�8N^��B�@����q�M�G���2J�DQ2��.{�Q��u�gտ���_��1[��Ϲ'�����g-_&�#A����2iMu!���5{3���Bt礉\f ���/�1>gZF1g��N�d~����%��4��S�b|[�<w�m����PrTL޻;�r�ov�Z_=a_ﰵ<����֍/�{ʼ���^ZF>A3�C��������