��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]Zɬf(�'4�o^d5��o5�V+�����YE�٘tv~ұNVz��!#I�PWa���T!fj�T�(�Q�P�=�׭�[W������L�9��0E�K�M����C�N���K��N+����@9��x��ѠB��yPI�v���#l� ���F���aK�:���$l���X�2O^�lhp�F��������O��uY�guI�$�T]B�M�Y]�,�<��:yہ��4T���=�?�P��k*\��)�M��D�0t�� uI{F�2]w���S98�;�V���O$�&Sq�Lr�eQ��X@�"��F*�`����>x��o�mJ�2^#�zO
�z��_>���x8�+�����RhZ��[�pm�Ғ�`{ ��t�T{��ڿ���k}�0�LB���[]��	���?׈�h��\Ji�'�}�{�ϭ�3~I�9Q�>��Ї����z�	�μWtʟ��d�GN�B�w
��94[&k�'g��S^�����.�����
xO����x=c���HG��*4��"�qs�\K�{�^p��qV�wh����|�Z��a�U�C��pUOi�~�`yM�pŬ�J/ly�E���ԥ��N0��0�J+���X,��[�L���|�#[��Vp��l�,��������@��p�S�̡����pd�}N�: ��K�㳯��TT��Fa)�ܤ[����n��b�V-�P��a���M��1xۗ�=���O#]M�$n�I�|��s�쇈�ȳ����O�4#g�����˵]͵O�B����"�r��%����El��k��LS;��0I؈��ƂZ�r?�3���-�or���0��[C�4��Y ��9����/d�k�� ?S��z�ț��qZ?�ṯi���R,��r��D�"t ~�9��� 617GW�E��hXq�Uy�=���us)�O���N��w����l6!�R�RA9liz�K�`��b��pX����������g��i{����|�:P��/�1j���ROlhrRoY|{b�����>�1�	�6R��J|i! �h�G�ř\~�z�ja/ ޹�߅�[C��3F�D���5{P��t��AG�ִ�A���<��`����\	16i��c�$jA[K����o���x��w��ʝ�M��'w�ֿ��������L^�E�8��)���"8��-�J1^�p��{���'w;�A�t0L�x�.32�o�s��ח��I���k{�%�:!�1������x�}�9���l6�= �f�ā�.Ǡ�������$_p�5�Z${�v|�g��3��.cԄZ�N
���d�m����0��O�<����	��=�e`�$�93�S�z�iB�=�M��� z�9r�V��>���y�(Q�������%f��3�њ�:V��NZ������3��*�^����]�����V��*d��8-�-��8Vٺ�U|������?ֵn_]�kA&�,��k�$�&gtYU-(�J8�[*�F^�FET(��S}C�����#���LE �����k���W%��Au�٣Od�SVFv�R���י<�C�x�y�5+�����KU�bT-�_f���0M�wE��i֫d�Q�y��Mx$�>�Z���.f.�(g��=d�l�R�#�k#�uW �U�A�sY���k� 7����;x�Ƨ~�Bڣ눴����]���=�d}j��{i\E�WK�z��`�W�.��YE]�u��ϭ4�:ܞ��I����ًm����%4I����墬 '�T`�h�tM2u�\�־�����^'�`צ����h���� �U���(@�y��<.O|;�Z�x�
��:�vw����2;۫|x޷��W��%-迒��4o����Ų����۽��-���bT!FP�F$�[[o/�kj<|�h�q�;��_��eJ3�o��]���A�9��3q���M�n�tLt3�j��)28�#2�':�][�����:�%��]��(0�n�);��U<?�_��Zҳ�qŋ�h'�b� H���Ȕ9�����C�Ʈ_t�[����l<4C�K����겴�|;K����Q5B�l�^hZ܊��x/�\��)|�gt$��S~�Z��Z�+����sB�u*|��ب�bJ��M���,�^��'����"(F|�ۉ/����� ���q މ��>BHH`)���,|���ׂ'�� c`���O�Zֳ�!F1� ��+�?Bt/����ƈ�&�CqcЗ�'a״���x\Mԝ��F��",,Z��s	�
6���� |�[_p&䀹��b�-"�!+`�~L8��.<��������\�T�Pk$�۟i�U�_�}m��Oοr��:>0K��va��96|=~�g#�lͶX��/@��g�7�h�Yp�ǟ,KE����u���v�����^D��>1{�e�S�1�FfpRc3S}?L�eN"K�m6)lH�aϦP�1cy`�g!	�d���������4��N>�[�4��r�B�|^��R�+���щ�lBI�6W?=g!�)"NR�V�sA�6&�u���]5V��(1�U2���\q�� ��J�+�z}�˘%9���ͯ��G���Y����Xg������>s���k�FKLY԰���!�DP��C�5	��w�m�+���W簠�6Z��0�0�c��z0ҿ��(�u�v��f�@��US��`=sO�$�a�.`R"�����q�s]S�ή��8������1�%�����8�N$���.���Й�7�96Y=v�"} .�!��Gΐ�ٙx8Z����W�?�5߰u
��qV���cH���B�ϫR�ξ{��4�hhn�e�@��>�3���_��[�X�j��C-{��NҶ����~N��h�j���)�V�:1J�s7�_D ��+�'23Xχ��t�pA���?��0|�l~4�+XR��Xs.]�k�7�H��
�N�bJ5F���9���������b�������2�w��(��_�nO�=��dP?C�|r���VAK����dtU��~n �C����:t(|5U֪E� ����L�������^W:qP=~���{��_vA����hJԣ���;��~ie�/�֍��1�M롸����J{�	�K�+|�;�=�鷼�������`<���Wx�sb�����e�� �<g���O�����Hr��z3ױ�=��6��8��45Y�`�cZ����0Q���%cm��Z�>#