��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���1���"ء�o�*�w�rR�Ɨ��c��#�����1t�U)��u�'x�Н��3���X7Eէ�±	�E����u��~?V_��C(<+>[qH�g�'����l�&6 /׾�� ��C���>�K�%+tݗ&y�	&���W'[��5�����f^4I��4�R6��J��s,M�Zr��"?�����a^���?j����&0�:�bF9��
�)�k��w�o7��2����g�b�!Q�k}N����2+/]����@���h3��9>�<7S�Q��<�T��A�
�#��ݛ>o����3K�$�d¢��A_���E2�=!X�#�G7�=��06�De�fvӿ�oԹRj��?Y�0a}X����� ��itN~b���K��2Z���d�[o]�����`4#4,y�95�����~-���^��݇{�e:«����<5�Jǂ5
<m��P�`��c��5�삱E��>�Rˆ���w��D�	W� ��ˇ��Ө�6`��?#��Y��X6� w���;S��`(��l����T����G �+L��`9����ji�'�Z��?YG���A\ �5ܳSo�,pDd"ÿ"����Mַ:3wa;�_��b䳉�$g;��]��9��h��7��b���T֊P1���[�|���<�J����h�H`�,,?c�9]}�l�ʛ�@WN�)� jGL�n��d��cK�*�.���8x*�������5i���[.@Su�o�fq�~����Xf,�f�\���Z���:��j���0v��t���/b>R/�����ݖqe�6
G����"��;�rݫ��U��Uq=�hp_�4|� s+d�,���LB�2��;`�)(pu�|M�n�B+]�j����2�tHy2����4���Z���NϘ&���U3��W*�������	� xn[������/�F�텪�y�КI{Y�g=x��!%����~=O�-�Γ8�s�A�i<;T�  ��wyrA�7�)�D��\�Ϧn�Ӧ�_6��o�PBl�k1���9=1�
�d�����JY�G�W��Ub1�Z�7��-�E��Hj���塺�	4A�^�E;)����@݊�B/zH�0sKX5-�N8����;_-�����6b�@t|�q����E�F,�¯Ȱ���9ż�( �88\=���+���Ӣ���<;���M�!��@�����oa�/�Q����Y�xo!�[�Q�$i*.V1��j��"K�v���x��B�u3�b����L������A1z��LQ[(� 6��V����q��"�@�ʘ�p��
�z��-�����xN�h���&��P����G��=�{
��)����!���v�&�yo}�S��ذ��]�rZ�L��
��:�T����i-K|���^Q���}���E}�!�3�/Uh��"��퓝e�˝��Ůcm6;`�Gh�u����ۺ=ԛ3,5�_��Z���Fs���,_