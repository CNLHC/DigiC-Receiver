��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��M�ۯ*)��k;L4�u6�oErK%��;��A/�������)�j2�j�&��Ukr�w/������>�hנ,H/�X�X
`���s��"���(�bAfϡ���x;x� #.��qT��T�zw��ߏ���.N�O&�	��+�a���+�7X��f�Ʈ(='~���VBU�s��ҩ�K-�����<�[�0���`=xhx���Ɓ�w�'KR��X������B����o����}��~�8hm�\��%̲�����O���bK��Z�,�鏥m�^I��y������?}��R�F|1��&9�3�7*��vGp���R|rY�$0�>�J2PA�~Ï���?�j��Ob���;��m5ñ�&�e��g����m�2\<�3�R�u��Y׌��76�NJ�]�>Y��k�w����H�B���m&�Z�_ŸdI}>��yOwj�%���3�Wx[	���t(�d �F������X��_�^�����{1M9B���|"�����A��CฦT
�;��X
 O Sw���$��Y�m�}���</���y_����I*M@��^3h��^���͟z��u�ф�j
�Ð����M4
�?2x�s�@J�Vdք�\���O ��:nW=���GJ��#tQY�`kfٝ�؝?c�4w��%��I�A(De����f�������H��L
���Na�P�>�E �����
S�b�T��x�W�}\�ҀDT�@g�����۪��|�n�{�"6)a�f?	�dskq��Ŗ���?�4m��t\���\��NK��t��V����rCGSj��T<wX4��#>����H��?LZ{}oN��!�Lo��ǩ�䘺�SF^fFFd���U���K%�/��Goҙ� 9�o��������ƨV�������M[��^�d~��C^��`���t��R�t�Iy�AMt����F��t�乷�Cn/8��َ��Ӟ��m�
�:b�Tp���I�jMBfPD�%��Z�I��M0gWV����L���E
Uڡӣ����fV*�Ha���d";Xԧ"�8��ͽ�4b�vq?�5^9@�vp���J'�Ǖ�G	/�zܛZ��X��H_��	2�4 �׫�FcF2382�u�^v|/�\x\��l�S#�6y0��s!���I��7�+�mA`z���ӝ�z:�9�\����~�V6��!�{�m�M��]^�F������~�-Q�w�&G�/ ��N<�X�Ĵ��]U:�e����Ѿ*��k�≷�Uk��N�7�H�'��u �Sg>�x*��j�]�#���j���l��T8|�p�a���ƙi�!p�{KY��޲����G�=�^�o�()�	���|�[�+��7�)��b�����ū���$�lٓ�#Sw�G�x'Д=���H)�;���32y"[�Ʈ�X%
�rX�?֫V�F��$5�NI��^+)�4�(�g��,�ht���4,:���+�x�e�
�9[FR'�8�DՕȞbI�1���)�~�]0q�L�}�k�:dʤ]׃y��Gm��I��^&ˇ���E�Q+��;���.f�#�_ezqWg}/�J�S��=��]W��'����P�:ŭĒ�r�k�;�(K��l9��T͙HҌ����g�4ǬB����B��[f�]��?�U=��Ai�T�o�d�7F;���:��Z�K�7y��6Ft%R��q�89�N��H�D[���7��z'ږxv���������ȍ��� �!-�c&��52=�`B�ИA��D立�`�T����5V���Å�R�'�H���`���jp��d����Oj^�S�ޮ��ɳ���	
̿ӓ�7m7꽜� p�N�JgT���E]>?{Gk���[���^��j[+m�$5_
�) v1h���;���3�<��A6zG$����M�äWag[7����=�xXw'�0�{�	�2R�[w�t��1,Co�	=�#l��c�ϑ�"����9�s�)�?~���5�4�C%壅f;^2�1�b����br@ɶ�Fu��n{���CJ�
X8���P�<�s�����]�D
��V��u//9A;򾃗de^
����L�xo���MP �Y�0Ō�YQ�e�_A��A���C&���*������L�-�}��sq�_��l�J8���=���Ôe�sn�W�w�QG���5�����If������7�\��}���s,I�@����ޖi���(,����Bs>�k�kK��>��R��}�>(����z�i�ܡ������@v������$��Z�´-���m�x�Rt���E�-�C�!Ic	�2����FbQw�C�s��MIDD8�WU���_��9�{�X�eѿ@��x��m�H����7Uߠ���}��y��~�C;��tJ6.$��Y�ҰK��M>�X���+��Pƒ� �}O`A�=!�
λ���^P6]�F�"�+!?E>
U-�Jgl�q�e$w&u���@��̩����n$��qgs/�|�㝉*�	S���� ���<��X�{�[m+�+5ʚ����W`x$�~h(��X��W��g�tewD�����@�Y莭u�,k��b �C�	b̹n��(x7nKWF�ڊH��M��Ԯ�A���$򈌑̄F)>Ѷbȶ��=6��V�y]�WԬ�m�[���<u�$��2
pT1f*��lLf�<�C��������;[r2O��49ݝI�<�p��2.l�R��zM��7}� C� ���b��(S��*u�:
]1M5�9]�
����:~���58�U(��ֈ?������y�{CT�Oƹ!u1�*9a;xD���p��uչ��r�7���t͝��]bz� d���zG�nhH(�藯%ɦ�>��C#;Gd!et�����#�ꝹIЃ���#N~���������|��ⱊ�M@Y�n噂�C4�c���'���δ71fɓp��/���Gv��ݖ����W��b�X�[Y��^�4[�-��
2u�j�`�|C�q�Œ:h�-�ZC.Ps��P^�'bD��#�Yb���q݄;2F���D�CdN�qKi��qK�A��%��zm/�	����zı�!S���#���U�=p��I����s��x+�#(	(��s��ݵ�z "�~�v�w����f�,텪4�8��L��P�j��T˲q}(��P�'�7S�?�̀��{�{t��ş�%�9<VU�,���o�����R�Mbc�2�������M��\�����NQ�Cd)������Pya�B�j�or����z�%�0�W��,'��V�'!��t:2��{�0S�d�Ri&�����D8�B}��Ÿ�����Գc�>)|��M._�9�Po�OY0K�w�8"���+��#�̢d�KT��w�?j{�iZ�*+�IjS�]��B:R�u��"1-
����}X�?�tﾉ#��j���%bT����j5�Jf�2rB�wq6xag������O�����*/(`�n�i�����H
�k�PE.��ne@W�Q�qCyAl��7�Jdw:�\��n�x�b���	i��X���6ۻQqq�d�Kf��y���-�,�o��xl���\3�VO���Q4A��^�sE�pH���G�i�x��q���lr��v�e�D���m����]��6q��Lcۦ���=�j��z�E	� ٫�Ll����0�aR�o�5\o`hFo�šN[p��d&�S��NvT�<����gS)�;��À6_��:���G�~�$ǵL���3T;S����5�H���yfZ�.�}I�*p�n5�����������j|�By �V��)�{wGU�O��o&�Vd��P抟�>�@�)�\T�ZLF)œHY�á˽���팟�;JZ�FKE�R�{���	���$@���}@2�Q�
��.I��ʎ�+�)�l�Qc�����k����=�*Ծ&[�lB���=D �"S�.�oՀɢ�;�D,�f�Y�
KW���&,ٱ�X�@����_IC��9~/�}��(l���|��F�|x�uʯv��L�AH�w���4³ϫ[b��7ab7��*1w�`rIm/뾾SA/�g!�,tJ��S�`#�Z�j�~���`��lK��5GJ�z��6e�)Y�����6��WmZ]�ޡ������-�����9z� ޥ�ݭ�no���u����B2�׮8#+(K�nϧ�R�uo;ثe#_=^�(Wy
X�aIv��N���& ��5 bc��\k��j����_�_�QZx}Q��Vh�SM�s�`B�`��X��/���=9s�礰������c��ˤi�R�MD�{��t�W�d�K�Cms1�H��i@4`�_'��Y��@���{��^/$��' 39L&՗�Ɵn�H�'4 $J �����Q;r����|�Y��7���9�w3�hk<��6&��%D�S��Ɂ�ZO���k��1��C���_�R-վ	�]�X3h�~"8�/؍���	���[�g��ͻ�5U�[�WU��9b7N��:^��cps�Q��]�G<,O9��c�z�#n^�x(KutcK$x���ލ���:ȭ{#䀹\�����a�mWmrH��!N2���73���n�I�~�Fs���/S�t���k���U`�Y�˾*���6�vIΤ+N��8�`y��}�J@)w��׹���&1�\��>��	��˿��\�q�����(�X������u�,w7�ɴ�A@}��{��g�Q��pޥ�wy묿.�f�g7�\����	�]���TV��i?!My�n����I��T�n�NKUO1�#��� �C��G��`w��Bސ�TC�v�_փ�&���p�V�0�/p�j� K��TM�)��U��O�;��q�.�Z��A�6�qdrg��ҏ߹cW��E��pg���9��9<�B�*OV�t�N�}�'�2y�P�,ݡk�����/S�&HCN\��,�x�Y���`tOq�jF{�g	E~��顉m�H��F#�E��7zR{���y�WÇڧҀ������fsF(\#V�k�c�:� ����%0�����F4fɯ�G���4-~�֔:+���x?��;�G��y�U�=��d��`bU򝡇[S%���@e\����0���b��x�w=_	�N6(I�>���,?~Ľ=�&>��<���GI�0��p��}�a���"��;���˧;�Z��^_��ʿ����M�z� ����!����De:� n�}{?�
��Q�M7̛��+���C��7\�k���O�u�@O6hv�L�4�ZP�Q��c�	X�Șh�̀b��s�	-h�%�1�f�o��P��K)�R>Y'���9ô�0Rm�Ŋ`6�U�;$i��R�9s�"���zn�ڴ�{@1o����f`va�sB�K׭ɘP��W��W1����2t��:���Z����ڬ6S�C���L!K���RBnie��3����@H�*nM��l���W]��ZmQ_c�wo�A'��\�K���������}�8�E4�D'��rO�5LC:xO#"DF�rU�ݗ��L\I�}�����D��k��U��թ.�zK�s�����d����YC�_��IN}��MG7��NV�iI4��iF|%Bb⥓��梁��m�)+kZ���+���R�RM�|��3�\}^��5�=�t�e��w�ã���7x!�wyJ�����Dj��v��D\�{L�$��@�p_߿�}G����.9��i��a���%�a̭|��V�;)�ꇻ�F��:t�`Af'3���A�ڐA��Ė�yP��γ��9-#�D]q1�[�S\��9�"����\U����k�������T��ˠqO�6`��^�����̓�Q^�����c}�4fNo�͓�8l�,~�3�/C����TM�x���Z`(����[���o6��6,��!8; oyw�;_�~W��.�����8���_��8k+��6V\0n6z�7j6��>g<>e@R��0U������ ��%p���œwGS�����v�B��Ե�f� |��!-�)l��K�[�a}�F��:��[�޻J:a�M��HꀸG��jC ��ż�Gc>�j+^?�W���IrK�?�!z	W����0���9r!c�@<��Y��2�J��	�E�G{��ќ��֓'�����k�uZ8�~	��.�Q�Y��;R�bޕk��F�r�S�)��V8 �<�2�#"C��Oɭ�a�fFO�N.�i~ݼ P�򎒎����t�R.0��m"�
\�΅о
�����s2�W�����b��yw�焋|h�:�V���qK?W�2p�#WZePU�W����ڢ�:G,ꁟԪn���d8 4��2g�:����L�w~� 	����><SO3��|(�� ����S�� ���?���UL�I��Z�5O�S� ��ѧՌ�QAx�>�ˌR�΃��Ș7`z�M��d;�ⰲ�J�J��w-DHf�c�]�w#ƧN�>�?x�/ ��'H�f3S�=���:�V9jf1����ڞzGFY4�BY�m��Zq�X�,�r�ƅC_¤�v�O�rV�AZe(�bb�OR��J3<�N��K�Be��{Íw����qEJ<���\�:�oZ��=8Ͻ��A������Ə%�Fr�O�J84Z-8�bUDѯ7��z~����*�bt��޾r�kI.��yGx�@�P��Z!zH���m�<��\�]]$ �:[!k���^��@������Th8S�%K���vj�en�kUD�Xk�B4�߽#Q����E���X�����h�n8m
�J���\N�n���炔�.�8�x�@ti���M�g�����`��"�D���&VC'�Bx?��չ
�rO<Z�:O,�WJw��.��]��qI'��Y�̟� J�'����c�U7jӐWv�*ղ�S�YT�/~�y&�?��qiU�ݶK��g �Vac+�!š�^-�L�
���* ���|A��?ة|;eK2oVbn�E��p�u�zP�i_8ٜ�7�������M4���dBj%K�>��0�B�</�[��:�O���购�Mhx����ss����q��|T�37\�㣂�Y���ۤ6�[��h,�w��j�UM��s%T�mcjXVj?;�j.�vY�t�)�J�%t�������t����v���oHp���o��8AU����F��T�������ڥ���K&��Z\	��j��v$QQ� ��R���,+_h"�U��V��av��'7\մ8��W`JS_#|���eGHs�b�	�<�oFMᷞ� ����M�ۖ�j2``�KP��+�9mȉu,��TB�6u�O��9���ِ;�+�f!X�cX~UP�eAV��y�h�5����Xs��R�Y?5����tL���4�Y��U�;�5�g��F���P�&�����:}S��7�RØ�j�	D���D���o��ζ�V&��)����E]T����"�)�ke��obM�M�6�=�U@���5���R�#mذ�/�0(��ϗ�9����ͧ���/�I+�*������'�gꖡr,�9����f���Ʃ����"J	W����q�E?��.mK�f0���]x�jd�9��=���9~>��(5�^��c�f�`x
�SVT�#���F�_����v��T:S[C9s%�Ux�2'{a�lz�k�#�Ќ��6���.�����V�)�j�
�e��W�����;�,*4��U�E�f�I�,W�s��|t�-C�A?�ІKbưU���w��d9le'FΖ 1�y�R��4u}����z!y��s�fԭ���,�}����O�"oT��m�ni6G��B�b�5+���ꁼP'����.�����3�X�$�mE�3�s%�Rq�����`Z���o�}������Չ�$=�����:-��͓>1{��_��i�6��4�Rt�(A�y0��
�)�/�V�[Q܌z���(7�ji�FBXU.��;���d-��rˉ���"�FX�r[��a����I:���m�1��������К������CN>��p��Sv�D)RKR)��jhtS�C���%Y}`$Q4�Ą�C�io$���Q\���=��d���cN�+��h�C�On[�j.�X~����v�����7G����@�Yb���w���k�I�Y�>�ztCLٯU�z~S�ĩ�S�ΡH���n��|�|���^�4N�{�r�mQ�������3��,���p+:n/��0��9Ϗ�3:h���� �5.�y�@I�+��;���\���T�L���*��&�0r�,[~���0��z�q\?Z��}�@#D�\�Q��1t�,�W��ƙ"�(��ꧼ��l"բ������R6����ts㩽��%Z_,a#���[C0���˵o��f��Ĥ}�~�����Eu_ʡ��7�[���174�0l�;#�M��nI�v�@�+�Ԓ��9��**�Ut��ݱ\�LvDRqP#��h~f͵��*V{���7��>۔��*���n�[���L��{�wVs�;�}�i��V�yI��'�1z�C�
�o�'P��`=��weW�@��5<�m)�p�W�$�.M/]��.CD�"MX-+L��������YI���0��n�V�ڸ2jtb�\NV3��wH����%�n~->BӠJm^���Qa��nJ�C��>�V��ũ#^n4�-D�$xR�&���LL��Q7i����=����c��l�V��u�-�R��1�^���G�Zގ��J��Y�]�3G�7Ʉ��Ӿ(4�5r�n�jԓ0ɺs8z��+��y���ZY���)�L��))'bu�>��N����O��&~WpS�{j�j����XDՓu0�=�9=��7�UJ�\L�q1ug/]?�E��F�/�$�b9]�W=g��[5|n�$��P��CD��8���D�#�����`�D���N��,W�gS�����>;d�<+/A/4����m�x���^��g;�ᱏ��L >�h������
݁��0�
 L�L�Mt�"�\���A+q�)nk�������}YY5"96b�͙�+5��|�)X�z>�k��H��eh�ƒ���ø���!X�}���/��a�ض�NO��".�K��h����'6j���䇼J�$�|ȡB�.���/}e���s��W�F:~)��"���q	\< a��T�4��F��}�B�U#���������S��,#����y~�a��Jd�܆����&�>'O�薱�Ăj�����0�#��DU_{��)��4�A\ ��|���E�j�����0%�oI��ׂ])�����8���f����V�Y�o2�*AEi$���s#��{7��V�?6u*���׻��!�����1W�G��Q+��иe�{M�[��cO:k.��O��m�
	0������ ������ s~��	�t��ۆ�(`	�������~�Jf#��W���E+����f5��8��`��mR�r	C9�����WBsum�_�� ��#f�Cx�>�qd��+1e�Z�#�pyXR�	�ܦ�PX�'1ʋ(��� ��^!��@�����%�z�O�g�G�����]��M���Q�p���l�&In-y��Y��{�FԦ���SW�8L���Φ�B��S�����<җR�2�����؅!Y0����3>�GoNv�����;��sn�EF��b 9hQ��n���ً�cۏ�_ϻ�#\��s�*pɩ��1�oW���~��y'~0�u�:`���8ADB�<!����.4S<T�ǋ���Q��r����؊�J5�5O�1)gM�Gep���[Ոa'3ջ7�S�>��.#\q��&�>��pː�nN-N�D /��1w �j�D8�k���d�Hi� ���J���hY��4��-��hi���p�U�ቁ���=o �8��eX�R߁�kmpf��Ȫ�^c!��w���l�'�������e��K¿���.�pơq�f� ����u�T3Q��N�\C���$�A�B��3Y�3.<���m��;WF$�. ���1nO��O�Оh�z����jG��q4
�VQ �1���{kw�R�+��<�,��A�-�:�L���O�q̑�g)yW�`~����q%�wT����FR�v,��)�-�l��e>��x�4�a&M2���L\���6!c�Gw�$�#�i�#P0H��d(u�vۻ�6V��7��KLHcm������`E��	A j��f���0�ފx���0#���!_	Gʨ9��8�ځO���b߽qA���{Փ�Qҝ3;�`�8Z��s�����5�EҤ��@��b��@�xPm�oɯ�x��yx!�d��Uqy�U��
���YU�*�znj�9|���Ų����-��"ۯ���%t��i�(֮�%���@��VJ�%n�gٝW����+�����6&inCA�e�7��>��ԍ�Mq }�8{��T��8Z�{7�8��2����q9�W���oy���Cäv�q�c�I�݇�l'2H��*�1�O*ɂ�c�y1 Y�*��*�f�Eb+��7%�z[��h6��%��<k�<�G��fO�=p��2��ݾ�S�ճ�؀��,\@n8��i�/C�,~7\�Ma2 )�c�G\h3^CR��IN�@���H����q8uAs�'z��N�oh-6s>�v��<ʶ�U|��+�V�AO �GC��.�Yy�#-���Z��tn��2�)%C��r5�/�	 f}YkHK�NZ�t����̃���8���:��;[����>?a� aO/������僅�X���:�#�����A�یw��"��D;�[��ꯪ�m���.�nj��.J�E��t���e����׊cZ��Ֆ�h�l��ϲ<����U��te,�hB��1L���=&(Չ���,X������u��i�@?���0� ��G�=�/{J�L��~�+v���_���9�4�ZO��U����~������� ��[<䀭@(�)���y[��#�^�>������EN\��C^+Ye1���I��(�7�#�%J�p�k��BX�����gw��bP�Y�\!Q{�S��)����%�&j��p�y8T�`��2�m>UX�n.�n�BqMa��|��>$�g�b��W��I=K��j��0��3�̢��1���`M����`�1n�Y���_�����٧xD��лk^�9�__�_� �H�)��<#Cܵzo����� >Y}�z�O2�uŉ��qZ\�f���%����.�V(ve��\����>f)�lH�\\��K*~�x���5ŖX�3L�Zpz1�⥧N�Oܮ�$�Л6Q#�,�
5ed7v�X�"z ���_M���iH֦��
�zR"@�Ty�h� �I���jM���5�v���&T!��ЍM����l˘���n�v+p[���2��S`����k��B��n��2�{���
�W�S�[�����b���zRi9�`���s�G�Z��*�d�;S������
���Dm��%=9�=��Ȫ\�����C^残��#�����f��)��Ϥ~�0��G�u�E���ix^yO��_�0�o����*.1O�����8��a�p��� :h��j�[qꈼ|�U��Jj�D W�lھ�G�Ð5bd���#��t��	FO�B��7�3?*'�Z��/ �TSn`U���o=(WRi�P�KS�,�9�kr�=��Z�6k�8A
���Xyt�R1M6��]O���Cq!Wz71`e��ˋ����B�Y���\lgf
$�[��CS�2�]3^p��L,;cD;�9F��X�,���ᗢ�vJ/���R��^�W �̼���$�P(����z�Lq�"bgR��τ�����c�e=�L��A�pΊsՐsT�Vj�_Yr�R	3
�q#+E�ݗՄt,B_;��40E/{��{�$�|�>��1��
�:��3�4Xߪ�Z��a)9�5�d*����^��QY	O�A�pbT�v�߶"��B<�,E�ؽ*El� �wf20�u��9�9'5,4z����N�rtA�F���(�ə"*�;<�;`���4�ϸ I}��ȗ�~��*��[���
i�M����vqӻ.>>�)|n<N��=P���)�G���z��+[I���2� QWĥ��X�������dG��b��)I�\h��m3뛴^���%�l^3���d�n>��K\#�~��2��'奄�Yh���x��X�<�z. ՙ(�� g7�.Q��J�}�d��O�2ON�e4zwRT���Ξ�<$�mW%��^��P���M���2�X��D`��j�v��N)_�s!�/5��i�|��h��R�����
�-}��,v�[q����J���/>F�#V0_��;�z��F�x �.E�EU�tȶ��I:�{�i�yƞOW����ad���=�ط�7`r��ǐ!����3��̌���(v���Y�*����$%�����L�'q�s>���[���6:�%�!���K�D�gh�B�|��@[����bw�hf��Ĵ���_DC�@�v�l�d�.�Ӓ-4�+�/}Y�5���tDc��`1 V^@���$H�Z��xz�.!� ��[	����_�k�ֳ]�}�V�2W��ޮ�:K$m��d�1�P-gILы%�PBC���ue���.i�T �P��n�֭�6r�kA�e�j��r�pkC�JL%�^��j���߁�g{n�	��E�Ǫa��$rw��������hJ��������惌�������Ԩn�	��,={|#Yj��-\��_}���!t���Şx~�v�J°�-�����S�G�T�A.����g"s�E�=�"����� I���L*,P?ul�l1�:�.",�����9��.������bp�z�=��O)��T��f�G��i��#�p1��@�A���6-_D��M�C"I#3��
�S���,HZ➠��>>�s������?�61g5��W�8&�=��p��Qa��g��9ߠZ�ӣ�n��m�9��׮��(Q�x@���v�B�3<��>1�)��c���쉚��������H�i�dk���J�[����7���}�)��"B�-�ƺUq�o�~F��~,��@���gf�~���u����OݽI��/D�^q����?˓َ��7��[29�8��k1]�8��@���^��3�Y�u�f,q�K�h8��
����o�4	�6��;��M��9�ӹj�h���Zf��Ei�iR�����y9�"�p�[���|���M�\+��Vi�qC����E+v�ǻ���mZ=��t���4[w�k[�:��4�Q��팜��i՜p��ǳ4�'b�������O�����6�E�f����ێ����Z�ffD6ĞL��ITz��-;�5*�|�@ȱL��}�`�e���C
�8�M5g=��y4m��&0�;����P뢦�����Hܗ��o�+����������A o4t.�.��'4��*��I�S��ݱ��C�$݄�tF#���oX-ŭ����� HAԒK!���;�ɧ��D�n�n��͓a�&����&�-7���d%��S&�3�"{�Ǉ�NE������*���\�Ժ&e���g �L����_w��`nQ��*�� ��tE�"W&b{�&ۦ��Dr�F"m�:C����)m�*�M�����4���I+�7Ȧe���Lߟ�Ma�M�>�)���[�As�F?\a^��lʆ�~�f�ň�r��=)M],� Rv��`X �}���G����0��~�F=�*�����J$������4�2��+���:~�yf߰F�
 #XmկO5;!��r(�i�*��j�\|��y�C�+�^�}�u�����n��EÓ�wx� ���m{�_A�;b��] �̨��x��] �A���U��&�d�A����I)��;H~�8�e��S�wI
Н�Wy���qg$�ʈx3}L���]�;�y�$�����Ώ����D���Z�:B���:mW\�M�I
�s���#�lv!�R����6�N�����z��W�H�T_�:@����q9�s�A�ʩ�v��4>����Af�������Ί)����NI�4EI�����f�:It�;h�ˌ`�ge�aޜq/�m|��8K�}�VV��\��q��d+0���J����{�k�i�%��ʅM�) �vz��_���*L.�'����2�|����g�/�˧��`�χ�+"�8�HB]2�a��V�/�,��*&��qq���2Z9�c���Q��}14Lڍ�6�K�.���;Wd����8f�[V4Xa�r�^7��5���a� �����.,�,�)*11�Ƿ$h���� 9{m�'4��n;�:1 D0ߎ�u�Yios
T~�d8��IW�㣄rl��$���49�����|l���J�7�� �c	��:<����CD���8�$O�*M}FR�_-��ؠ�6�ٹ��u;��q��a���)����.B$��SoT�[�U �+S��
d5ͮU.>x�F���v�?M0���]��R�<Hx�"��n�{o�z�q>g`F���A3;`���fn�jv	^��/��v���);��I^�(�D�'^�2]{�Y�{}�O��W�M�y�Э=���:�Y�\������N:َ�����]��:{O��,4+Z&�D
\?��.-��_+P����цէG���s��q���|��c\�Z�����%,|:�?�7/9�pަ"���bgS|dɤ� ����˾ZS������	8�% �C}6�la��b�(NC. oU+��iV{���l"y���0^�&&4�S��L{������� �(���n�7}�({@f>��h���C�v{�5�E�������>������6�z�%:��,���T�����JDegJ �@��F��Uػ;�'H�8=��"�.Q�n����;Q��%����hD4�G�m{��8J�l	�B!VP���ָEH}�1Kq+r{��Cw$RE�K�m� ���(ܢ4ݳZ�����p��kJ� ��q�Vj!:��{4�_S���ŋ��T���	�Z���K��].����8��;��؏"(��	�RxO��*���;3\���i���R��XSfx��*u�j��z��#��8�#!�[��q��������'ާm����8)� ��/>a�gf�rg�ֱ���
_�4�W�������@��Mo������S�=��RV sN�Ic��D���+q|��%Dk�M�j�Z<Ν�d<[M���h�`�&�V��D����@)��`�$�ҩ3��t�у�l'���F/3��|='C�wp3�WІ��J�B�I��7����e'�A���]^\(�e��a�2M�ǿ���l0��8u\@��_3�%(�J�lZs^��v�!*�IoX���N��*�,usy��,H'BXs/�7î��I'&fh�U	�V����I�@�+�HSR��P;�N=uM^�&�*���*�[�ĺ�e0,4������=5v\ޫ�}��1�ި�&5�e��<˧�7��ن��.|H��
%i1�����\���3�����He�P%z�G������|Y���t�H^cYTy�$�(É8$�	�	�?\[���'�3�^�1�����vĭ'Ԁ�3p���1�V�� ���l�J�x�鹚�zB�4[�Sе� ��W�p��a'�'xJ��?{��j	i���^~�V�q�w�E��S�?1hcW�榶���<��q�Qk����m��"���]��J�* ��ȗۿ��`�5���R�^vF��XYБ>�#I�[�A}�����L�ȵ)|���NB�F�����;E-8@�=Ef6���7�뽻���9Gɯ�9I�
�Q�J)/ȯl4_ۢ�Μ|sA��OA����/�x�c�k`�c�:t!N.͌���DCނ�g���"�F9��W�Dn�G���C@�sEy�@�
y���_����������O�&���.�Q47ɱ*��&�@;^��}!����Y�e��{��������}�I���L��w�W�X��n�6�:T�w��!���|�]��f~:�C���� �-O�DDsQ#�Ga�2��֍��&J�y�y����)P�\�R��8Mih����r��xjL=Y�w�<�]��������0�i�����y��q�Y�۰�}������P�iD��_�67�6Ӫ 	���rO� x��n0�[�\�j�9: ̪�L�WQ� ���ۖ��g�hdГkD���yH��gf����<J��<�F��B8����c���4�'mEi�t�P�sX:P��nh1ƾ�g��A�O� 0�{�4�T�l>�r0ƅ�잧�(��K�yt ��z���R`$��4��}��[��ϲ���k~���3"؞0��-�8������e#Vs�� �	�A�(qj�Ƿ��yM�[Y`upY���6�������k-'Pt��v���\��V���q����� �J5��IyH����:�����x�m�5�쒜��a�L� E��v{9�������!�{�h/�EЙ�C�-�i�}L���!��w!�C`��O�� �S����i���NYL�����+��眩a	�z	Vo7#G��Fw��a�DH����N�{azEhBjr�wF7 ��{-�2��'8`�1�QǦ)UYFY�Y�����#wI���Id\�jA��9
�7ұ�r�]s�ϧ�[^��a&ʧ[9�9�Cȵ��g�@nu���-�Dy���,/�$~yi����(��?1��I�?
W�EDA���pQ&&��1?��q�@
����I6溎
6���+��-
�Lx��/��������6n��QDH�|�Z�)����b���,� xD�� ��H9�2���V��X�,|�8~� �|�����4���\������W��	[��AvB_8ڔTgr�z��q�ϵ6�Y=(�R*濂����\�8�Nnّ��|� �q��.���xh�s:Ë���h"�H�_����o�V����/�x��"�UHZ�6B\�3e��^c$��:%�5���D��� �ZR��a;�Uq�Z��aL�m� � �Ay����c� s
������bZ��0�+�{�Un/�q�43D#�t�x��z���|w�!ԧ��.�F՘��ӶGK�~O�b�]$�^,�},�,�cS��*����U�s�s�ꣻ�1\-�,˦^���Z�G*!���m�'���G ���$��%f3>EW�&��+��؀*���'H�;4Z��FO�_��^xm��B~Rܑ�<�Թ�щ0�Fy�+��Ȇ�Hƣ:�N��(Ӂ�I(��!ם�q�)E4�F�% ��87"�LN ����F�i������G}/�Y쥶�S�L�0He��\ka˖�6��Ҏ;�J����r�\�۔G�[d�hd���B�oc��B|F'�t����g%��"½ۭ-�~����/�b^�+5:��ɵR�hކ֜�^��'�6Ý��=d�W2'�S6>��.��	�'f��)SI��v&���1����
~]H��ʵ0blJ��p�Ǩn�*D��ղ)�i��P��q0��~/(;��� UĉJ�VM}1��b���`MC0E���9�~���9Q5?r�!X��g<p|b��K�Z�3?���0����$�f/Suj3���� h�A�^�uC�Ǿ�K���Co�V��nd�CC��(sf��u[F��oH�J<��+��[a8�^{%���%Y��o]�~rl/�A1n� ��y+��Ib����}���}[����sW�u��QI�\������<)��*ʔ$��+s�^�\J-�ۢ�� HH��U��a#�LC	��N���o&�<�;|�����Y<ҹ�JZ�C%�.Ƽ�������w$���.us;�u-q�G��". �V�=��:Ь�Ҭ�FJ�[����?��}?�.i���SD�Q�x���a��1��Ug��!����`t��O��˿g��J�eZ�C�
�ֵ�E�L|V��f�� �b���Y��S����`�GY	�쇢R�5@�ڳJ����6��i��.}��2��l���:P-��D{߹h�����T(qxq����mE���p�%�D��V�}�r�%�z�$x��P���'�jN�ϫ9�Fw +x�;�a����A�����'����r�򚄅CbT(��̙Ʀvo�y�!��FQ�����f���#Ą�
�����n;��x�]RGuk����h;Hƃ+�����o��ͦ����a�K���<���oK��(���,uE���4��&�v钸g�7W��nk�A���[�U+e����A�|v�`�'���n�;U�@_�YVQ:���a1�zUW@�e!�*��}��5�d��2�?J��c��o�[T��*0%Vi��Ƙ�Ȋ�-0z���{a� ���J�����:�c�!g��BT�4��S��eř��gZ��o����:� �.�+HET�zv���ׯ�����N�#���
�/[*��d�� �r�ឭ%(�D�۾kq�%8q��-�ٶ׬/��z�sLl�!:�+�&R�C��#�t�Pnn$�"E8�3��n@��mXg�5���4���>V���]s:���!�9~5�Q1'�H ������d25i�� ~.�cR����`��3kr��t����-�$����w��ɯ�S���G �z:���S����e�H�{v�e�'c�r��s×��Z��F)԰����G������­G~@�P�f4�CN�l;�G8�@b��ť�N}��_���4�v�Nk�c���=�+���D!άغ�X!�"[[5{�S��K���PQa2w+�����`�v1�p\�V옺k6-���9W��N�q[A�i����L��������M�$��}���E�k������f�c�L8�t{3I:͋�,P�o�ώ�?�l�=y�Pd�ڂ>e�R�(��G��ѽE�����dv�����]�a��'�v�hy�V^��_�X�M!%Y��y��|�{������կZ�i#j��G��������ƣ��_7�O9�2�$��{�!�W��o���e�� $.1�脗p5��?/F���dWi���\�x�j��1g"���ڞ3�=�C�D��8�� �/2(�J���$�!mm�g����՘�$nW��׊��Ҫ��Nȋ���w�̔����GśE9^9^���ɒ@É��Vn��Y���v�ן�
�����`�ïTl�C2�%ȡ"�G>��'A=8:<HU�2�QpD����lB����Om`X�����ϓ��3t�)��%�g:��[�ˆz*d� �]vbp�R�(���u݌=���I�Om��bܗ�eI�X}�E��#m�5nOD=и�`�D<�����ڍ>�<���	��F�ͮ�vqϓfm)������)���痀fk�J�Pb�����Q�b�!H��{��;նk@�V[>0�z�������/���������~�����Pk���ʯ����nO/�X�_��kJ���5�)~;K��,�w�+xS�17T��Yz����fC��^�9;F��'x�o�	��> /W���Zvd��D:ݶI����J�O��'�`� ��$�N��%1-����ZP���<Yt�P!�`�@�����8o��'����'����I��aD&i�Rد�0�(5����y6�Ȭ��#���;"j�<�-K��<�f��O/A�j��\�@d��B5�Z�ڷ.��i��l����<�O0�ѓ(�o҇�r�$���[�#�q��`�U�0 �!�No� Y�4liFi�@���=͋e��Q\�s����?�Y��s��ݏ��@�<Ƃ��d����U{"\�|j&g�SR���
L�6���A�n?�rE �q(�9e���ߙ1���xZe�B�@,��  �:��H&�s�\�E�DMɳMV� �p�$.��[�ݦ�����?��/�^��(�ǥ̀,Y[��幄x�^�Ycva��ᆩ{�޻�-_�,ƔQA�!3�%�ꎮ��hw+pf̺Ԗ+Djh��:K��3ƪ�H�]E��^�kY���،̚��!��l�t�����|6�W����~�`�R#������`�7�r<�)y3�ؗ\O�C+PL�VɈc�y���ff�[����k���|�4"���>�0�����]w`��Z�!B�7��o��~j��K�{��e�s��$��"|v0�Ɏ��65�My��yx�l�b��n+�5d��?l�a�	~����� Զ�
���ş��4������6x�c�T�H���X5Y��t��/���B��PWk�KyI����r:�je'm �A��\�x��g�}
=�^S>]��{��@��x ����[^�{��W���"�ͨT1M�YF	A��f���Ʌr+D����&6��웚v�FҮ]Ś@޽��ڰp�����c>��T�Z��4�R#[�s�a� /[���c�l��;��0{E��d����P��Ro1�V_�[�Yz�C_$(@|S���5(B+BqD��X4q:�l��4��%V�����t.6"���O�o6�4*�"���!T��e(|�ɮ�$[';�@��j��D�Σ7��"ƛ�{zy���lV� ��_D��<���)+���L �*F��jj�Qjnf��=ā����T����f�K;
��/P�&����8�j�P�� Ͱ�[ô�o1�}ki0�����u f�Tl!�])h��8�_��@nj�I �&3 ��K���H�+)��' ����L�6Ҷ��/�<_;H��EL�ʤ0j{fbn���-�����Nk 9��?������hd|Iأ���|�u_�~�YrQ�������wH������<R�7��i���"�2�;�i���U��r4߲���,��;�ث��*=Z\���n,�'�B���R�Da�=n��MP���R�	��>�?�x�e������,*��HXQtK��B�__��+3fm������Ǎ �,R���m��r�D�/����þoS�d6�2�{���p�ca<\�tG��\�(��
{�Mt�ߝv*#)~�����Tn��zΒ��R#6�-W�I����+�"er�nY���D8����A9�#�7=A�L�ff��?'}*Kbm�)���������]�3���1�hC�ԜR�ae�׈�@��N:d�#��?���$��Mq�i��O�$���
�mA��$������ʣ��������PU��B},O>*��Դ�ӡz���qf $��w��a��E�}Ň�kh���2����4��?$:ɚ.�/�Z�rT*8$�Í�F�Ey(�
�S�	�:w�ӿ+��� �}�D
(�ϒ��r);�)����2���1  5x�ԉ�?�^�n�gK]�F�k�u����3#a�	"����ǋG31�v�	ys�Ɏ7��_��Ｄ����T�,^�g5���p[:ԙ�p�t)~�~3Kۜ� ���X��Z��
Ũ:��������uh��/����.�;��N�����7�\2�w�D@�A}����L�7�˶\�|����}{1p�=zF�9��N�I/j�3[t�t���Tp{�Ka�g��>����s�T���ilk�!���T�]x˼;��$�Ι0X�O������@��TL�f���b����iz�w!�|���Y��Cj��;���D{Uk�M�:�=>j�c����!��d�����8�Ze��;�(u�'������m�gXɤQM�>`�����iԾ�ۙ
D��`����b���[e(p�a?3Cr�yC���2����Y�1�l�+�#P�C*#�<�:����DN�(!�⹩hErp�P9��U�v_���͋ߓ6���HZ��pN�}�O�`��P~fG��Nd~��Q�[f��,���f��.���Ց�ym�S� �a��I0&˨����g��kqU}o�����,*w<�+�\0L]?�C�xG��!Ǽ�t���M�8�-l�{��Bǿ�I}7'�~�1��Q�u��
�jW�pg5��靤��!���܋b+]T36{T�c��v-3;z�je"��D"?���4���2�G�RTS��s�엷�L@!�|�nȑj�3���g)cA|��e|�*��?�c.l�� �>`��|S��ysG���&?%9P��ܜݛ�P߼�H we���TS�YV�}/��^Զ�Mp�-��[@3����n˿���!ԇv�-�*�ĕ���H>V-�}���:#�N������Z���4�2�n�`�Ho2F�h.��$0,���L�q�]ࣚa�R)�Az�>��Fܤ��8.���K:["PU`K�Y0�9R��JE�5t����Sφ>}���af���$�j��ԚE&�4``%�$�5;��ѝ��q��p��\����_7* k#�Y��'WD�2���fY��W�w�j𰗧�E��/�3J�����q��~d���?4��qM�|��Csu��5�G�n�
�������_l<�%��J詣S]����w�U��H
��>��y��B�M%���_�#H�G"ߑ�� �8�5�$f�	Q'8	g�U%�PV�z[�� �БS�C,׋~ݏ�����͟���N
�Yj�J�V���3����£��Vçnۂ��]c6 ~mt9p(���z[\
1Xa~k*�} g	R;F������Cj������좹��L�g�h#54�,�&�Hk�=L߀��K�z 	r:��ʊf�ԸT��55���z��fE��UbX=�aQ~>�(�=�`�9��/?��Ȏ+8"ǚ!���)'n�Z1C-q��չ��q��ə�mM��Q������Y�����֯"z��t�N�(��j'�7� �j2��K�@�xN�����&�Jo6�{�?=FM�quk�:�R���<{W3`�	X��J?�;��
�;C= ��od$X+�5��ȋ
����yt�[��Z:�WRsd��4��Rl�n�ٵe�韮Dt��_o���|Ϸ��f�,��/�GUSO&����}{NZ��v!Z7}�KӓJ��n8pL��{3�C��2Uh�'+JK�u\�#�\5�'ē(���c?�H�r�:P�.�ê���C� qE�D��/\��N�?�/�Wr�NPeYF�+ ���Q�^����O�ҹ�JH������S��=�F,P?]�r����05=i�底ao��X0k���	ow�Ǝ�gFVE܁�L��N8��Ófi��S	�h���$̜�	|��3Z�7�r����A]���iA�	;�� �5B�����?(����H(Z����{�46��{X��<���v~�)�ķxm������X]mZ��*AI2��M���ykC�C��l;V2��Y�x�v�����D �]�vnc�k��8��Y�� Z��9h����\��*6���Ġ��8?V�9Et���"ZJ"��׸�Mh���zT�K��x����LlN2�!}E�\���qbL`�+p��&Ln�Q�~������e1*Ud�!��
�x��ѡ�:�=�e0 �ϚE���6Ӿ{K����/×��v��I&g�f�d�U�4���5F
Sb�b>�d%���=��1IK�$�pISfp35�P/���8z'{K�o�66c��i��Sk\�"��2R �<�fG��w��.xB��k�p%M�P�����7@��-��n[���#2'��r��$(���!e0�a����9��7�"��,x�Wm�/|*���*��r2�0Ļ!��+hY�(\�5#'��o���Q��S�u����_2�������y$��s�=��(2U�I�$B[�����ć�+��\]��X:�i�<-��{
�GT�)+e.E]A@����n���m��yib15�#��.�:����[W_����XPO��4^�_��7���d��'OIzO�~���HaH�[m���R�u)Q��n7||%�\ƱF��ϱ�1E��#B}\:A�W"!;�yG�(	���2M��ߏEN��:�e;š�V
hѿ<���,x�Ѷ�����L�ӈw������f�) ��0��x�z�!�jG��|�!���Lf.���^T;���A�t��^��@���/�_2�疦�P��)�P5�O�`2��C���]�����[-f�s�;�eY����\ݤq���[�����W��V��"��=J�XQ�6��hn⹚W��
Il�W�+c�or:�  ( ��4/"�c)~�j��`9=i7��[�������ϕ,�c���=j&�L��|�\�,��p%��a44>pa�,�UJ�g��a����u��zW�����S ^��T�D��m���_6֍���G��a�v�NX\�����0YZ�^ -��2���w�̣�<̥�p������4r�����k�����3	h6��+���O�%�kf�tzϏએ����1�oD<̎h�Ձt��å�e�B⽗��OҜ��B�P���t��,r��P�F�����p�p90��ݒ�jZk���>��̹K+�����)��S�[u���u�w�{v�`ZΥ�����Tar��%�]g��I3E1)���9&��͌���������&�ry�\�t}�
WrfCddV��X۞h��� �U�^aV���ԥw�k� ��t�������f���!�������kk�]Q�rN������H�ꒊG���#�BƑ�^L$�ٺ&"��4��G`?)��0���1!A�I�f��Nx6u��o�I�n��r�ݰ�<��}!��y�a��*��> RS�#J~]#^���kPJ��_�!�`��P����Yb��0׋�|qkɅ�s.��&�\V�Ipս�����	F;G)yM��s��ႆ��Ki��˳W�eO$9r���ro�n�K4D����������G������V.����(_��U^O���ozg""�@� ����n(�V��v#��LU��k�Z��ЩuY��,�A����Ǥ�]��ėQ��*��~���!=�lj�K�Ļ�#,W�04�*�<ߘi�Bd7�t���mj1d^L�hV�Q�sf:��|ƀ�.��1ʐ�T2@��Ws�}l /Б�����h�A���dUp������c�63C~>��îl>4�2��]J{�*WT_�_O`%*��]&NpCc�h�0�T�_Б6S��*�aeL4�Z�,�d�����>�V�g1A��Nl�e��5��|NjB�@-ϳG���פ:���xg7U'����9 ��f�.z��H$z�+Gd�+�ag���cL[}��7��Ș��0��.�N���=LM�D[�w�H_
u�ַ����%3�/V�NzFL���8P�yJX�������Č����#E��)�d+��V���]B��q��fq��\G����#<^���*���cCQ��%'Cᚃ���s�T�w�d��5�?�����NpY5����iS4\ ���Z~����p�p������8�������Qo�H�j�P3��ݖ9B��/�\	6% ��`o��V$��|����~���~��?K�s)OL��T�\�D��^F�*vM�� �O-�!x�����Oz�0�8������[�rN)������p�����T��ܟЊ��������R9�@�T�Q�Q����_i�*j�d���t�����;9[�v��-�����p�R"�Y��^��|8�B�8^$9��}ҿ>1�ju��E�}�ϸ�(��jg�tP�gX:�!�qy�@f�IR���-�XX���4 �$n�'�ޜ;B�tߪ���C^6��A"���h��������S>�������?/�,:���:��֚���QTk����DŇ���X)����LEc��Y�Pe:��u����q���ATZ��ZP�6��ukf|\�}erm��%.�qY�+�X�!��9�5�8Y���@�i�ޢ���g�f1;r��jsH���l��X�����-ǔiֱ��V@L�N)���,(���b>�w�,�Q��Gt�Z���a�Kp�K
�>	� �.s_�y��/Q�����~\H�G�(P2��U p�*������������7���y��4�v!�k$,AkC��A5qFc�T֫Wz]�"��-��p��DokcL?��pq?�PP1�/��B:��&~{��.��d�M;8�o�v���M&���U��i�r�G�';M7"+���"/�It�E�59ߺ �tu���i]�^?L�^�h���e$��'�2!<3F$+�🙢&{�~sJ�`�w����dp�}рR���h�'c�4ĵ�PHD�([�if����0��ř��O	p�k��.K��{����_ ��+ƽ�͒�&Դ�Q3D�
��$�hc���ю4Pd*��O����D�!:�b�&[��4�_��U��	��sj�U�l��s�O�����Xʢ'eTu�.L��T���nj��9��<��*�{�{f�o����?��s�Yu��-��00]C�������&Q� {�%�ӤT���y+Q��B�n!��כ�ރ����?-�E�pxa��\2y����\��E/�8=�$�V1\Q62n�Ԝp|h�bOG4!�1J����A�^������;��I�C�$���O�T;��j���5�wP�g�CֆR!�3���͆�����5��
�l@n���br���*�8(������@�����i̵���:�ĩu��<����Ɂ|5�7@��)2�~E���hD7��hL 1����b#90�w2�>in7��y��n;��dჼ	�6_ �_0Yq9a��)k@]Ĩ=�z&�Y��nv����vm�ZbK�k^RW����g�<_��+0S�*��A�K4i+�v!0.�h��]5��-���\$Ŝ�R�-�Q}H�y@�ch.<���E�W�R�L�LRA���υ�ʾ٤�p@�Y��"���=|T���5�]��&�̐HK9i�HW��b�6f�%vKoYa��e��_'�>h��[m��R����w�ս�ݾm[�<q�re����w��ۯ�{����>|\{&��F���+��`q�$��z<ԛSu#'��B�%�k B���-0�/Ӄ�S札��e��;~�9l��Z�}�C�����66��e}�Xy"�>l(ђ�J'hzm��*ox�ZF:s�-����s	�vߕg����7ц`��й�Ø�� -z����o���'V�����+��Bpw��G��� �+���·k��]v�e͂���}���В	E������$� �?���7��V���|>aN�-����0G����D��Oi;�ތۗW�NtN����"�|���t:�#3yAQU�=�C���9�Y-mG�k�y�S�ӜzRe���e���_"��g+/Ŋ`k����,2A�5���u�WWu��y� �-�[��K�AKS���H`r�k;ȁ}�$��6C���n��Zz�����@�;伍P��ƂW��4"*p
gN�׎�����^��p�!�QCU��K�����Gam���o����!Õ%��+��β�X��� �C�b�����Uڝ\C,*ѕZ��S!�i|�>l��Q�Fe��������F i ���պv<Z�`��C�{���H�c�^�U�����]`wH i�T�yp+�iX�Ǯ9��L�nգ���c�{:��y"��g�Ml�D|F��}�ORO���<�.
28����]�.@�]���J?w#�-������{�gU�f�p1��斒U���˶�.HP��c�T�E�I;>��[k#��_*=H$L�-����f7
s�i�?hߊ�ӢSmU�T	B�d�>��ׯ}@��uTZRnQlϱ"��ohv�E˖F��ü:�AE��[�cg]����wk�!�{����k.�RR�hKؔL
�XI��}�?{O�L�� ���C�H��
�����\��b���R��i�B�ۦB\	Wn{x���ڻ����mp75�N[���?X���#D��3���)�&&^���9������پȹ&t���.��tW���ַXQ-%�9�p���!_]��*�������i��v�LA��>X�6?m!�ϐ2���b.74t�>���5Y����=�@���7P��+���z�y�?Z��`;S��U�0-�	�cu�4�+�m���:��6��]s�(vg{��uobY���|�����ȵXD|�����"?��."���p�7����I)�Ow�S������	{]�6��#;�-&d��Y�������O�6k���,���������ww<����8���8U��ᰘY6�P �n�x�i�m���0�t����H���736}U��[� ^��㰋�X�������$�<n_7��`�8���a��ךsZ�+�B?:��a��3�0# 4�f
]j�+������8].������gE�W(�9��{��i�\�z`�
�F3��m���z��@��=-�X�j��s��R�_(=�<;)$W8љn���d,�OZT5�ږ�
^���'BX�C�؋i+ݮ�i���ՄK��>���Y��o۬��3{x�&�i����1d��J>�kR�����O��Ǻ�j}�ʈܽ��@ԒNk�M����pX�|�~��R1�_��eˢu/�M[}���NʵإV���>� �cT��f8(I#��T���t׍t�_�<c/�B5�Xd�43qF��58)t�5��I��]3?���9iX3��tK�ʏ�(�?�h6��9O\�>l�Z����f���`=�Q��s�I��i]��-H1�V���\<�@�Ts�P��y�d�qx��g่ǟ��1B����X�l����V͠�A�k����gd�aA�����H�,}��Y���#�6���*�����^�<Ǘh�V�|�]�5l�Sl�#�����8�v��/q<g���O�&�R���g�b�ۄ0{l͘�6y�xIw����p��,�i�
�_�u�wZK��k7�T��;F����ɒe\)t�v��_Q�h�#,�V~�HD�W��"^g���WcRث�DW�^�d�s(�ۂ#)$�|zJM�/���?n;� u��.��5�7t�槂�;Z�0�MB�������?�v�L/�Б�!B�`���|Y��=����-�!� ��q�C�71�[��$ϤIF���>�{#���g?�����:[��)��ʩ��w����Z���iO�l�c9�E�����������`�����Gչ�+,�b�G�!Gaj��g�&�?���ݽ~o�7g�}$:j���|�O�^F�pK������ϗ�ʫՐl; [��!^��~�oÁA�t!_����પ�[���bp��+W�����2�!	PXf��.�k���P��I����	=�P�������� 7 �E�B�Ou�<Ld8/o��pc�������ָh�Ô�h��^�"��d�����3��Bp>���;6��,��	7}�0��f�Y
�h�>��r!�����<��G��A���C�]`��7���]9+'h;�Q�KG@���<�5 ����X�%u�X��9v�&������"�㰜��	5�=$�z_vBu�o�2X:Q�M���*���a��S�%*�LTp��9���p���-(���P��n�cf��pE]P-O��;߈���P����)W��[���w.������s�&3iv�_(@t�t�|c\�Tn�H��*��;i���ꂴ:��LhtO*ѯ٩��b^A�.cp��,��Gju�0h�8u��퍢�K��^Z��[�`��9��(�VŘJ8P��"���q¾�z5���ױ<���w��ĵӲ\���y�Y�?����f?��,�i� 4!�T��w�G{�*W�vJ�D_�������)���z-�ӊޑ5���Eۂ��v	g�q\�.�=�#�=�]䕀��Ν@&��MȀ�h�-�d�����tn-(`��N�DN��@��_��&���_��RC�E��e�,�Ww����N���>�q�ǋ:_��qc�e�7CH��p��+�+p@����>{�wc*�N7�^Tr�4�$ś��``n^oLU������Q ���_��4�7jv)�d���sT>���W���Y d���S���B�X����G��ִw��ոx�E�-%+wFPs�C��xc�%^A	j��L'?q�[Tp��;3
>0����qf�w~oW@�����������M�M�<���L�Ϙ8�}wPH�{O�.��l^�Y�\s8�{��.[�y��<�q3,�������i���Ybm�ݐH�&A6'z��tOY܈(c��s!v��?ZL��tß��	�����!֦ڛ�\��7�$�ʾL��G �� ����*D�0,Յ��9l�m�!.�5�KF	?��f�٦�LuT��-q��v��cצ)�1��&�Ȍ��
�/l&�֘K���CŬN\�o����������/��zS��b2�X�R���1Y�5N�5���ǜ�y`#{��[���(])v��Y;\��Z��K$�2�!;i�A }ش&��-	��Z�A\KOwM���F.���Z�[��rƦ�5P
ܟW����|��l��DY,����ٕ�o�hJ<[��[*�W�>��w�#�K!���V�@a�I�-F���NAR���f�1�f����d���J� �ZrWm�qϦ���O�q���}���9��Z���X�Q���7m1Ɏ�j_��)��<YM����&B�r��f���r�!��5�ɷ(�����دK�6Q��/,�g��h^���B2�>��Ѓ�=�|��d����)2Ց>n	:��tiF}��F/Y$�e&�C��H��[y=)��o�Y�_Nm�׃)J`rT��؜�	��IcX@'��GtBI��n3��E�G�K*n�6+%�n���˫ܞe����2�9�"a�`��B�N�ɏ"�)�����_�"�Y\#���r��	����w�:m��D_���"e�&mi�Z����S�6]72{��=��"�tl�����]ʣ�������^jY�aK�9�79ľ*>�����Ç@���ͮ�p I�ޭ]�؉����]�ڏ������̸�p��}R ��}0�c�����*Q�ih"Ȯ���}@�@���iTaEԲ=�k4�/�I�5��d}�X!���}2�sȜ���f �c�>ڍ���u��������r]9V\�e�`��߁ l����@z���w�3�oc'ϕ]�k�R��(�V]|�<WW�0�S���+Bi�S41�ҡ�������pC`��Ő�dG��#��g��˦N_:&% uU�>^Xf�P\�}��_v����6OeI����ݧ3F2?G����ޟ6J�T%|��S��C����29�c�Q��պd�a�NO�G�&B+�b���4��ǿ@�[>O�����Mo�~�?���s���3-_��kj#���ϡ� 4_T�7�;�Σ���Y��+���jߧɨ�F�5oqn,���h_�ۻ���=飶#�p���a����U�"?�͍.}���$L�:� �z�x�ı�z�MZ�<!�����j�>�af����UB����2	�iqڥ��J�b�2�qJ|9v*|���J^���8�SD���ɖ0y�%W�,{�f�E�oj��r�.)�m E�Pz�LZ�^����#6ٱ�BQ:)��bu+*T����|7O�Y$ŕZ�nd�.C��m���Mί7�P��v�����ù�ჰ�4�d%����:��}��iP��+b_o*�)���y����Z��!"��c���|T�\9��2��p���i[Ku|�"!@�mAk}���g�}b�G2�8�h��n�s�k[�Ϭ�����&ڭv�j}j$�����^�d�fv�u�+�-m$�7����[��R@��~�k����K����쭀�ҒV@���eY9 Ӝ_ܮ��ǋ���˰e�c���5�&�W*����n��.�گ��K��|$.�5��1�;�҃�y��m������}��S�.����nY��"��ŋ��4�٘e�c�����pai
"m��ۧs7�6n5��]�~�`}�^�T�(r�c��h�=����i�ݷ� �Y_ ���$�K�l��ݣP��Z��X"�d�CO�ܢ�1n�Z��E���S@f�L�|�c��=?�,p��"G�ij,�:���>����N�ˈ	y�E��sd�uC'`�G-1ĒI�+��6�S��/�����ט��l���L{~��	c�@w�!W�7�u:��Ss�*�Ϫ �Eư'��ΘmS�7aW�$ta������
�R�#��?g}'�&��\��~����Kq��}V�2�||�]iP��%�T�Fz7ؒח�LŪ�w�"7�P j�0;�Ʒ�
6�}�{�jc"㨉u}�������r��z��V{�j�Hf�$�r�-e��Y[Dލ��(9��!8�j�%��M�v�ˠ��-k'�?�vJΑsd�
�I��T7����8��頍�#�Vݮ>��"h�gdкK���8n�-L��Y.*�ƅ��'��f�1M��5A8�aF�R�vC�{��-ȉ�Ɨ���i\��ike���.�A5�[����X�+�=f/,A���1����5���CpO�?9=A~Md��%����6�"�:���U1n*�p.[�e�5�q`�l�j跿+L�X�c�y&�*ѷdB��p�H��� �̓�^�y��gn����n��풨7�N� bE��K���]]w���AM�ӗ��#���zs�ܡńdݻ2XT�wR�L֨�����<.�+3���z��O�V�N&�c�f	�W�^�z�Q�yG�Α���+���b��+�`be�L9m
�.���g_�J�;��ş�x�u�YDp�*0������șsF�r������P28�ɪ�,vì��"&Ϗcz�5.����HR����W8�; z.�l]�H;��i�d9�\-�[����*��K���M�h�f�9;	�4���+�95t+�F�ˍ�ip�N(�	��h�����J|FK��mJ���tK5��y�k�s�݃��.�R�0:T����R�6�i;&��P��i���.7����Ƴu���dP�����H��gѾ�j5w����\����2�t���tWWj�k&0?� q�A������`��f5C>��\Ë�YƘk--8�J��tBJt��Ed?�N1"�ġϱZ|Z���@�S�H�d�,�z�?�x��
�~3�I�#I2Y*k��@6�o�o�g/�M��M0<��7���pp��%Fk��t�ħ��=���K��c�7U�L����k��Id��^�i1xz�ޗ�=Re�J�g���f(�����5 JZgO�[�m�_��wJ-�i������x7��u���7N�_��w5�fW9_[v$��K�lK�������C�u?�$G������8b�{|1�y�7Q�3��wU�$�7*��V���95�Y�􎑏���q*v.g"E}ml���m�4W���b�;J ���jo�\��hB0[C\���U�
�2%Z���d�N�E�Yd��e=�ܾ��`�>�M�`$`-�AK�;vW�AYG���RzZ��rN�B�@t��x�`�:T$j�gk�Y�� U�CK]+��'��*;yzEpP�ߖ��./�+Dtv)5㗌�.v�V� �њ��\Úi�m!�n�D��(H�*��iޛ������9uEs�ۤ����@�x��f��όM�ҁ�dwW���7Ȍ���𛹡�em��g\�H�%VRn�$�h6�0�K��������@�v�]
M ���#��h�0�|���w�M�?2�\'_�(ɗr���a�-�[�tO�.$�TR�������ᎀVU[���n��k�"����D����~�g�4��@�t>��v;K��f�� qa�"%��`ט����xhpv��E����+rn��ȅu��<�k�I�9q��o)��X��"��x8ː�f��Sa@�c�ߎ;�[-J���R �ִ�f���H�͘�I������Q�Η�P�]��#h�kP\�]��+�D�ܾ�6P���	�/j�PU0�E����ښ�r'����vqB�����r�u���>Y��c����r�c���B�9<�jh���X�0��;/&����NmjF
�b�g�i��A�T����CÏ'Y --��Q�v.�=��r�5|Ȟc*��H��=��wI��рd�Q���p����&~6�G��3���7�%�jX�qזZW�(�~ɿ@
����FQ��d1���3Ax	)���Aw��v���2���6v������ ��b)�s$�;m1���V�2w?*�{B�#�k2}guD�������;e��ϩ�����[Υ+(�t~=w2�	�v��4����þ�y��&���Z;�-�":�8��5��^�H��U�/��u��0���ɬ�G@Y:{22-�+ڂ��_�`����c�U��*Jm��P�sv��d��\6!��WL&OQ��(���s�?�1�������Āj��A�"���F�gO�O/D�p���_���`��
�G�IH*�
@N~����6�q�(Q�(:J2�=_���y
�z��z��f���Ƒ�F{]�dp���i���R�Y��D%���%]5fGǕ�J�'O�D_�;����ZR�o�mD�������f��[��Г���� Y�+�sC�A!�c�=\H�[��v��� ��YzPۼ����6.����{�HM��Z��U��r<��E�	�-�[��c�k���.�M׻��r���@0�����i�|jG���T�����#����hE1��h���m�<6�>����bӤ��������N/e�O�V�����U!�f��M5��$'�<�*!UNa������n2%��ۀ��c�]ПZ��������C6\�!|4Q�T��u uwF�y0AopV��fr ؤ�������7r��4�]I��6XכAC��N,2B��J������:'L�.�:���d��C*Ɋ�6+�Jg��+Ъ����K�tE�),�趕��D���k�������Dd�}I�D2aG��Q6�r�{󔔘<��U�8ֈ�y�R����YǌbmBS�g���Uѝ�EV�)W��K����+�w�ç2"x;j���t��\
���P���İ{(��'�O�x�88�Ŏ�/�U4�S�ҍ��K�D��T�kݮc��B1l3�bw����mX�k`j+{}j��6N�l��xo��. UB��Z�*ؿlT� !ĆpUC4-��o�u��]N>4'�"	�l�X�V����o���AF�t����:���r�A�W!^c�/�%��Q��<��Fd6
/��GV��6���%�J�p����a�F����E\���:N��Ĕ8#g;"���-@t���2)��P�K <q� um�d��]��=m�0�v/��;l��T�/V@�������h�J|(�Ke8�%�e��yF��B���|��'C� �:>>X_��E�@�#8��!�������j�^Ч��:�����@"��9t�������"8���jq/�ޗa�Tg՘�tZ��bh`k+���+b4Y��2sn4��(%�.�Q�wߘ�)�&����(7�Yml,�l>�?�����r�U,�nh���4Z��9D+t�?��s�
�J[�j���6�)�14U�|�����ޅ��Y`�zW��r
m]͸��\���J�3�&�|�$2)S�]���5U��5_L���Tz��F�JlϮ�۴��Y���q �/�A$�qk�j�aO }���}mDs����3��bgf�R�I���pWؤ�l�A=�^'$���S����}ݤ�lnL�A�.��#WJ�U��+���kC쐮�Z��B�y�cP.��[�?w=EG1^A�ߌ{�Re�wX��z�y��@P�v�1Ei02<���x��o��r��.g�b��L����&pƚ�/�1Fe�4>�2?��<�b�U Ob#������@j�x�6�N�x{�!����(Yr���@%첬
*��H�{&��,�eZ#�1fWG�z1�`f�U��]��L�����n�M�І!�e�����|2x�����ِ�V��O���x�~��E���>؋���헥�+f]>��C޶��Y|�S��f�Z�^�X��WT��'P~�����ɡd�q��X8X"Z���'�d;��,R�����qΗs��z��s�Ԟ��A	D�B9T0�)�F۔0�k��y]�]J��p��at�O�M�ѹM-/s1E��XNʦ�}�5���撪h�
���$e�aW���P݌M�{�I���p���'�=�}UNO�|��E 2w�/i�r�{��\9�z���i9$�!H���k����N}�����;Q u��5##�H�	���鏲���"�Mq�bt����wt��\��Ò����%�����R�SE4ݮ�V�X_	�%6M$>��7�᠒�� �����CB}[kJz<9��IĚ��BL-;�_L����G��q�@���Zn]�堛���v� �P�p�_���V�I��'�U����s�`�����!�=Oɇ3�6�4�?����c�c���8z�^\K'�hxD� �F?���_7֞�	�<j������!�D��*WՉ]2QԴͥ�Gb1oE���|���� }T�c��|�'-�r�\3�������� �5H�bږ@(Y}:@Ĕ}ga7������B���.��Wr'ڎLxM�y����{P���6����.Skq �����1�l�؁qv�V�q�����)[+6���}���n3��h��������R���vH���>�^�]�?S�6���H���U���1N���W֋� �"V����3�?"�����$)}-��lΧT�t5nĆ�:�G�{5V�c��~�#x�v��3���qL�g:�LF^��*Ꝼ�֍<��v�}�Pt�J����8�Z>Fp~��L��XԖ�x����6��� �Ƃ�3ù+���;�P�."�����D�\D]�JM���Fv�mý`�<ٷ�W�QwA=4�G���)��	�s��돘Wv�R;��ϭ�I�����o7�fip�}E�W��~n��-�.W�o���v
�K�0�3��C����o�ȌWr��σ�=+��\�cқ����x�X_ǘ8��&*NQL>�ނ���j�q��Ph ��F��?��Z�r�S���E�ڠ�)3q����d�����a�,���"�?d���~���3F�bT���H�<�B�:��a�2>hd����{q~�͢EL�go�Զ[�z[��8�Z����.tA���� �׻�X6���f��Oح���G��cUm��4LF0��L@�X���|:3�L�L�8��~v �Ӿ3������r���0K	�A�j(�!��������5�h��p�d�� o9��@t���4P�GDb��]�;mc�SX	����м���':s���-ޗ-�8�e�xg��Y<����	��Z�:���q[���+~��-���=�M(�2ĸ�@��x�f�0��>�=ɪ-9�*��Nt���gJ�|������%���]Hp:?��1���$�lq�K%g-��P�>�)B>���'΂�����0�!�l�J������J� &֮,s\�{h��$5.��E�m�V_R���6�hZI��[�ۘ���'k/{!+N��Ks]��s:�
��P�����
��!���yg�	邂JtMj,�\4V�@���H�������&6`݌�F���;�N���P�$c6�4#A/�3ʉ�
W@4��cD�0&��������7x�Žw3�g�ͨ�U�Ra������e�{7M���7��"���?D�<��~(���;G�lW�v���
�T�.2�:ՒEXɞ�{���->j�<�R�J�D��$?��N��c
vQ<j��4�AA_��Q��D=�Oݲbw�R_Ѵ�V@|T�^5�N��?Vj�0{�ʜ�w�	�Nʶi�l9�`ΤYۗ�SH���,�P�N�&�K���@%�M�34. >�P�'�f��O�cDf}������eGIm�A��=.欷C%YW�|d�=D�̿��2A�*�x��Z����)�m��3B�l��W�
|>k֚���F�T@2 �y��=��xp.�X)�tۯٜN! ���hbID����[�OU-$_�l�]�Q�kdz����隃\�#��S��7ׁ�u�n#��Me�
*�m��7���lh���J��@(m�VB6�Z;�"P}��إ���Kq�����*d4 ��I`��Z�b0ܟ�%�Ø~��'_��G�Y�:%�8��]�����$KI<h���it�%[���ZDd;%�K�iʐ���M�@ԃ}��.,�9��:��4O�Q�d��b�>�=��.�r�����z)ok��>�#�^����\��^s0']�$��Hx!��%��u�B�u,���Ȑ�膌{��x���0���)�;A��X�;� u���!WQ+M��xK��=��p�?���
(��od߆�'���FG-W�\#���ŭ����V��s��z���M_��z 9=�ƫ�k���:�2:�fA)��p����3���s�AzA(<�J���7��X:��-��mvy�\'%=��7��tF�)��/�@(�j�	U�Vo%䮓�#A�.�8�߶i��C�А�$�#�㲧��F����{H�	����y���F�'��쭾�5�3�o%��_�U����k>7�if����M삪\�>��<v$@i^yk/����(*�T��7�w���j�:�yR/+��Sej�����`7��Z���'�ÈZb.2�y]�"�z�H���~~�w�0{jDJ)�Q��p�=��0V���~=�I���6~��FpD]���ʺ�mdY[FX;rS�5u�'3�Z$Ct�@	���;�ۏq�����I�~�}2Svtq[-H�2ce����M�k������)�!���Qt$e1~��=�b�h*� uq�>-�^���`��Fp�>����%�'/�9�Ag��/���=��s/9���6���ū]�ﯖ/o�\��o�/���S6���}�A���p��I��A��{��lL���K������0�M�3�CJ�_���r�	��m����ڃP�aD�F���%�a�3���r6�����&�Z~s�$\zÜ�0��"�.�ߒ��}@�=P}~�$:�����~��ˡ!���⎐���K�x}��p�|�~��"Kc����y�
�tFԁ�iA�;�a��������
���T�Q�#��&�����Y���9�bi�:�4V\%�� yH6@�H�#1�~j��������!A�ڿ �T�>� 5�%�@N�ߑ*��8��#�P[�R���r��7��>�\�����t������LAN�d������L]Zjw��y@�V(F�0�9x�Y#o������f:��3~c����ț�@Ҿ��m�hV��8�.�xc�J~FU�/�����,v�N���|M<�R��:�c?M���H
f��q�`��j�˝̀��:3D\�q͚����QL��(�u��bY�q�Eс<;tɢ���l@_ƥ�=�E8�+��6�VN{k��N^)��'��g�:$e\�X(>[I紻��x����B�nix�e|K{=��5� ��spVq��^d_0W��D[�����v��*�����wM3R%���c��nA����!���@6S+���2�����j`ļ���}y�X�� g��Ο{����y�J�s����%��}��`�A���'�/K���I�Po$�8����/�G84�J��tV�v��+lE���R=��6~,�`��~駺��6�7L���e��5!N�.w�s��������UJ��:�a���#���zB�ys�^��6�Ơq\)
U��+�=u�צK��Y8#lNo���[��ǖċ�~�i�!��@��������okB��-t�̬a�s�
ɉ9�|j�IUK<82׏ݒ#P�,��e�7E>�!����}49�{4����7B�[Y9iɃ�\�	 �"\�?�MV�ƾ��-����X�Pb�<�2@c7ŭ�������������T�����A���/��BKU2���J��Il�U\����Rn4v����qr��C�ep�?�b���=��г@h/2�-�]�|O\WT�y�-��R��ƒxͤ�G_��Ves�\T�u�][���DF���_���	[Ԟg�b:���Ą�6�:�)#�V��}��/e�Yc���6Pj�#���Fh�YL���L��(|BbA1;�4�����S&�)&h �kN��l�F��(�h�7�%c��uՖV��Dt�U~V⿫�H�K-����ѽ�f��6�mK���`V�rd�	�vEX���� Ɣek�IƤ�r38l�X���E\Ղż{�kÁk,��م1]�]��Q�.�m�-�ٝ�$�|^RJ^}�E�ԸX�gP��x����������k��'E2�Z+I~#�߸�)�]�}dq1B0�ܙ�v�n��$ ��M���C���F@.+���@E�HӚ��xϴ�&� #�wf��:��*\%As=�+�B��R��7^P�=�D�-�S�J�WxmAuc����,��4]���{&d�j�Qua :�u.��b*,]Ƣ�;Q� n.� ��"�R���`�P��2UdCf{\z� )�� �-��W����A���_���6�O?��L�[p�� ���h��&O�f#��>X{��A����r�i�O4%�vd�]Q��Xn��7���o�AR��q,e�-!d[��'gN����f9�T$��qA�qoL�y�����օ�q�s��.�=e�R��=��N�Ύ�#�o�b(Q 9-i �Ց~U�<�����߳7h\�{�)5�|_dث�^�&ش23��Y�w�~?9��M�j<|������)d�uu����0���4�>6�`	�8i�cUȍ��W�қfa����ǫ�Ҵ���_.R-09L���TP:� ��Rg4РZ=�q���4V�o�T:�K��{7�� c��K�-k�QC�.1s������<��m� ��͛F�*>����)E��nW����|�ܕr{��n�g2�����P�f��ƜY'�3������MyT��/D��9x!NxUÑ�е沮���E��3I˘t�W�q-��=���M���� 2Q7�zL�����ɵ-���?X����8D�B t�mYXVf�e�I�F��O%��5�.2���:�}�} v �,�rh� ��#0�_u�ڧ@Y��媑d�R�A�m5�A������~���/<�j!�팣]��x\��8�~+{�avh�b_����kŠς&��\\����]b,J(�~n5�t��)�;�TOVz���޹f(�q��6��.�'�9��"D��P�CO�g��g�C�ۿ���y`��Җ�"�Ԍ���o�	�Z�DW�>�9��D�1V���T�ʙ�#yC�w�r��L������>iV&�r��oʻ K ��%x-�>B��ɏ<�dũ^�������g��~����*d�������)ns�/���Ƣ�����S��4U@B��SF��Ʈ��
�ʕІ�kU��G<A)����ѽ_�u���C��V�k��}b��q��s)}/�N-.�D`�5���PNR�ؼ�(_.4�`��p'l)��� �
�HO&�����׺k~ˀ���2��[�]�{(��"e;>��A5jp�xm��
=l]����wT�����_L҄�h Ks�ؠ���;�Ũ��=/ӧ1妋9]�-8�����A$�is���?w�*�q�%[<%W]���ߓy����Y�]�Ȓ4{y��K�t���l�N�V]k2_t��"Ly[���3�7ə�t�&�̔Il'�U�ţ#=�4�*X�l��m�����Q{�'3��S�0L�9�'ظdh��Ӧ��%��W�*�Y}��<��q:J`��P�H�j��Ƞ �T����.�H��)���ʒL�Jy*4>�U��O.A.�������^mb9w����#��Vz掭Y3\յ�� x�M��?ܧ�^n��K��9H�`�[,6#�x�vw��߭��i�zx�勎P-2�R�o��(����[��\�8	Ɵ�sE��F��Asm�kˁ:k|x�_�i�G�C���Y�勫��� o��k<-h�\�=jH��O �f�
NVr�����O�ά&�?ip�L�'�|R �;>�1���&w�˄��cL�q�RA���f��+Ո��+�������Q;�m�=����.�1L��j籒j&왋�i�G���)I�1=1�&;S�\$m;��;+ː ����v����ح�L���3��C?�R��ې_��s3��=�!p��J5��~Nۦc���r�[���}��PZV��5q,�>�W����,��xLґs���w}�MfRÁ&N^[S&*�ye���h{5;�'$8[��Ύ��Ȧ��W�eá�Gl�#�:vY�eJ��������uF�%X`,ט����	O�Fy}����Uݬ5��#�-�}�d׸�x�]s���BLf��P+}�E�5��Ei�*Π1��F�֕��#�P�D���,ȗ���ئ�DS���s���#R$��bиI�g��u4�$���U}�����0�	��l~)�|���}{o�p�kE�������� ُ��~��/��sW���ZSS��':z��Ix�m�U`�ȅ�����6Gx͕��䱣W��fk+�pHx�@RN�L��i��z�j�D)�h_��ʩi�ޚ��&%o'C.�ćHWƎ����	�8Z���U�@�uG��,��p���mu�b�:-GH[����F�?�hA[��ݛ��V@���vG]�&�*��3ZK,6�.P-Ep�J����NrG�/��i9��*ɒ+�ʿ���h��<S��T5vp;�ht���� ]�����0S��}����0�gY��Qs��̡�^�J��w"���Zȝ[��Cr������f��`цkP%�A�S���,r_`�"��Cz�u�b���v� +Ӷk�N����=E�͚�⃾=�@k��`D�E�v������9���@0��:�A[I��pD���ڿJ�[9�cO�U��b�9��ƃ1��)Lto�x�����T�sV�S�Y��T��
���uߎ�|V;D8��و����+����q!��>�ġ�*��wʼ�JL��@��%�� ��;υ�o #s��$5K/��gxAl-��	�%���P��Y���J�0�fBW�3*������n�F{��|4��$�nps���#B�۬Ov)���r�|��� ��~��m�;L�]��Yc�� ��g��<�͛F��}��/�� hc�N�n��r�%����J�0������شegqe�ߍ��jG6��Ba�q��e�1m�t=3(�wz���l�=p���X^�{��� +�Z�`�.G{p���p唨[�Gi���R0,� c��ggsn���zw�����E�kB G�
T�����h��GK��]�8�D��Y��k���y�W�&C�_8����6V^�V��g��=�0rx$�� TԦ���-h��������� }���	KA��D����+��})X�
�����p�T%|�v�'L� �����1F��\=AA��J�b��[��2�v\ϴ�:u�u�]�>�b�?�@��S4꧰@G�n��oL��<�a�����iK��?v���<e(&8��(��j��*����2�%�1���s@�jr�T��L<�'_�Y�4�H'�2������k�zj*�,G��{ܞ��" �˔�3����hVu���`.)�![7eݦyC<�{�5YJ�?;q�'�{~w3�Mc�|��t�h�L�U��Cf^2sŻ6\����g�0��Ͼ�o>J�k����k� �&��!;`�r��9{o�x`y�_c��}JkHc��r��ƍ^�rq�>f�/z��'Pe�Wwz����Q��?��<���������"�+<���u�JV�^���1A��e��$����\�!�%p�}�1m,du`�!bS��s'�����e
�_q�S(�mb_�ub��
�v�!�g��6
71p>V��K����0��.�I7��A�m'��i0�R��U 6�+���=�U^r����VkYn�i��.0D�A�J��"�0�C��/�o�e/5�=nh�/��������%����uӐ�(���� ����.�맳��)��П_ҋ�VDIa_$-�{TX���Fv���������F����;�e����h�&ȭ�;vs�a��d1�{���[=�?�4/%03l�j$������|:�ۀaLk�Q=&�������ojfIQ���mĉ��lT�"í�E/���SǬ�qJ��KTp~��ݤ��Sc��:�#�g�$�
\�l.ڊm?�7#�s<���L��O��qx_a����jm KuS��a{��y�r8ȅZ���./�%�J�Y�bC6[!p/_�q�D����O���O�;ց>�r���糜V�b؍�,��������Η�K7����4���#�W�z!Hj+��Z�m�Cg�fD	v�(��_sZD�>���tW���A��Ј�;<�����荗K��yu�K�_��{�Ƙ7��Gw`O=>ޥ�@�2v�$�q���ᵱ݆4��'�TXj�D ���t�+�X7>�h]`=���r�L���/ۢ�ā5�MUG6o�*��9�I'Z^JU֑�27�1���E����\��E��խ��/�t}	�r�ˊ#B��&Y��;�D�(slN1���6�@�il�^��ӯh� ��3�[���;��
v������%L���K�!�z�ҹb��!82�4/��j���+���58]r���=u3sz۝#=�JD�4M<s6#-�|�<�L�����󬬜>g�>+�b��c뢊	�v���Z�]
ݶjE���|4�*�i����DYy�����Ie���I7t"џ�o]s����Y�֏�l1q*��Ȉ2�?/�ǙV�ih0����e�8'�R{���d�l�<�UJ���g�D%�O�b8O��k�zIX����\r
[��軧�!�,���Y���Xv�p���ѐ�%��m��k�����=#M	��\w;�!1� �>
�2�,<q��Y*w>{\\j~���b��*�T����szD�0��B��!V|)|\���oI��~8]��Ģ��ħ��,j&}_6zL�ڍ䒋{3ĺ�4*;�2^��>T�`����[!V�4��!6:��z۸j��
��H����;�)����E����[N$��4��U�����.7�o�dܨ� ��E�Z�og�z's�·
��A�$ky�YXw�T^{���ا�Gs1��g���(N��#r.������Ds�����~���	��Ȫ�&�гг�G]#qVG..Cd�`R����mԲ�un�����97m"2n)�rv��t��VE�7��2�\�;0��M���x��̵��8���ΙC�����TH��yɾ@@8*c#הR3?@Z��E����qף�9�a'���Z��W�� �P�g�}��(�"b���;vJ/��)���X�-�H�_F�,p��I�&:�
X�WI�u����-f��c�	��=�X��i�&Zڋ��l%��#E��F�R��x��{v}��Q�+c�]�B��-c]�4��إ@Ϗ�mr|���^՚�F���Z���&Ҩ���߽���5zܰc$��q6�s�Kq�i2�ס�8S� �3���a�HBl%�\�v�K�[�sd&&l-z&����:;m��\�~�~�7u�i�Dd�(�j�:WW������z�n�NS	q��_&h;�2�9\Ms��m|�j�����'���D�̥���hg4s���Ïe6�V�q�����ϯ=͝������r?�$yŖJe,I#��ו���Xcf]}H����.-��J~g����1���#��MDsl�]�IE��uB���́�43u�>�L2
x�v�	<.·!�N<� ���-�B�v�8� ���9W}��h"j�<g�_���E��sW��*p�4�w�Ɯ���C�����éZP(�-$�w䬲y��ݮn��D��Ɉ?6��AǶ�Q~F}
$�!5#�)?M9;��|�<�S��(�X�:� ��Bo��;W���j9Svќ;��w!܅Ȣ���W�^��j�K��)
O�-�򬙞R��P�Vtb���R|�y^���69L`�l�[��)��q[�ƫZ��cU��95�5{V�	E��j]�M�M���L..�W�6s��Ҕ�=��lJ���nA�q!���;���N�� p7n��"�I�w��
G>��6-����E��u�w����`]/����5�����kn����]EQ=���d���������LUpk�
�xQ��Kr,�T9^�����oL��� �?ٓBAc�"؛
��1�p��X�aJ��W�0�ϗH<��)�8>F.w2V�[����N�XĹ�qw������@2
qZ�Z�n&���!~D��{�S26��#)1��Y�ݨ�����O�R ��$սDD������~�,�	�%�%wۖC�!_VDb��xơ�䳤������ki��p���[ޞd�?>m�P}���b7|B��毕�uR��S-A�#~���Z�ݓo���e�3�Ȋ�,u�fH-9���O:�?��@����� ��*p[���Ғ�Ӊ��js����1C�VT
�C�Pv0�svԊN*ބaŧ9?�i���KV�	�T��+���NZ���Kf�%��'��౯�w�1C�����G^�����`!ǌ�B�3b�.j���"[7E�Ǹl�'��[U:�ѣ����d6���.],G3+T9���S�;dyk9|�CnIhe�~r��������:�R�n�7��c(����#��]ͩ]i�rWS>\�,Ӎƚ�o!5Q$�u��Yt\h)��+�b�Epq�]Z9Ps�q���o�s'|n!�}��z#�nK��gSY���ǥ`�("�u����S�<͔��`�tN�rqp�]���/�xɥ =�����CXT���Q�(:yU��mH˪'��J2˰�	u �̓d8]%�P3N�"�M��=*���i��#�\�?H7v3r���|P,@^��.�,{~�M{)�ץ�����;���#��tn�0>^V����59�#�;�2/
���Ĳ�׌Mu�?����<NA��:.�|�T�eP�.�c���YK��^W�� F��1_����B�L�:t$a�n�T����"���O�n�s���Lg�jW.d͵�H���_��pq.�u���Jq������Π=$$z9���ԓ�E�+I��Nl_mW�To�毻Fg�ߴ5O/F�h>�?k	d�ȴ)��^P���[�M�
�yܬ7��z�^��G�g	X�֛j��' ��ж�j�Pp��P@�f��2_�K��EԲ��1K�Ve����}�����.o����M�ٙp�t �8��Ŋ�F�Zv(V�&X���������m򔂩��O�08i��߰�R��:oЭ�6�j<J��M���/�5<���>���,7��:�UE��;*1��i���-�F
D��nz��=��xL��T�@F�}��ܜ��'��0?!��
�M�r��B||�u/B��	�؄�;��܇�k>n��a�e�@	�haSg:���x�:�������#V�Y��u��vyjGB�>:�:5{U]�n%�:��<�!�)�W�M��ؑ�ț��7�Φ@JS��4�:Ȍ�OO��fg�q���~��͞�����Z�a�Q�۔>����o��E�suD�� �[��Ҥ=��vb^��8�X���ח�o��]���3�P��5���} Eͬ��;�ԟ#O��eV�GlO�T���~3]M�`��2.2������l�}H�kz%}]R�5ף1e׵�����D� �lj�I��h����5	�[Ŧ+E�14�\���U�6
N�H�S��OC3�ӹ�	�W?П�s0:��t�ȣ�ْ��5�<��M�̲�#O�E��"�C�*4���Ӷ+��{|��VP&�J�IS��u����oh��5��%62�bF6�b2Z]o�}�N���E5ƥ.��+�n��
��������#�z��43�IZk;�)��$���E7��D��ކ�j����s�B������O ��zZ��L[^����Ղ��!ۇa�ڂr��]�mCͨ�
�vD
�$ ��#�8v!]�AѶ�r���iM��H��F����yC��~Ӱr��=@١���O�H�Q�a�q���; �8�iT�&X	��;p�$爕�W�ו��f���$��`�xA>����")��|;�"H����?ӣ��ƹ��ޞ�Y���6x{��/G����l ���44�ý����RS�_��V���W���j���!����+"��AdpI�9A�b/��L���b7��8M$��}S�:V�Z�$���G	pu^ؒ���O%�櫛>[�Ix�?���C���L̲�� R ��_C�7�v�-��~Z�í�JV!��C��2d̮�ƾ��]6��4�GR���Y�
����=�O�Z邈�0��:�b;�{lm$ѕi�\RP�����o�1:���|��j
I�ۼ��#�s��)�!bա���� ��@��l���U(X4�dbl���ߒE���'�c�4:�\VNl�}�]�O�ƪ�f_�%���ؼ�~xL��T���g�Xu�]����r��B>���%y�v/�8o�qkQr�h�c�JJM�o�>LEJ�:H ��|���.{�E��w��Q��9�I� J���Iv���(F���]�h�l�5h�p�)-�/c�bk��.B���ˮ}d�1c�pz���Ç���+@�|�Ta��=��B�l�܂�x�撊�ᚅN7��""�k锪dW��[a��Asؔa��H�a�H����d�#�=
�c�a$�~�.p��u3��߽=f�g��t�|C�V�L�G�ԼΩ�q�k�E�(���ںN�z�ƎZ��B$E����%S"������YaϚHV^c���R;��L��嗞�gA�BG�r�OdC:���)':"T�7d�'w�q�֦ڲ��~ny�/+UͿ����\H^�Pd�X��of(@fh��B��ʮW�24�-�@�8���v	�%����d���w �4�B	�d`=�ʫ��8��M k��}����Q���`+j}�G�˷��H!����q���m����R�L� ����b?�O<H.i��� |S�����QVÙ�����OiP���>8e�j�	���S�9��u����0�re}�ist��D��s6U�㭧>D�on��GV=�GnE
���/UN�����5kb�@�$ڭ �:������I�h��v�K���6��K&C	+1�5�u�Ҷ�/�<D��W#���d��tן�-�+���e� ��*��Q�ܿ�h� "�hl%�s{��
����T�mШ0�2OG2���Eٍ8��E�W�ʎ�cz�w�R�%�Amж���Eʣ�ře*�2Y��������HK� �C>b�;-�VAu�:R	��d��c�M�����sD��D�FKR�����k�MOc�ED&N������k;����P8���N�� ^\6��Aveh��N���Z��yd>m�`�2�ǒ$���4X*���e��z���-B۹�#��C��d�(�m}����)OÊ8��w#��|`��1v@51f�F�����\$!x��u�鯀kb�w��{��7�JAr��y�_
u�&߿L˿����,o��|:�t��\���L�]�.M��*�8|ǆ
҇?�N�x�[W�>������Pp%wmd�Z`�p���H2I�r�|"6{�z�*�շ�M �&�/�z}��dsY�L����e���7����(b��d;$���x�w�k5r�m_ �!���^�ּ�q��?��屋��>+䇗���Y����lCk^�'�%� �Hh� U"T7�W�+�\ޞ����n}�LU���a�>j��r_�PS���\���P����?�?U�[1��a��A�t��F����'�92���^�"7و�8��f�z�H��Җ"�EČ�f��a\=��1P�*�+��.6.��Oj���m��̒�h��\�������_%Z����õ��H��YZ�a`�q�>I�����x��>�3��K=��é�&�UIO���Y�uz�)�"�����"x2+�-���N-Z�pӞ��i��qo-�:z���{U�.ͣdP4q۵\r7�>��*F��*�Sy��0�ܷ7.ٖ���]Q&/+��8�t�;	]�_��1�H�}���ý���l�H'����=c�(�E�Gm��nz��_�W�Ė�y�!]m��a#��oK�EVK2�#����y*�Y�7{C-�����~�xF�	�n2��
��f�V��d<P�dw��H萦��ϋq�i)�yw�#�B��z���~�=!�vW ���Ι1ef��7q��Hۆ�!��jME��9q���8)j�����o� �q�M�U��OH|�/�u��r�����'�	"�3WR�մ�/vг�҉w5.�0���D^:`O�r�*XR��Q�bm7N��H7\��q[���dj�L�#E��*~u\NP�wk Z۵T�ܴP�2��-���Q5<R�qK������e\y��_��}��A�w�E(��f{mw���S�^��}��v��%��d���@ԕ�*߱\}����|p�s��æ���T��8���G�c���mm��"�`��E�"@o���Gu���\��C�V���?����A��|��~�0l]�|�n��,�O��n�Qrn�GHt��:u���jh�`�|�M�i�U(�o/�K���T-�#�������[
<�~�B��vZy�8�.#`��扒�.%�D9�&��|�����B�X_��X�u �k�TN��j�+�/��?_2Ak���ߕI�BK۩��-�t�8�W^'�;G��i�BՀ`�2�`�>蕷^̞�u��R��0�`�lû�ɹ�Fj�#x���o5�Y�����������4BZ6��Ti�I{W.��3���~傭W,W\��e�T��(�b��3����_��$7�ݲ�5�+K�t�;m\zE� ��\��> Y���خ��lBF}���!��/i�[�dD�;bm �4��6�-��eI�.}�6�s�Ź(�DW�[*&E�'�TW�.f�]�g�i���̈́�J��H_94�4�����_���i�(׷�!�$��U���[��a.qv����3��������Ձ�*�9$M��	�3f�wo�'<-���6���^�F��m�Ł�뼂v�Q���G�M�Iܲ�j�4\������{�*���	G��R�׹A'z&����G�~aX+�(�ʮ�(e��,��uq���ਘ7{+�E�����,߷<�J�꫉�(j�"�EO����zR��.3��	�#c$��r�
^�T+8Y9:��J�??�VO��-
̭����esVaRhz����PQ��:�I���6��-��@~�kxq&��O��yةtm}�i[�>��{�_(,�O��9l7��.Ȅs�����������ό�s6v���������
�>��ib;������11i����RH�,u$_4*e)~��o"ҧ�@�J�M^X��7h46 �@���������Ij�	7����9��>�뼸�F�
�*Z�c���ǧe��[3��#��_]�O��^O��S����-32L��GƇh��Z$j�{��1�U���B���6:\xw֡�4Lf U���a V�n��\7T��ci��ܺ�is(��3��q^����س��J/e���D��I��:�>Q�a�l�}\m��-9:)L7w~�����/{n[J��@'k>	l'�gÜs�~�V�E��(�7ɿn\�gM�(�7���Q�4:#�@)4T��`zu\1J��x�?��4�ݔ�{�c�j�y��ug�<�1֙�\�-�NE�7��/N�=@�ϋ?����!9���v[���	X�z`/*�����5���������fPH6SL���[�[��7#ޢjy����ҳ1���"�&\�(z{ ����'"R���X � �Y�yGb_m��to����x���sǋ�l̸xxUA(sl��_iY���Ҋ�M�C�2ß�,�cii�FĂN+��M�������` ��
	��X���U�;ʿM@˚���$B2�~5e�I�%�x�����wk&��i��t��[�f�-���s�:��6��J�Y��*m�4�1�����V�����4wc �V�1��j\������_f68�����7���@��h(?x��@�~��t ���u�pƣ��-ln,P���C4����0ʱDj}��2Ԗ[I�(����Ѭv3��'y�%"$�]����R����C+@\& ��}�O�b�2@�*�Yxl�:�1�&�i+�_:K
TU��z,x,=vI����}�b{XS�L\X�'߰��^�f������]0K%a	�n�I�}qa��c�~�*���"
op���^E��wO�����}tĽ���S�2��o���ԗ����n�Ή�&�jƖ'<%T��J]bs��-�PYT�48n����A2]0���q�z�=~�<����%6�1z��Ð�~;'B5cdf0#S� �'�����ɝ�'�Jʠ�P�cnЉ�C� ��;2[��IC�G�f����<gB4�X��_�����-�͑�Q�4������pCG� G��H��%3{x����P��<��ݣ� 5K¹������C� aU�J�VڎW��p����Ģ�tу�TS�0��S�K�Y#$#��Hbך�8�1�n;����N�qMqrw���w W�.B2�aEG�?h
�l�S���$�4_v��D
�%�D�V'��Ω0�Z�Tչuo��WJ#R��%�&������yw�WK�e���i�{S�	Vr�7+��ӵ;��+�����w�q6)�5�-g�|<����ڑ�Pj���u���̈́$��~�@8/�`Ea'�@?%-�OR`1�f����eBb�5O��n����F���-@��pTMh���R�Q�Q�ƻ̦������"B8w/��wI�h���}<�K����q�O�W�*w�Z�s]���U.���>�J����P��Bo�AS^�Tr�_��H�nsm�����+��6�;�:��:��,T����E��F׾)TV�� 8��"�q��;�R��D�6���f"�h�q�+����wq�%ڟ��E�㓔��J���9��VG���[�M��F$8���%�Z뛇��i�ߡ��s�T����6ն%�$����w���ī�RHyt����U�'��i�ɹ���"��G�^�ʷ��C<�/�~���s��2�X\�r���THp���t����,`P����(�����Dz��5�/X��+���^ϖ�q�<���*�Z)���͒�k�_��*��_M!Y�f*�
?���J/�<>U��kX�?n�����jjiL[��@2j��������Xb��%q���\Ql��fͱ���a�_���&��T?�i��(�X��J�."i��p�H��\߁<z�3�9R& עj��ڿ�)<��H>�m���XĶ��e���gx3�hnQ��I��e{��k���1��'��w!���G�I�ԟP��l�J��T�.(OPwvA��+���-,��wUr���9�w��Sj�:��� �qޑ=% ��{�GF~�@�-��k�p����Bȹ2.�rXϘʕ/�#�o�C�T{�^%��/ǔ�������i6���b�>�g%�n��b������0�ϰ�����P�L:�����]�y9�<1������R���gh���[s��qU�q,�.B P.�,�Ђ +�
�!���W�T�	��˻�¶C�'N�P�?�4ӏ	6���!���u˹3�dZz�-��B����\�ہ�7������{qd��x�j[�GL��wU�7�{;!����.�h�CT)P>�i&��v�?�-��#�s\��ckT��*�a_��=7i ^�M�S��y ����ua6B4%��+Ͽ�H��<���1"��>~����b�lXE�-̲ٗ�G�n��К ����bLݬ������O�[�0_�G]��qդ��Z������d����V<�#��'~_�Ω?���
�8>r�����7s-xE�9CI����U�����v�;8;H��@�(��ySW�p�M��:g��+����Z&2a��Q����J�J�����y�����t �RN)��v���U�	����P_
�<��np��*zD��_u!�z\)PӤW����x�s�t\�ě��vj�-�|�����8т�T�\�K�~�����Za�-��/I�O>�Ǩӭn���7D������3���RF�,s*���J`��� ����c�l w'8_�|i�(���� �<L;���S�F�1��P�k�I#��B�Nvd�0= &^{v�u{L�����⋭ ��=Fb�������J_��Rt�z�������;�n��n'�]�%֫�xRl2���_���]Fa�d~�t���<���2r�Nv�pf*6P0k��G5{�����^�؂	G3%��u��3ǯ>��ſ����|�	H��͎Z�.o�^���3®�7�~�rz�:Qq
Q����p�Y�D���6��%V*fra�Ѽ�S�BP�����l%����&~B�g$��C̓o0}D#8�<�72]
gW�T%��s?P�팈�P$u�Cg�8L8�N~q�dA��G%�g�4���L��\�ulOj~�r����J��zࡆ2,I3&QG�G�=�eUc������	`x�R2럚��j˷��@o�A��D��]��9��Z	�]�G�g������(F��
	p]=S�����^����X��n\-?��<hM��]�q9�s*Q�?��95BvO𠦟O����JBZ�U	tsu����v���ɜߞ��ŝ��QI-�8�=����?��)� E+6s#;Fܹȉ?ʞ<Yk��qu�g���і���<@�0�&Z��}��|������� &����Z�OV���Z)�<�0º����!�f�\�#�lfr,6��E��BF�����\B�^���m�`����J�O��Y�.��M=���d��@ɓ�lW8���A��/�!@�馁�ů��dE`3�AK�=�t��g�+9���Z@S�n����wF��3���N.�]V���8f>�u��k1=�?����܏d��#�����>�t0.ͧ�#�8X,3`�� =�Ϡ�&���D�����T�(����899#��RR4U��b�P�8f+�o�w�j�����T��e���͠�������0�%̥��V�^aA� ��%	�Y>��E�7A��zb�S.�K;�*��dnEcO��(B��t�\���`D;AԪ�Y�d�$�q�=#���e��q��i�����S���w��HJ����wB��
�dC$�xV�1fj:�x�h.�_A_��B���N
(�������H����s�c���@^�V;4��*�,�T���\�JV��PW;���tri�����"��^^^�	�A8*%á1KlWx�>�V^,=���}J:,��vv�5����[G����2(��̵~�넹y�(Z�&��+�C�z�j�T����	���{2��]!�"Y�k"E�%h{��z,�ԪӀw��j"��T'�/��9�]4����,�%��3��y<%��G��<CZ��8�l��7��MU+��~f�~�gm=Sm�_��u���Ǡ�R�� �W*|J�"[�Y<��FgV�����e�(f�)�."&�aO�;	�������į�}���O0�3lB$<� ��"���W�jv.K�Lxm;*�O�pL�q�Lq�Y�Mf�删:��,��o�E�W׿[�%X$�A���o�H������"I�n���A��{�W0�wʒ��m]^�O�Q)Lz����lS	G���;JQ�v(�ܯ�(e�;�E���˰�qD%]�����ߌ
5�C�ZR7ޯ����+�>����!>� �,����W�QiR"�"�2����c+�%�%<�� 0��7OR?��S��MMt�����(��⽀� O��c���	�U�]B>����J���r X���9�8VD�������������嚾�L��F�Ol8�qQzQ�IzGɩ��WF�l84��4U�
��u;�J�q�ȅ�dRڠ��q"�IÁ��S�f��J%ݱĢ���h��b-�<W��*d��K�x�<yE�b��I�_b���
����eod�������":bq��S+em�b�ߔ��E�2]�ks� i:I��Z��:��C�Vqw�a�7Y�X��E�V�Ь�<x�};<����K��Y��ߨ��%#<�L��Ґ���j�^r��I�'���D��J�Y�2N10t��1d�1CE�����u�_����n�ֹ�֞��<-�?���x{#oo>bf:�+��7����u���) ���h���D�س	|��NYګ�(.�Sw�ž��h<:a�0��e
����u��0�T=���|���Ӭ�F�����06��|˶����w�2(�4J=�I���C��I��6a^S�iZ	`��rpe�X��u�!l�5���	��n���%�}�B���uZ��^�y��4�7?1rx�!@c��������%E�-��O���&����A��*D��j�3��g��j�$)�1i/~���i^�J���=J<*��{ei�P5ƿ��qk1G=W����/
Fd�^u���:�_��'�q���+6�מk���u"f(;�W��.�9�9���,��1ۘ��*��J+m}G`&���`���g�Xy2���@��?�5����3�Kn�"��_
S���c�Ϣ�I��r��}-���.���k#��h�P(��/Kذ�Et�b��T�|";�l���QNR�h�#���{�0�����������Y��j��Cѯ\V$mqJ�;T��Z���S�(1i���[5-{��Ȱ^)p�������TD9P�����nC��Y�{��9�*c�%&������COu9���:W������y�K���-��e�v4�C�#�P��)�>����5	!�.x�DI������r���	8��u�G�ݚ(�����BJQ:U��x�D�D�~f�c���7����������5�:��D�Yɠ\F��2&�P:t�!u�L����z�����b�w0������Ȩ�8N���f}U�����`�q�0��<�C�燑���m�!�d��������
c�D#���OEL$���)5�jU���/����?κ}�� x�Mqٺ�p�g��:8;�'������0�����u�B�0���p�}Kl�7�	#^�6���cO؎sQ�)�=������c�MΝ]�\�oPW��Z��.��:n�G�+�X����+}%w�\ lf�}'OY����zk�VMMZ��*Y]$*�rd��4���-FS����A>�����M}�T����Z� Ɇ���\���G,m�;e�,���}&��,+�N�­t�D�� Og��Q��^�i���5D�����;yp�	w�,��VW�K�I@�H[S��zg���6���wLw��a���|�H�~�3�5,p%B���� w�s��"S��[��T)�6��*C1+�It�&�ݷ�h
��b��kN�!f�A�n&K�7گ�G�|�(���)ܭ65�`V���T�aY�z���˰Y�I`��Y�1��������l����4|�eL^z}-u��$��n�2N*��9.������cG�5ЉA�k����,Q�~pb��7'��k�J�uH���)~����Yf�e�v�rP{e�卐[�@�hv6v�z���i��[0lM��&fb�fq��u�G1�F�b�[�	���N�1Z�FMS�̥B���~B�����B�g�%:m�էeԁ����, u-�l�K�YC�b�P:^�/'�XKԖ�W�5��Y��.i��L��@�}RI�m,�?��y$Z�ր���x��^��VDԴ,dm�LZ���2.��ub�,..d�`�%����!6�x��rϟ0em�������M}��}�Sf$k���;=pKu��_j�X��eo}8X��t�&�I�U[�P������wGc!����]��@]ݚ�v����ӝ�pl_����6��9qV�V���xX):�Mȏcg�]'TI���wCha��M�(��՟�cH�#�U��?.t���!��LD����7�."A������N�p]�+J������_J`
�'/�}���ʊ�֯K�~K��:1�m=�^ ��o����c�&�0K�;ٽ4�fv�W]A����� c��L��Q�B�q�����'�քۺ/��fFl]�r����V��EG�4a�@Tz7�z Ā֚��f��"��I���Gh�O��ܖ�3��ax�;�'�r6}�z_��*9F�z���#�l"������m���]T�d'9S�@K�'bˁ��ʰL�,�rO����{ͪt
o�ż���`���G��z��}�Us]����c�0鬖�=������;���;�q8�	����hO���"�z��p� F�~�����t �ג��آ�8y31�Yw�5�C �@](D$�:E�-��<u\�ۄ�ϑ% ��:��0�XG t8w5�kHj�v�b�y 8�����3}��U��Z���k�=65���Jc����{�9Ey�F��Xk�`>h��yB��	E�����&����o�Fa.zr���[pq�'�M�Y=��x�y�]���W�פ�.��k����v]|�ޒ������n�:��R�^�#
sD�E�0�~��c���V.$u�c���چoO(��C�k��dX&W'�e���}jq�М���$qX�xNK.�����$GFTZn+Nu�$�
�u�tG��,i�H�Bg��
�>�Z\�ں��:׾��@�A�면	4���ຜ�z�~#����C��CR�~D� ����&�=	�(/r	���K�B`���5��+��64�S�oU�T���ϊ�ej��YqǤ6�d�.<&���z�E���&�;jmnl���2�����bc3��SH�7`<}�O�����MG�Wۃ�)׀�"�a|�P�x˃������]���NF��IB��v��U]�����ny~Z��V%<]�w P���Y���y-�r�C�lm�V�)m/
�@`�cݟm��t�	lI��>�|�*�y�ns"0#Ex`e�x�a���[B� ��0v�k��b��xG��\�~�I�p(Sz�'��d�$���q�#�P���^��S��<�k�˂��|t=�(��*N ���7�#��02�4H���2`'�̏�-��
���^�ӛ-˨ٜʓ^_�B����~�/y�YR��ͅ]��N�	�r�˚�O¦��:����{P�o�胍�9���{��^V�\@�^ ��A3�V����	G`��c�Ɲ�?Il�7##�����\(���,���Y�lr)�``m֙��!����l��@B$R�~˧�*�P��sI@}�	x����3Ў������0��g�~9��}L�be��K5T��k�P�g�L�c�݁�ݮ���&M �=J�'��9@������[��6�gi$/gy�g�J��B#Y_X�Θ��lvP���&?Α�+@����2Yo���8,��b&+xS��K��m�fj��9-���������Wt�Ld�Z{@���Ʉ����my�	��D�66_p,܄_v� ���um�� �� \�d&Q�1qt{�p	�5!��0Iڡ[� w6��4H��_�M�m��͗��Ȑ�y��ɓr�y>�&��������,Hj�����A������T�����:���Z\�P��W��xo�{WQ������&���W�Jɘm��P������f-�_B-K7���{A�"Bթ��f%v4Mu}�@�版��	&c�A�����'\��ԙ���wJr����'c��E�����.I��'��)J�<eJ=5���{�n�$�=��Z]d!/w�|"�@��d�;�{��}ª#>�� ��)�ݐ�&(
� _��}�r׀����gXV�=]��/��EA���#d]�pU����A�6���+g�1^�ǋ�{�װ6���KJE�[ԙ��0�]��q�4�B�Kc���N�lC�ŧ����4�*����Š���La\�N�?B[I�N������r�m�_���>X#���HSN)�)�����Eޔb�0^��5kG���)�TKwA�;vq�k���IeCE�g�L!�ɦ���}����C*<i���S)�b�ķClD��WV�{�?eX�1'h��Û1��3T�����,Yo�!��Ze�.$LJZAW�.�Ŀ�0Do�=>��׮�(R'"�EA:3��^�2��a���Ϋm;�/&�4_�kX�{�j4�c��S���Te���´��$�����q^�Vm�P�q����7B��JI�Õ{��vH�Y7�������(�6�7,Ԟv����	��{u���(:�v�I��>Gi��렧D9Ԧ�b��ǭ^m%lB�ٍLX�	}2�u�Z$U�N�~4����l۽�d� ��=�ݰT*��8��J[��EP.q��k=f�ܰ�&z9>�?����U��2����Ԁi������s�	�V��Ոr��f���n�����9Ji���؞r��mQ'���f��޶dy1B��?�9��ʕʫ�����m�L&>Ң�P'W���@+T�ׅ��~��Q+�)���vn����@������i�)��M҃,|g��5��F�$��0��ee-#�y)�lfY8J�˛)�����5׽�W\ZX�S��j�aXb,M��5O���m�6���rCB�̟�t��<�'O�X�r�d�{�>>\�`�ά�Oȫe(xk�߰�*1�%��&�ѓ�6bF�����H�9��o�2��z�]O��S��U^H<��f�)Pz��'��b߉�͙���a�ӈ���U;�J�^w�1�H�EU���~q�t8g,�d9+�,�X���l��Ŋ���40ٖJ�=�}��$S���.{�Q��fI�3�<ϰ\%�'��/�*�W�F�5\}�9��-��&�؍qR�eA�70���6��
>��eE���#��R������f`~��6�=o4�8�M@����<S�Q�3P-�������I��c��EY�gN3z>����	�*��Q�m���ǭ�0��aA녹V�*b�v�}A(�0�Tg��'ў��5?��m3s�[n�=@�(mz���H]p��I샴�!{�ċD� �z�/�0 ����*?�I�bC� _�oh��2���u�gd�!�º���'���K똊��"Q��^������TG&~�^�.&bܦ�C�$�`�q$8�&��`��Km�LD����Y}p<��i@OVU��k����M�B:v�����W��/7�DC�#��fJ���m�7�W垩3�}]�b[�)�'��b�(ƒ+㘭סɆ"��R?e�>Q�|<�]Q�w(��]3ٞ(�e�9-��e���W\~�s�$�Z������_Q<k�#�H�А�/�.�m�NB2�\
i�t0ULTk�ѭmĴ��g�$�Q'L�2�b��K7��_�N�Dj}���2�z�c��6g��-sF����n�����Sr?zb	~�p�����ck�Ѯ�Ot�@:A�2�Ԕx *h��8,��XhT�D)c�a(OPs/�Ď�۳Y53i��S���8ۀ%�=�G��K��r�jb%��^�����;N:�k�;����2�w�Z�[k��F�/L��A�\A�)0��o�Q�6��{>|y�2�rc���GD��{;��;PD�����G�wZ�,u�@�!ؠ�#Ǖ:P��c�������s�NR��͵����j��n�"{2Z��Y:�n�Eb��*�
;b�����|���V��C���3�F�����%`�R���I�2;>u��3��J9��3�{�c��*���3[U'(NU"�E�a�����E��ؤ(�(#3i{l2��ų�QD(֠P�,�v�1p5��$�*�"r���%i�����_&�~_� E�[�zZ+����5���í�
MC�Ҡ��y�-*��D�-��ĜZ�;'g�#�'��$R�f�1p�^���Ʒµ�\?@��t�R����f���}q����T�F��k9i�(c���ؓ��?6��M�@�೥��o��Hn4�L$�F$��lR�>j�o��C�?��M�j���Ɩ��X����U��[��+#k��F��&޾q8w�'*QH�"8j
�3Ǻ���n�%̴�߂ቁ�(�����L��q��®0��X�f#ݘ@TmCT�g}�3�Y�]3R�9rH���k�K��Kh8�:?�L���`���#��T&�9�/D@�`Բ���_����3�������d)?�v�^+�z���;7�ӑ�aP��i b�������	HEdNǌ�y�i(�d
P��fT�l� ��Xn�ޞj
d����V�1���P�۵6.�3�
U����1��/5|���B$�@z�_j�H{��$�HS|U��Ǯ\T�27(�;�EkM�ՙ=��&u4| �>Vi>:{�L�J�׳/NS����Fų�����qv����g޷	~�Z<t�s����gRS3W�+˒歐bP�_)��IM��WSR
�6~�2V�PQ�	x�b��A�(W�=֥�J��~��Yꥎԉ�O��Q��HQ1�%un�ׄ!P�lA�޿��j�X��F@�����r�R��!�4�^y� o�C�4nq��^#�n_���\V9�	F�h��*�_t{��wJ����kk��|����O�"��6Al��0�R���B���a�S��Sjs��f��9���#Xޗ
Yj��y�x���TP� ��I��I�N}m�d�Ǫ]�b7�$���M�=��.�չ�J���/�γXU�v@��wa1�MXYL�����`�x�-@��/:�-7֥q�#�!��֩��6��B{�6(� ����\��/9d�k�������u�un9��^����-jFOӍ�I��o��x���NN�J���Q�&�J��� h��\fw�6��C�}�׼;�k�~_ZP���/ǐj��p�/��T��Guc�\C�:+��!6,�7�fZ��c�?g���|3M�LKO�mZ�_�vA��S��btg9�N���h��@�w��e��V�S�g�8.��<j��?�^ ��jTz�sY�נS�Z@��%��k� �q����[�&��W\�u��|�T�s��S͙����w�aMQ]t2E��fV���f8&aVT����5�x�lޖ�@���I�@��w�p�J�:>O|�!Ii1��M`4����5E��,�����;����,����9���,~=�=��o�Q�zv�-x�Hp����N��#��Z������\�`�g.fD��5�Ƒh(T9�SexFo����.�rg�HU �%A�\,@iC�����G�?x�����wj���07T�v�����YM+9%9*��v�Rh�|A�S ۨ�}���	�n�����4v���Zل~�͋�';R���tR�t��Ӈ-0�����wB���ݍ��Ԣ�_���p=�~m�c���oT��X�
5�lT���xih�P����9AM�B�������<�\'����3���6V��3hlO@���S�QR�:{1�~���8�!��!�3w,�}�|M���s��Dµʅu
4�CCX��9�Y�A�ꆨ��D�^t�����گ����^S�6h�w�p�+�`L�ZAja����j�t��XZY�JT�4:@�J�R����XYhB�1���	�S.v�-Orӑ���I��r� AH�����y� �P/�'1ʈ�ߓ��h�u�O�y�����(>��")�kB�Xݿ��ޛ�X���rT��<	@7G�O���But�-`������`�:�ܨ����C%�ቂ�@��'ճd��\��%� ���U�����������S�6��[s�R�`K�C��>�����  �}�6�Ϩ�i�"�v��>H�mL�G�)(B1"�Xa�*v��9��.Q�{w���ŧ���45񅸨ژJ�$��_eFf2G;���wS-U�M�P��
�O����w9� �YqL2��[�N�$x\��}���('���-S��H�l�t��n+�TZ��v�ֲy�n6���ڠ�=�g�Pk�[$S�r�R��g�	��I&�<�nI��E��jC����	%s $��6n�<�H�]������3����_����;)3��=VCH���O����X6.[(ir<F 4N�L��Q�F��Шoa�`I7���Ҏj]CuM�U��䜽�������F�[���GTI*��=�.�����V	�=n������0��~k�n��t��c,8J�S��'z����mD��G��=dzm?<��]PV�kI�l��6̠��%�E/���O|+l?>�€�1�v�A�]�B� ���=ޟh��dH@UO��Cz>� V�`噡o�4̢�MO�JQ���Q|TH�
 ��N>��`d��贏�/��n�b� ��W�N��<�!ڦ5�"�JA�ŕ s�U��B#������V-�K����t���K��`\6�7*Io�ʞ釷�pM��Z��2�����>�o$�;^�%4Va�40��W�TPċ,X�U�(��x��@���}z��M"�938����G�E���u�U)�c`E��$>�v�� �LG�Y�lׄ�ho�2��Pu"�d�T�7ߎKB��3���y]��q����}Z$G�j�u��M[�-�X�'��>甎UZ�7��	(du Q���w�M����J|�i����G>��aš"�d
�CyH�l=��ņ�?@34�c1���/ۍ3؝�;D�S�tz�ˊ��U �9�,Տ���=.�A��`�i���mU�{t����/����f�9ʔ���w�d$B0�iC���S��̍�qBI�_���A��t+� 7�Ls��)��=��%:��Sh�4qyF�<i5�)�Y�X|�xg	F����U�&{|<a@y�w��.�VÅ�k[�J�>! �XwB�gP�F�g[�_#���o+���¸*�p�f�o/�j���uZ'��~��H��y��iƍ��|�G��|��j�;��?vU~9������5a�n[��F�(��zT�0�;c{�4����8^y����ϻ��ST�m��AH�C�n�3G�d���y�� ��q�B�A��e�
��%�������ީH�U��-����b#1�SE�Ҧ�B����[�sr�sPbW��c����H��2������*��>^��az`n�^<�X"]g/ō��)��������O�8&������Hb-6ɀ�a`�S�~N2cs��)[��EZ�O�u+��-p}ԇb�c\�̫0��a�Ǭ�}�~"����&����7�������wG�8��p�e���$����t-=VAZ�ĢUֺB��$� l��6�@R:���0�cH̢Mm�����wgW{O(�{T�sf�����#%c�-〤�{n�(���>�З�A��q�
^R�6��� Qa@���ݍ����WƑ��:DqsT��獚b{>�v���:Wa��_�\���HmHV��А����p�D���c���D��Ψ>(���L8�W���7��B��^���w�|�A�+6C�@��>�&���6�5ƙ��f7�PĖLO\'v/LsR �i���jd�H����í��)��_e�2E�
J�{���=����N����-�ɫ�
Ny��Փ�#�E�C' őF*K i}F��#F1�����hE��LUDv\w6S؄�4t�����R/�^xA��C�0U$�?�����J�t�����ѝT���$��`���`�r�P�T{m������������;�����ڊA�s9�E�/J<����X?*�(	aO(��X�o]�����J�B^,@�)��r{��±l�oA�R8�ް��̝7��3&��0�y��U�L5��m��>K;-�=M�Ιfd%Án�V2|H���J;����`������T�'�V�>�je��u	�"��|�c�kIO��иAw�����Md`3��u��K�ԒϘ���aY�k���%(6T �?L����G���n޾+��8'�ؚqK�����x�vJ�����c�]Ġ0y|�1q���S�&"���绨"i>�[H�َ��;3�^uq�R���A	�I�r�s��\�$߱/�O#�˔��]�KX�rNKE�.����w᧞G���W86ؐ��7��5XͿ�*�U��t�̙��i��o���Y��D���E6U�$J^���i�#�<- ֱW\��<f�A0M������Xz��!�m>d@����E,%�m���m�����:���g��=�4�z�R6�}�l;�|7���=ybM�)�<��*�gL`����']��,]�����\߳��3�XőG�-�G@��C��"ǳ�L��MI��w*>�����uXg:kk{�=��'� �jm��� j����C�u'�R���u�>��,���9����㡈a�~�����f��9؁n<��[˟p�[Ȁ|��L4΅rg���p�֏�`}*�(To`�'Z|8�\�J���Er1'9��Sn��������o;���:�x��E���×�P��e
ٟ����+p���]�^������@��:l���qвU*�?}QH������HƂ��E��Zl�&���̧]��k./L�_��rip׬d	u8���C"�I$��yPK+zn��_1\�**�+�1���M�c��ְ^�՟�7*���
6%׷��ƥK�V�"�����kE
]��^iN�}���Wc!J�e0}O�,�(�뻬%�h���3=OO�L����s��'_�T��2���3?q�P7ňUI�W��N˒�=}[+ͫ�� ����s�-��ۤ��R���ӯ��?�VqG5t��Fl�-���fL�o��������e֛c��E<A�(5gڗ|?�'9@����T��"���!��Q�v��x���~{
)���7={^ɯ�\ݓP��\_٫�[bd��h|�>��Y��ř�;�Uz�����A�}��@��;s�P/.i���\��W+8�S�^�dJ��f@��8���j*dc*���+���[�O��2�6'���t��h,b��W�p=� x\�m�8��,+u-�g��`�q$*1���hs�T�H.��w�������F�|�1���_H����ڮb�C�u.A*+#������? (�|<����b�z[,��nk�u�v7�L(ޜ�=JRŢH�UP#n�Y�ވ��"���v��sP6���*u"q*,O~��[�]tޜ}ʮ��p��s1�l-�}�/p��9Rv�0�y`��@�zq�_��:ɴ.�C�8(T��aW�of��`P��~��"ҿX�
NJ\��ŽB����Ŀ�X�k�R5�����l�Z�M��6,��P�K��TQ(���
��.�`�����[�q�$I�L�G:����5���	:8?��]��r��-_���mn"Ҏ�5���ǹ�a�p���X}2�	�� w�b|�E����fA�whqC�`ΖS�r]�~�g�l���6��킫��F�Ry�4��<��Rw!�+�F\��&yX�1r#:Y#"�i|��l3z�Y�h���{M%#�Y3�7��U�����T0�.���	u�Jʗ� ��S�ߨ�I1�y�NiC/E�����sݻ6.#�����_�E5S.�Z?�2����%	,{v0���D��BoiJ+��R�gઅj�	p��FD�����2<F�&X�����~�[�M����[�_��KKr��}_�?�r�߷b�F���:茄�@�3��1�&�*��Y���\v� �Y4����=����7�٬q�!�g!��?%�L۩aWa��HPz��H/3��d�c}n'E����ڥ��&��Rf�Iq>����	�!q��9(���TM���{���4 �T�é6�M+�NHŝ�K&Mᙛ�0��	�iw�2�K#ɺ�8�R���!�,\��:_��1���K�[�z������B6ʟNͯ�����.Y]�L�Q��cԎ@l���	�BRXb���;5C��g4eZ�����!KtE�ϑ���pW���h�;��������̹��O$�*���|�0+��(��\���!ӯ��X��҇�d;��3��i7�8l�[O���Dg@�!	�;\�{�)� >���.�ym�����*��s��K����~b�4(R���@1YX~�C�e��\)tY�8��g̈́�ʌ��m��U��1��/f%F���{R��a�r�C
)с��ZbKh�&Zr�}�t=�_S{j�/|=��T/�{{�����{K9�p�#ey�$\��d8��L�폚��9:u�?SɠZ�]N�s���dv��-2Yy��%a�6���>m:c����pT�Z�nA��1A�tQ��\���Wl��pAw/^3g�3n�,�,���dJ���W}?"Q�!.���߹K�|6Q�h�	@3h����Og9E5�h��$������昜�M�m~�<nr�������B�bԮ����]@�o͵�%I��*��b1Gi�(nO�Wf�����-�.,a���%������G
�3J!�d&ϯyb�K�W�3�N�=��K,�*�g�ղ�J .I�}���K�p������������twt�V��.�E���i��u�v^j���Q���2xcm�	�s��rFF��^;�C)�e^&����ޞU�Y�����q��εYnI"p�P��=Gхy����\�ͥ�Ij���4]`�Л����d����oP�o
�Mc�6ˬ,HhdEA#�.S�?8�M�0��gi9�j`9�֛��9��H��)��{��8�P<zD��8��V��0�Y���]����D��UbU٦ #� |e4GK/�b�=PCSߪH�;����=��*~S:#��dzŊ$��B,��]����^���DX�.'|SYFK��Aʌ�l�As)��[V��D�x�D
��=}49�Oj�Z��4�G��K!��x6��c��Z$�ߴ�&6g'#h���9�׬�Jn�Җ �Za˿�v���A�ƃއ��)����K~���;�Tq��FAk�b:�Z�x�@/� ijga�L���r��s��eL|�јB�v&������FN��k�~��p��hr�1����ƄWr��/:2�K���q�Qfۢ�f�(3��yi�f/-X��G��9�h	3�N�6�;�-M5q����k��`��)hՁ��?����R�h�G�\�����m�N�R�ZY��hl�R�s��OC�ԟ��p�ڠ�Zq�=����3�!����� ֭�z�5����"8�`�f�
X���C iW��;�@4�e$�-\k�O;�.�!�u�?صp��G�o��yx��� /c>m�l��w��-국�l��gϋb���-r!�V���@Ф���y��� �ʄ\��ҋ��`�h8.����wو�VYXK=N�E;Y
�`����zS��3�yd��U~7K�DI���d�C벉�+҅�QT�)�I�al�QT��):ma��lAo@-w�e��95����Z,7��߿��'8���B��}Rޘ���a����	��w���R�H�%�����������Q�W����4�Nw(-Kk��Wk�l�Y��I�m�=O��������H�)86�ͮ=����OC�zA�{��	�(�V�iZ�h#-��}�\�U��p�̑G�HkK���#����pȑ4S�ht7N�;|�N��E�J�����q�ѾA��x�����Mr�u_8kН7�}�>���M���>��X(2�r�
��G2�cc��d�Bֿ�E�����G�5C��n�$�1�Hb�B�a+Q����*��y��)�~�6@3�+�BϠl��UZ{X�rT�⸘H�H<ǁ�k�-wl�w�A�yz��`�}#�|vi��oJ�N����|k�?�O�C���ȸ��7�$�7.�=�6���$�Q�l���%�I� "hG]"��U{���gY�Б2�1U�����ۊ�Ո�A������B���\X��W9?|k�/�	�� V}x�`�e�f�,��T���@<������l���/�� �$�~�K����LG��_�>#h�.������|:v�❥�z�]*A�H��O6_�Kj5��i�l������s�ш�1Ï���6�f~�sjF$�Vzi�|�p?�/�7���o�)��S`Y�׳�&�T]�C����j��Y���e ��fwL#b������=�_���P�LAFkP!��	�@�a�[������&<
��[���l��~od�cbY#��7��IX�6�~\���(&V�L��vo�i�=n& h�2%:�%��o��=����J��fK�Y���B�`����y~�b�2�jЫAH�]�7�^��i��jkHL[tE�n)y�E�9Ҫ,/�����>�"��S��s�xd9�*R;1���\jHr��S������,�O���C�b�V��nz��1d|z��ĳ����ǆ�@�C�����V'�V�"�{�+i6���O���ٕs�`o˅�@XT�%�3p[���`m/��o]�4��^��o�Ud��C���u�JD4�+�/�X�
�"M-���x����}te����]��G~�ԁ.*�W�5�Ī���o���^���!u'��X�6COX#�-i���V��&��@>�j���}��rSt?/��&ha �X/&�]u���3�bZ�m;�����xǮsO���?r����\���k���B�L���o��sM�i-RC���>դǬS��:�'&� 0�؜�u	�^��0��~o�8*��`w���)����tÎA�ˋ/��M7������=^����%}��_=�Sx�U(�v�)���w� ���ขxR��
tX�lHK�D�k��^x���!��@����=��|�l]]{���Wb�c����h�i�7\��fWqj0�,/M�e�:� 9�	�Q��$>�a���:�u���2u}�ڳ.P�� �"��#���F���Y�*�9�NO���Qs�d��n0�?�P�EV�W��C�x�v�^��\���6Υң�x'B"O
%5��
�'��e��o]�1��.Kq].!����k��zݱ����ɺRcZtܻ�r�v�<v���up��FԒ\{߃`������)g��Ξ��YJEwd��:d��Oh��q�h��i>a4�t��HD	xC㠟N�D1�}.���Pj�Й%��Xe����t��� �UK������_ؤ%L�ǀ��l�8���NF�n����,����<�bpf�6
O8�p� �)�ځ]{E�z�l	��[��R@)���ƛ��S��f��R�rZӋ�'J�8�Ob�wW н� HG�m�H|\@�!ںJ��Ob�w���zoܳ�dY���ߋ�z\v�d�-Y�_:�*�caV�dk}n�SP�R< ���7��5K�̛��7Ƣ,��jRa/�O�'���&�J8�p��x�_�dw[�I�6�����[k)/v�.�3W��-�^�������X�xh��,_B�^�v�W�t��풲f����̃�Ҙy��F!����Fp�Ok[����2xR�v�>��B�LiOzN��kN�=1���\6�XپT �-�>����7>`��Bq�+Tj.��������?��7 ?r�g|�>�$�C߭����3�7��G��t��!��L]X�>�2�*A�����@���N�;������߳�w���Q7��^WV�Q髋g�������AX��u�1��۞�=��|"C@J�K�@1�fl ��ڡ~E4|�ĺו�>��E�d0}D��`_���i��q	_V�hEY�B	߸���:ǂ۞K����e���WwUU�>�rz��C�����l���2W��H ��꿹97sXo´�,ș�JFb�j�]��g��$Z�$3�����PD?�M�פ�1�Re��L��]��>�6�q7n������Òd�u���ߧ�n�p��U���x��/�#%���)��~B�7�H�)q��ۥ�d�%'2OE��I��-H���aQAћc?����d�H8� ��~b�?k�mÄ��Y�Y����0z�"���;�'+�T�"z.m�/�����o���ǚ.�P�4��i�B�i�����Y
��ן{$G��:�`��Eڻ�jg6H��4#E��ǃ�t����$n"��,��������˩���c�i���,��f��S�����%����|�m���l�Z����L`�isyP�t
�)⟑�C�%�"����3���o��C�|jl��̓�o���j�ߋ��1c��g��,Y�èڗ;�em�+y�w�X?�3�I߳�p����dT������Z˽����?�ONK��n��G��mgq� Ibz�>�ZĚ�ʘ��CaZ�; ����ߺx�j���� � �2nF��H�n\R�4��k��gV��M�"�[5Y}P��9�V�ي��I�aS0�W��E��}V�0�~�
��[p	[�I�d�4��2˒Fۺ�£�şz�����u�W�~f�5��,�P�io$<k�W�V���uɥ�����%I8��撋��_����}	r��;��l� �[J�]䶟���ץ8X�l��<R�r|g	`F��v��������u�h@6�"�e���7�A��v�ó��RN��;��m1RM�����įw�
I�a:Q�G�e�T_(4��8)ߋTʭ;!u��Xw�p�[-(Ew��W$?,4V�'���>q<��p���G�,�B7<�"�A��#l_Ɣܲ�Mgr��QS��5s�{��,U
X1���ws��5r\ ��:B���
�^"`�7ŭ�l4l�ϳ�F�|�)�Rʡ��A�-�zPJ3�l�u��H���#;����yF�jNX�v��[���É�ZF8Bu_�����G�����U�_a9~G��{�c����EL��0?�ΎğĤP��%�O�<U��(����ɘaR)T�3�6ړ��MϺ�����uhe��>�In�f*A{Mϕ���-���>�S�>�7���Cpc|G����H�#|#3x� D\X/K1���bUy��"����2�P�IQ��%���<��V|�$����w�-�h���8mtש�E�����	t֩$4�9& O��+�9����r)�c}o�Ҡ,�i7wRs���*A3��k5����c��7�஘��$#�벌��3h[ʬ�~Fe������.��S��B6ꄎ7��ƹ2�rEgH��=��������7�Gc�*��&킼F����C�+���0җ�ƻ���ي��ýa��-#?�H@Q�(44B}+����0/}��\ٕ�L;ΆK�F:�r�Cc��Խ_�U�ë,T��6|S�]�
�w2�#{K�'H��T����h�dXt+�)�1�`��_�DR5��k >�7�=3�D�<Vp'�`Q���-9VA� i@����⬘`)�G�.8���&eS�Yg��h�2�Y>"o����G3"���,JPP�Х���@;�X1��.' $���ꀯe��#�I^9I��AEk�<��C�R*�LU��f̳8�fu{�(��vl�g^�CQwC�!itً��̿���[aܗ%)���&�"��P�AHe�i&��X�����}�꒲$U�������A��!8]�a!J�;R��y,����1ˇ͡Z��ֲ���{�E��(��JܑUz�@j\_Wps���0,��N3Y:%O�,�Z�q���[���jd��G����_	�K���������������G�7�i�50Wˠ�Q4�~X#��%���NŲ
����o�Cb=r}`�9�� [{*�7�Q�<�8]��@�UO,��j�f��P/�?����bO�����$l�g��� �tQH�`�V�MR�į��0H�*�n2C*��F���_���ڲ�� �N)�ԥ�(ٙ�2��(T^prK�VU�V@��o�3���%L���CO��L���t7�CqW��K ˶4��������+�g~׷q�'��[�b�ʍ.��'��l�r��F�4,
�=[���G��z�J]�'���@;,l/��arN0T�y�>�<�/���b�߈~�#�e�Vu�losݶ&2&��pZ7�"5��I=�Tߜ��ܟJ&M�ff��"ܝs��sc�l�
V��}�/�T{$B����Эl���n72~�&�d�����F�t��F��쉗��3O�۝�����v��^B�0�sZˬTz�'@��&�qƲ=�.uMe��M�	F�4����m��?w�Mt���s���mx* �pwKo?)'Ε���~�T7���㬯��gAE�4��Q$?�_���, �E�v�7C?�ݙZsk����`v���~�7uŷCG�IAM<!��{��I;�+��ȑ
�������i�,��&V*��� 82����Q�����*:�������2ᐓP�f��0_���\��K�w�nb��$���d�Pk:�G=�l�f���:�~�ƃ�vqu�]E���ܷ��q[#�j�WgPѨ�����f@ ׄ�*��v�Õ*��+�:h�o��D�N�|�����U�}n�LΙ~��t�!��q���t����"������PW�$=<��VI(jV�"�|c\��7���ⰴ�5^�q�`}J��$z��4��HTo�)2�> �Į#n����L�KA��`}�C��?o�lͻ��d>�h��D&��t�@�2��	��ͅQ��F�o����]2-���(���ҁu���9�D���$�lS�	%�J�@#)�O�wQ��bX�� ����;EW�Nxp����5�ަ�̹	*!�iW�î��#?�i�0$ ���,̂��׋�A��q��|��ju�a�숯��D�D�Oڼ�[�f�C�MlvgjQJ��m�T�Ru�q<�|�Ё���ǾEuix�D{�En��'��o/��T�1͔�l��`C�=�F"y0b!�"<�m+�5H�x7��n����E��4O��+9�<f�u~y˧�����~�V��Z����,5r��z�Ь�����(����� �>yb�����{x/\�(�1�D����E��3#H�2M�;H�7; 5d�n���w�n�!�&%>�pҐ������	Yә�yC��뱹ڷ)?U�S$���3*�zl��xO���a�d �>uR�*
ͨ�=��k \�vA��ۢ�2UB;��ء�[��j �JW_��{#Ձ�=��m&��n�n�aк<�~�����.at�ɚE�oU�-zs�E4V���p'..L	�[�����]ɮm�8B*����j�i�;;;�-�`۹��6#hם�:*Od��2��p���FTS>X�h�X��Ѱ�|�y05���ń�m��Tl�y4D�H��&n����aBb�A	%P`�։�
�ւ^p7o������L�0b��23��5��WZe,3�e�@D���&5����v�(��B���β3���x���6)H��[�����x��� �'b#ݛ���(��%�Jh����,�:'`�]�Tf������s���3�q�6!;Sj����P&�,_���L�"��g����<��u��_���#b��0'����$1�4�9C���=���NIS5����p��K�\rϖ��^aJ<#f�L�=P�8b:�6�7�k��*�$�-uTx�Z��ͽ���Ɛ@��@�Z� ��E-n�@�|k�]e0��|�Xޝ3e�����sf��:���Y��n�̰���žG�ya��Qo�z]�U���m"�_�!+�,ɧ ��VV�>����K]�姞r���%���F9{��P�%I�U����W�i^c5[K��O�>z��B�&��^j����;���?-��:/�Ib��}Z��]>^�ofi ��$�4<�Y=`MV2�\ݫ�	�g˫�I��D��gU�(ő��u������̯i�]��m�Q�G-�P)��P�_-������,VO?O�_,�'�W�1�W�����Z��h�0#T�9�ru�� Wى�q{[{����� ���%���l��rǠ/��ȾI�ì�$��7�`���x��?ԝt��5��0���&�!�&4�PI�3=3��%�o��	%|�����oܬ�9W}��Rʬt�f ���Z����v� P�y�S�^�r�d;�P/����]�.�C/l������`��W�彦�a�NwR�D��A��5�TC�K��J [v g=W��:�˺W����]L%.2� ϋ^*�6��띺v��\2�X�?^�����Lڽ<�����_�&ˁ`�mo��?��M�>1`�).�6����\Dnkꄓ����
8��]�u�����#�ɩC.�g�B�i�Px����;�Cu�cǃ.<!�͠�7��7^�W�_ <~���%�����d������y/�=(���&j.��Y��<V�8���}ˢ���mF���b��q�&~w�0*���bM]@�ػBS�h#w9�<��%!�w�*Y�h*�ƅ�.���h�7}a	�g;���eѷ�Pj��['�7�|�\n76|����#�\�Ar�T�;�!����~F�s����_�}��W�rVh��+��kjܴA'���|�kעF
�9�;�QZX����qL�� 'S���\t�K�l� ��})���2��<�Sg>���Gd�g�iڰ}4�eO�T�iIY�\W7�eV:��������W�S��L�����?���#�����"�fdc��>Y�����p�Rjq�|M�m�7�����zI=0�	�."�2q
���\���&r�5Q�J�K��T���
d�g��!9Ę��R)�\d��h�\�U�=[u� �&�I��`a��[�zf\}�d�ǅ�b�Rz��So�Qq;O1�Fn"��H�5@D�6�(V��<AE�ls������8{��*�Y�0�.n��;zd�H�Ɏd��ލ�*$6�������F�,����7�?����#��Fy><7B1ƯӶ�Bk��}�=Y���HMg`tf\��3V��nh,�I � ���\�(��O#��L�3<���,N=Y��l��v6���?�-�<�;56		T�Z��3��x�W�˅ph4e�aY�}g�毆+���Z��C���P�hz��@}H���?�5=��@��*6�fs�g��2����t�g!��7�G�^�M᧱��b����a`�ʱ�B��6���6SХ4V�P&	0��QV���d��ᄓ�=\��"�E(>~y����W�t��nƭ<�*i��Ƚ�0`g*�&\7#��j�7���������t�&�QJ��]���_�YO�F��9~�\���L#a�G�)ㅪ���V{�d4p�t������l�x{� 9��^�3u%_y�߹W�5Y�N�\C��6"�
��&�╂BJ��M��2@�9��Z|�+���E̓���1��!��6�~�c�>���s��l�Lū��IE&�}�|�_G3P�/�y����K�iވe�U ��{��%cgf��Q��	�%�� [V^<����2�8E��|$���p���v`:ږ�ٗ��Ш��}V�ڪ�e��� ��Se���{��8~&!�Qr�� "2H�uЁd���>k�+13�q�U�'�a��%m�w#q{r20��;G�g#���\O��yB��Y�P����}(���X �v8�\�$a{�.������#6)H^V�k%ٙ�)nR�|5L���Q_�?���qL����ŀ�d�K��&G]Ѥ(QL�f��S���6>`�E�x@���;�3�;@�2M8����3�L��`�{���7 U7���)� �~r]}���$}�"�����!
�q���=eӼQ֐���j^�*d���\r芧���"|���4#]��F��kXΌ-��G��C.t�G��V��wϐg*��E����j��n�]  WL�~p�&e+w��4&��X�
>��}P�h�d�8Z�0��&���~'o����� ����RlDt:��f�O�@��K��N楇���B02{��8�B��f��8 �[0D�[%�I��2�Zoy��!�}m	0m��$�Ne���cf6�ZBQ3���"�	�<r����4��U��v�$)π�)m2��zlQM7QkF�0��V��W�ew��d;�̃+�ҏ���Ѿ֔n�j '�}�^���)Nm�M�I�9����*������'�y���c[���L���nވh�:ˢ�?�:�?�3�$���� �\��N��d@a+�����XNW���Y�Q�[Ψ��{�^��Ի|��ᣃ��q����sJ'����@�k��3�����.$?�0nu���[�e9��U�f����-V�h��B.����5wٺ��  �kL>Q�9�Y�Q>�˥�sJ�O�L8�V�E�b����akch2��H8�7N9}CNQ@M�%J�S5�����]�]�� <�:��<�S�s���I�"�BZY�q|���]b��.|3�pl=������^���%�1$��jYh�'�|��ʯ��Z#�����#{�֥�.)y1զ`����[�z���֘c`������5��> �RV��Pݞ�⽖1���u���+3�^�����,q�(�V���>���RC�[E��|����<.�[O΋~�u^X[�o�Hn���jX�C]��w������n�߭mo��$�Q��D�<wD&\��n��j�de��ѣ���b	�"L���E��c��^|�O[y��g�۪�z��D>�Ruϟ��<��G�	hST�˻Q
�|���:1h���ک�׿���1�����%�k����1�{�A`Q�����^g��˱�+\B���fhs�4o$�0K74i�
^�N0'��xշh/����I�6Ji�dBd��bz(k~�lɫ��m��iF��=x�\�c�b~�'��/��Bk�4��m(d�f�l�P���.8�c���n�RQ�촶� Wb�T�w�(���0k"zi�cs!ͯj3!���U�M~2�?��_0R��ހ�{�*`zBQ$J�)�Q.�:�I�Z~�}R��q���4ڿ����t�H�6�&��&�9V5��C�Q	 <|Ԩ_T�w�&��p_f7C�����k ��?>���#}�$���o��}@/�KJ�o1���H��|=Ƿ���	KY�ÿ�}%.(����Q���ɶ-�A0Ê���eqm�H?�H�7�D�/+�:�ҍ$e�4�mQ��y@c�~|R�D�7} ����{R 7?�g��_{��v8���|x<_���	��t�,5�q9��C��y8�Q�%R<��u���&��+.7�nO��me�1 B���i8t`�����8�����&_�ɦ�$$	�><f���"�r��^��׈��:zr����I�q�੸���<|o��A{�e`��n"V�뼷�i�4j�k���y���R�W���A�ӀiEn�ω2�Љ����ji�]�4B�4?�$L�����1�͖9���|SNT���qț�;N��_�O�G�#��e��d��h
��sH�\%��
:��X�?͂�'A�>K�^�q	�m�����.Mk��r*Q���'Ϙ��&�8��K�%���f)�_7_K!&Z��'곳i�jj�|۵�Y8�ĄǶ��na���=��J�����@���`���<UQ��謽y��p�+�G���6f��"�f��d
 a���zj^۳�Mb+b:�(�k��S����%���$;q�Zs���2�m�ێǚ�x\��,C8�#yb��{�I<�=��aA��{�\ +2NAkq�<bZ�_Q������ݓ���*)���f�F�Vq�ݚp�G-�ҽ'tҎ�M%�����I�h٦\�ÒX`GS�L&|�i٧��a㎂�c�������:�}���pϘi6�D���^?�	񳣶d1"��L�ډ��˰b.�U�rϣ�|;_��L��*ҿ�Sx�i6�i�~����F�Lu7���R؁��W$��oܷ8H�Cm�V$4�Pof���p��{@H3#�ο���Z�Tk�H�}�����}��L��:����3!�
Ös��R^��	ˀ�����t�H���� ��)��(gy��y:�â.��s�n�����4!&��ǤU:��[d=�`�ZRc��FRx.a.J�m7 B���b�.���-��4E���2�{���p��2��M���}+��[��¤�	}7O�!��$>
�fg*vE�Җ��Ƹ�VQ�G�>i�M����74��	)��&;�F|�ﮣ쐟��ߜi�L!��ٍ���mD*�(�7����e��`��ą�;�(PU\��Z��fIԔ�x��,��l���茢��������_�S/�}�u��hd����iksd��fwՓ��ָ�o��ԙ�EM�b�'0|��us�o0[���CD�}s�>���y�ZN�{kXzghՒ��kEҳ��7ĵ���ĭ�������J�u3Ӊ�I�.�cs��(�M��<�x1fW�x��4�(�H��Y�p'g�y�����~\ �v��Z���d�m���:`�J]��Qs��������Ad��o�{���/x@f)���K�4V��!�����1�/\�m2��-k��mԵ+��-?}��7�)M9A/u;�s�L_OCT�^��@�s{C_kܒt��o�)�k?O�M^����M炘	�P���j�K��Mo<H�u�oi��C�w$v ڄd��I7D&0��n*Ɔ��!G{�62�P�dm�̺�U�#'o�}z�;���:�'��Bg�oe�*�A�(�|T�/1M�P~��M�5���@�f���Pt��8D-a�M8�I8���R�M����� ��^�g?�����2uA΍n�`Fi|����.e��6�g�(F�\u���O.�C�ȵ]�����tL���E+|�Ԁ�}Բ5�^)����td՟.�/ tw��/b3	�&�`��2�Ӂ���䥞�x8|����
|o��'���]�Rh�k2!{��U2�>!(�06&�`��T�7��<�_�@���Զp2�+���k���}�Ə+����9TkW���G�Ohy܆K�
G-x����U�A����){bR�Q�4�k=�׫9�5�׭/b��R��k��M,����-�"T��O���*y�]�.ٓ_3�C+Q��Ǐu��zT�̺?���@[}���ѧx��	�u�9��o"EN݀�	AV�W��$��08���0���@��Ķ`.������'Z� �zUhkh��8���@��uX����mU�8*��Oi7�9���?_?��e�x�y�G��vH��=�q�\���l�a��3 �4~�]Z�k�.��)�����n	��m�(��ݕx:��bME�}����h��A2x�����tғ[Ӽ�D�< �О����{W�PC�u/��s<��>"�{��H������]�#�'����\{ԯb"�ē8��=���.�L&!���SE�KZ��-��+Ϻ�Y�9TՄ�²ߚ]���z��H:�
NJy�*\�,�${��ư���� 1�#�p+����N�y=BIF�j�2�e��C���Gפ;=��M�'ڭ���T"����dn@�!9͠Cg �}��Ds��Ս�;��w���G���v^���ge����l��ZQ�>�?�P!'\��x�hr.`�|��Y��u�n��y(���������j�_6�u�v�pEp.4�p0�ӕ=Ni(�CE���/B��?̖���g��+�qfW���B��.�\�5U���ܣ[���r6�;>ų��!?�S�F�#�=A[�j��egN-M��1qǨ�����H>,��.e�9h��V�� ����FG�lC�ʇ�8�r��4�v&ϼD���S�C�/d�ތr%��a��C	��[R���c©�M���pk���"}c�z�\�� �)�o����O��)������K�"��b~��"B��t:���v��K{;|0�+��A s�L�M��7����c�Cq�J�.�Φ��6}x�[�0v�`:Ef�L4g�q�� Q���EMN*���^����d%�@������C��!��T]ۣ�i���ٞ�Bԙi�eZ��N2��(�9�X���I�^3��P�\�j���NAk�'���B�QZ��-���5>v�.����C�_.�S��������ӌ�|q{�k"�j�L�9��J�8:;��Ų̏�]��{�'��a����CA���ҍn�L��Mȡ�x�b���v������Lǝ�Ƙ�gPKvsj�*���\�REy<�\Z�0ΤT����`����b�m�*v��0�eBM��o��c�߫�G��?�%��-��+=�����/e���m�Q�?��h�1�� ,�נ��H|FX��A�������A�㙗+ŀ
�b���e=%���[k9DIF��r���w���~{���֩P9J/|�pt��X�RW�r�/��F�����K"]�hb��v;��IL��$10�����@ZGYʙb�Gp�L������g9�CI�r1�U���V&����an�Yq0-e����݈'��W(�|��#�oMIo��UeX-k��Mr骸��������=�Y�P/U�(��#b},C0�3�D��j��-r���Ҝ��iL%��v�l�	�Gk�#U
����*9{>�9r�L�S��s0�h'����h�8v��Ź�X������A8��|�Ã٦P�@���DO����y��t�d8�vK��N�����X���s羹l_��;z��cӴ��,�9�cnH��(8�IǛ��@IQ���,:�Kl�d��4��{w���QR��!����F6|w��s�q8��k�	��P�? �1�B�����|P��b�,ܔ�D̸'�� YF	"	}u�nj�>8��ko8���S$Ì���*TF�C�>�D��rQ4���Lic.����㚖~Dǅt"���0Q4�i�h2X�{� jw���ᬊJb�><,�B�mTZU�'�a��/����Aw�j���{�~���K3�c��e�A�����:|[|�'8]���񤈽@[3����e(��l��F�u� �OC�C�d~lv�!QTl��X�I׽ׂ��dL��U2e_�Zu[qmA�?�V�\���I�����n�<���U �?��ɖ�垩b�&x��W<��AFȈ�?ǔS���%t
�Rb�a��Ro'	�t^J��d(�%3��vn�}��1��UoΈ��_�V�Q9	Lwzk x9�;�7�;���k>E5�*v�� �j|و�}:�D\�:F-��l�*���j�|6@��퓧]��>9�|`�<�$�>]�Tv�Q�##�Z���P�}��-5^[J�3+�Ӫ����li���Ľ�q&�����	i��GV���C��u�h�b k7j���F����ɋ���y�>���I�ޝ����y��sCKD���y?I}354�]J�h���䯣b�O
��T��i~g7k8��$%��?��(���4y��a���5�/��A(�NZ���=��h��c0��۬\��k!�ί�k��k����)ھX w�ou�����}k��Z��m^�R5/��2&z��^OhZrm_e$J���d	�*�����ݾ+�K�n��k����3�{�*�S����ـF<M@D|S<k�B����LZt+VΆxxE������Ӵ튛m�N����(����T�Y��b"�#�o>m�ϪI9����3�yo��SgF���V��8��Q�9���~$���Q�+� !g�����{�X��/��V�΄P�@�Uj�xn=�,�����t&퀱�pK�3�9�[�_�����Is�,;��F��0=�7�Tr�[����0��9����rN��yE|����d���M��S��V�O�j��.���;X�I>�	�P�끱��ZH�*��R�DW��T��T��O�s0�n|Y�9<;�����"����]H��i��dն�E��(�e9�[� �N@�K���i����Ty?Al�YF�2�p���wY��L7�6P�[�)K�1Ә��M�{b���w�Nl�T�[B_�-[��rP�%��䂢��l�t��or�O�3�+FG(��4��J�k,E����QR�Z��V��t��6E�B���R�
���s!C�"�0*����kTz����.�#K��.�2q�������������_mB��/.�_�X�L��<�Y���a�b����@ߟOM�ԩ{� ��Jt�	>�[�}������}�9Q��/�����Nꆈ�l'go��2@WK�dɹ�rT�g;��z2��	=�Twq	�en�\�|�jV�u� �z{���<^<̡��z��5����]E��L`w��2�
���̠׸RL���Hc��=7�~���ƓD}�o봚A���1޵)��p�A���Y�.���Va�F�q��8ئ�ے-RHJ,$5T�.���
<�c�}�	��j��H�c�&��|�;�[~�]���r�6���	q"��9�0��o�h~�+ۍ�\"O�k�c�ݙu�:{�mPjH��n�& �Rvp;hש���Q1T�������x=��zG�y<����B��e3bh��:���Y���)pc`����\D6}�Λ*���4�_�u�d� 5;�j�w�~i8EME�zӌ�������j��c�#�p�K��,��XL�æ�i<x(���@� ����l��*/����F�Dy�=�ڿ.@��*�`?�i�ŭ���~�}�W�a����!�Uⵓڴ�_��y^XN�[%؝\kI_��+GN��m���������៝��0r]@GgJ˙��ъ���t��r��*ǙB?'7"7����!�	��y��5�\,�c`��gBo��fl�����P`t������U�J���F��V�˻�0��}.��\�����tpTL���|�k�����5���:�on����ZVR��d=)	Ú�kmA�ŨJ4��S۫8�v��%�ՠ��"�|���9y'`7��#ep�S߯�����r_���L!(�rp/ڡ�6�u)
��r�m[�#�Z�����]��/f�P���{�Ob.��J��3Qjr>|�H�WF
{�|v��ǟ<��~*�G�\�a�ş�.�&^'~���q���܋��G�q6��5�Ŕc���e�*$�g��HR�)���;2�1*�x)��O{��ݒ"�tq},��V�N��d�3�tJ>b(�a�8|� �9�}��=�W~%�񜅤%��٥��gUT�V��`�����c.'FXv���SWzLX;A�ͻ�<��-���g�6^W~m�B�x(m�"f�w���H���T1I�'��&��Bn1���sud��RY��ߺ��&U2��
ځ�AӀ��[� ����Kx�8�O��!��+�G�bf�>��r�)�O ��d@�oYg���	�׊7��ֆ��;�r��D�3�-�B�]6+�X���e
�t�>MW+�yUh�ڌe������g����C@�~͏[,�9�D&�ֺ�y�2ʫ�wwD��z�'L��S��%�p�J��B�5C��I0���K�V�)P2��<}�Z/��I�B�Q�2E-��v�2�luG|+Л	V�Os+q��$�j.�yj��桚U�\ȩ5����rt1q��t��Ҝ� ���@��s�&�,�ێ�h+�1���ƅ&��R? a�&K
d�
�pI��?�H�����
���/�v��*�GQ����=����G�u�������lr��V�̥�ҝEJO;$�b���e�y��Y��],�[��H����.�}��9&+i�{h1�i�c)ne�]���L���w#��q�pMT�/1�x��|vV�o �CE,�x�>7���k&W��U�A^�~o�;ơ��t�\K���re�7��3��xt��L8�a�/�rԲu������{�}h䯶�ˮ��R���k"���[�JpS��8�����`(�+mcгY�y)�|Z���
����Q��r���y�F�+?ͅ?'��0Л��y���W�!)"0����U4��ʞ�:ҙ�\@��
x���$P����J�>NĞ�I��T�G��\V���Mw��)_E� �@⽞hn��C����
8'� ���`N�)�<'�	�����c���$�h�:�4~a��%�!CXa��Jgv{O<?t+��B̆M$3��%�.��#_B:� �>xM�i`�!yK���;�&�!�D�ݱ�Oxa��X^@V�Qtn�����R<���,7{�Z�nִ�`yMo�Q4X�ʃw�.��HՋ�IQ��k�B/���G������J2JϵWT3��q�Sg�}�X�Kբ���c@T�a�ԣ�p�A���ԴB�Wb���ё��a���We]��~¨����K��g�~�����Y�<�f�/f�S���v[+�=���;M�N��إο]��T�(w�$�((�;���z�7ke��l����
�U�jYx�2fC��j�z�|�Jm3��d�F5������ǭg5�1�T��0Q�D�H�{���c�����6h�3ϖ|�$;:09�<��/�H�����M���	���a�ksG�@�u*z���
C�ɡ���7��\K�ҘsiP��Mr׎�\�E�$u� yȱԩ�ax��	6,�H�7�X֕s��k���(������C����E�5��ܜ&=N{,����ݿt㡓�p7[����.i�p��yv)[�g�{$AU�'	������b��{;�ޡvN�Qzҏ�;J�U��g�U|U���S��� �k�Zv��lo�0��a�k,�����T;K��$N�m���6��f�.�.l�rJV�i�f��o�ylX��h�%&$��B��Y�=9�6��E܋g_��.��oVϣ70T���olL��j���Bag�쯊�?2��xK#������)h(l"��Mؔ�Q�� �U�d1����軁Є���u.���h&1���-D�޷��ě�1_M\8�\ISV�I�ޭ E�Yp��F.����A��[ۥ�����ٽ�2���&��*J�Ą$x|�cj�D 	�4�P@�S �w��H�Č�~@)�b��5gM7w��&�~ţ˃?�Db<��D>�1+fڶJ2>ѳ��ef A��L}�y�J,eS�}<��ܞ�_6�T�����D�;�\�(6��_����i��Įf���N!nhx�ʪ�ԡPrx��*	hMvg�%o�i���:w���j�����O�Y�o'+?4L��m�~�'����yo[�G_��a�%g�	1:h�s��څ�6���a����������&�Th�}�dG�6:��0q\X��M�G��me8�m��K�nj4\�C�c16������Q���(e�-���pF�x��Cz�"�/��@�idekZ��������M�KZ~b|�{:��a�#�!�����o��- �;ެ	�=NKX��4I�����'�+�c\'=��Sw^ V���B���3j��P"e�8���ҙ��"��e��^��]�i0�N�P���( �\���/���Vx��8�'xOc'	��Y�PT�
8�,�w�cU7��Zw��z�N���8s�V���,E!�� �W}���}PH���T�_�x5�˯^@'�vۧ�T�S�����Fw�h�f�쫀�F������n;>V��5.��3���
%�`H���+	�m�f[Å�9�oZ	�/�V0�O�3��W��2������5v2>zV>|��*�	�u;�*2�I`|޳LC�O�`z��9L�B�f�����lTLD�O��)��Q�14���8:$��6j� ��Y���;#HH����X�8 ct�����Q�ȎQZ<��C�{�6��L~�� ���e�]��aC>b�������8�rlT��s�CmVL��WA��2�xIG��y�G��鴊�M�[}�-�`���o) ^��&���.�ޤ����Q�.
v�,�,��^��$8�]�P�A?Y�V�!T������;��ڧ�p���e��9QGc-Ԋ���o<�L_Eן�FTET�u��M���#R�y�=�d����ƚ���y���@�}��'�a����b$ q��b�"_y�1�����|��_�MD������Db%�O�e�2t����}=y��g�W^��5EѲڬ,�_8�Z19)��p�~�F�����X�,#�Ȣ�U�[�58�#b��H%v`���8{��^ �n@�6
�́��r*1A�D�Z1 ����n�\�q
� 9�zKy�R�Q��:'Y��#6W@�Nb�������@�ė�����Ո�����n�*�L��j��s/�cE�$�1�|��OT7`��nV�R��>g��J�U�����_��_�ՁF��W��Ѕ����X��)��י�{^� �8�}��-1����%����q���.���Z��%~ �rA"��FsD�:�������$[��pA����"lU�ֻS7�,VY^\��Ț��(BT<�[1�H���X�E����=���z��.��������TB	cP����/�G(?l�� a~F&{[f ���a�RD�F���6i0��\��=���6�N-n�傄��8^G฿_-�Uû�O��5������ ?y�T�����7=΄�Þ/�kw�e}�e�RSD1k��S�����0*91&
;���=iήT���Vz��?��~�Lw�X�v�7N�]����DK�U���~��� ��o��dVdm��O����[�J�!��om�GۭKA��{�[��P�:��*�Mh%+y������o�h���-҈D@?w�V3�Wi�Sl�\�A�Uh�[}��ӡF�� ���{gJ���v<D����
�"}�_z\c�� �P�1S�����8�ԯ��0����|ApK���jq���X�XFSP���>����3p\�l�J_	���-S7���I�H�W�mv<H���?q��OςO>������$�ү(���{C��M� "�ؤ$�ӌf�-Z.�V5������G����� Ð0��hF,Af<�9b�(`�>#�v�0�v��	�@�����cԟ*��g1����M<9��2��P,}�+8�r�֟#pI����\�XT���5�W�'ޙ��8C��m�-�.�a�@Q��JR_��+�\o5�9���5�B}_�Dߠ�G�DH�ǇVȚ��6�(R���%a��5�cw��0I*q�n�Q0�ǫ���pK�N�Z�V�	wTgo��b�o�h�y�g�ԓH$����>�����%��@�-��L3�Kx@��/��� ӌ�r++��f�
��:��f+���ge�ڳ�A�V�1���ܔ&��46w�pQ�<$7��Х�>��?$�_'�;��
`�n}��Ȉ�voh��<(jZü{V`��~iN�>s���yZ|{��{���?���/B�* �ZI+ķ/���Ǆ3�p���� ���K֤"�u_ɈM��ޠ��d��LExj��t���d_�Jm;r�z�r�)��=T�)��[d~�J����);����?�dm\��iIw��=4�[�:�CN�o�-�
S4��=�����`��ҭь�8�,
��e������[�!�3�k�A�z��#�V� �[(��kxF�m�3cOe�[��f��UYzE;v���w������k%-�SR�3=A�Cb�sq>`=If4����+��i7���G;�������S��9�b҅�!��oc팀wU��'*`��o��>b�PU��i)4*)r����F[�Ɓ����0^���5��
c�ġU$J�&P�&��#2f�V�[��V��kĖ��������XӼ�6��t��!����,�.�{R���D��L�5���u�N�r�	kN��w��v�y�&t �����0s�0p�%}��G(��L� O:/��Sl��"��1��1�j�^Bӆ`�%�a$�.�<rO�ՠ���53��N��n���79�\`ԣa�jfL�v@\�U\�K���S3�����?�Y� �|v�L���tQ���Nh�)��!f++�V��(�6�����SO�k�T�P��Y��&I#����#:jK�J��W��L����.��N��߀_�U���1�FH)�N�Cb�m� (~���f�b݀*��2�r��G'":P��ODri%g�ҏ��j'N��e��g� �]����(�B�fl����y؟��	%�(��Si�4� �D��D�|��d�,������[��@2����^tM%�����
��H�:��e<���'sٛ��S��8s�d� 4\�I�6{\�aTÓ�O���n�}X�X���kl�%Wy[�-k�}N���%��b�'`�y&���.������0İ�5������YK=*:�����J�����;�x����\�p�!�Z����F��%s���ͺO"�⥹��m��+5������o7�T����z��� V��w�U��	��P-2�͡���[�)d�f�MCϪ֫;�?�U��_S1j ��\�W(U0���1@�|�m�����T{�W��3	������y�vP�ϋ^U���5V擜f���L���<|9D���IC�yg�V:u�h%��7]1N"Xө�Wn�
p�MSn/o�4��%�ȹ5߷�E?V�U��񫨀��|�6���S�����V ���3��rT��v��ɚ�R��6	�c�L��g�d�3O
)#��q�(	_"�b�v�BY��]��%^&[�R64X:���/��n��~K/$�~������������ �  o԰*��x3J�U�$pCw���	h�����WWPe�jL�1$���6	#����]�`�X�1�`�	:���N��w�h�3N��&��o�G!�|���A��	��*F���I�W����	]�&�m������e���.��9i�����`��ҵ{�l2�v��7:NFo�%6����h H��.X��[=��Z�>Q����6��0���8N������mz��Xbx�S
릮�M�]
�r Fo��<z�eE��
�0'�K''�˧�7�p�u��+Ac$�[��hH?�A�_��A���B��=���=�2���Lú�;�j�l��&F��M�%�}֏r�=0��$#_��X�ߒ��'h���6�}���xA	��ga!X,���BYuXz���-K?&��y�׮�˩���?�bFv3�o>��A�q���m��wkЊ4O��y�K~#dO�<�c�"M���y�j�f��I����R�,��Gh�Ve��O��$q���i~?���C_/R���y=��6���eD�>�k7�8�Y�$�Xb�XB�p�ȷ�39�*�յ�P��9��kSd�vx���_�r���g\_�tP��M��%f�����èh.�*�_��t�Y��M���*!n����*|8,U��l��Jf�l�H42�q��x���=\q�<L��Zu֫�n�EKg��Ⲟ>Z� D]�%_`X*���G�!~88>P��?�@�BY� ­�Ef���-N=��1��n���Z�X��=i�Ej�d%�|6�]u�������JPO��m'��F�؂��,�s��p���Ka%�%�F��p�4��'a�	`�=�;h���Rj��,~�

���`�
n������"1��U:j�g=Oc|�Jဢ��֍��Ԅh��l���.�鹬M�������N�-������4f9�W�+�ӎ��K���ڞ� ��Q<>�w�o���I�y�yP)3������h��Kv[�6�e'HE
�* �Ji�Ȃx�>셝V3ܐ��)a�y?�}Ӈ}_Jī&MBLNy�7�����4缎7�t�w��{�G�Q����ѱr����5m�AxiX{�������O����zu|�	���K	e�"ȿ���L킍U3���l��Y�t�ԃ[���*�����,�۴v�����U+�9y+)��ȼ���L�ʴ2o���ݨ�����k$��u�,�2��P�b@t9��ikRc�Ơ=4�G4���%�Ջ7e��k�?��hM ��3W��݁�ǚ�C�9$!��&Q|��I�$A@���f��f@��0>���&����~')Vyѕ�b��8M+O���Չ9G�ؿ�P�&�ַs��Eyt���� �Y�&�;�R\W�̫�Ӓ��0��p�E�Ci���*�}XsO8p�]itė�	�.:��$m�j߂G1bM��bJ*���!���Yi�[_m}şN��Ps���Pg���J/�����es��m�����rKA�9�o���H�X�k�c:��TM���j���]zbM!��J>���a��j�YP09h}81�6�.����o+�߰M�y�{�)��)#7���u�gA��L�nQ��^����\^�3|5�r��Di���b|w�ѣ�����oC�	��>�󵧾ǝ�>�à���t����̴r_���WD,�­U�[`j� ��W���Ԫ�':�O@կBRyk|�b��d`/։��e¸
�МfL�ـז��lsF5-t�K4 s�&G���1&���u'�@�2ȡfYv"�.�����:�������K[.�9_���ntcNֳ����"�d���+n����d<�h�^��!?-]Ӝ���}uT��2F��]^
��j�]�xJuz�ƅ�W�XㄦK�e�wn������O��#X�w���&e�<��k��ϣc���^���Ild�-�!ҁ�R�xUS�Fj�'gI¡�i3��р���dS�� ������7]y
4g�iF.T���:�yS���f�F*�e�,&��^��A���M�NӶ��8�l�qQ�GI~�\݁�fO,�Im�,��6��/���|�*��*�Y�JYQu�x��^
�l���񿃳�u�^�AB�O�AM-�콟���"6���5��YhZ�����F�>�\�~���&M�k��`(�Pg�Mk��+3W~羱A��Զ����_Pr固 ���H��+�- ��Z��Am��)����>)��C��܀�o��T(�@CA!���&<�������	$�d�xb�scS�i�A�ڵN(<�X��#~�5�k�����O�����*별�W�sF����U���s��������P(d�8�A��~�b�KA/�غ�|�Kfg�#���&��cw==���RX�C:a�U[���Ӂ���"��~ic�%�����2��,�ō������Ɂ�[�7-=J6����`�&�t˟��#^k��^�#9�.{���OnX6�����D�X�MI��2\���]��&����7{��M�P 6����ȎV�RjՌ��݋��;
���� e,6�?��	hy��PZҔ��U�x��N��:m8����������Bl���z�ŋ"����� ���TQ�{(�>2%_��1]�bq�>�K�/���2�H\^}�e��vF��d=�T4�/n���Xf��o��YӒ�/�Ơ�Q�,�.1��1���x"u'F�ehu���R�'/�7~*��MA��n6t�������7�^�hse�,JzU�d;��}��hhI���;��G�F�� �]_m&���2{��S�hE��FAa̡�.&�Z�
\]�1�J޼]X��X����ּx���e!v	��-Ի"ޗ�����B�s|&�>5f���#�G]�&�u�/�>�� A��a��MS�[���.�A�?�[-�*��<,�^���`����{��*�n��&\ֲj���C%���I>95��:���M�k��IW��?�S�{ri�AM���D�c��.����G<�;~ؔ� �By�a��錅`��L���Jju:���,�$TZ�`?N�G{U�D�:�a�9�%X~����$��M`#�mg��~,驐Q��ӺR���M�6�MQAp�B�Zw�I{D�߮�.WѐQVG�96
I6Ƥ+��J�R�ly�bW���F�J
i�.g5���t��j�����C*ewj@�?�\4���4ïs���)�;.S�Uhh_�)�	�,������{�=�%r&:Y/w���n;�rS��i�P������{�FB��Oe*{�D�Ԫ.a3k�C�11t�p�I�Ѿ��$X��B�^���P'�����3n8"�yK7VUF� �2��M
9.�h��].�I����Q�:�9��X�P����3�M���Ρ2%��O%�6l+�,�%Y7���v6[J��[�r��W��bS|��D��Dl>�M�.�c1���+�yF��n��Y�jӢ��M�W�W�W5]��\�IH�_X=�D-i8mR���FG�w�����Dv�f7U%}6��ʃ�x�S�3C�
sk�k�̃�u�si�R�� @�^%՞���D�S�&���_s��G������|^�js���hV��rĀ�fa�ݗ�^`����)>ǀ�YG��Xv5�	���I`Y��:����cB�Fz=]]'��Ш�#��������f�VO"�����`��ؠf�+�h��(�O����@I��v�?����ӗ<E"g��z��*�7��B�|_�L4<3��ۺ�Z)�B�'s;�YmM����e�rFs����k��P��M0���A�Z��=t�LUDF!y�ݯ%�sO�x �=���l��2i�̜lâ��ks%3�Ŭ}|�o"�U��"R����yH�g�Vd
�Y�ބ�Q�łkQ���,:06L�s�� J�2Q�O2��HA�Q�7 ằ�%YG���/蹪߰��}5R�7L�R�3K�N�l)�zԧo�����8x{2%$pQ� �{�,������K�d�`W��΍V�ͩ���c��#}��0ڥ3�\���0	��ߞQzcd��e�i:;�B!NQq7�(� ��op���)�)����0��f�n��3�)F�[/�:���-?����?���d�3�N ��Y�nHgdmP!�&��!��V��zA��g� J��<�(�k1	���IWmKR����*����7�?�cA��Ǩ��9��)&���gk��#�Z���ݩ+!տ�m�A5���c)�\ZnFo���=1�j�(��1�k�^g�J:f��I`��qx揧�E���N��]�B��������C�N��J�u�ڳ�q��K��jyd��|%�ꯛ��H�����P"~����I�<Պ�u-4��#'�bN�qZ�2���T=&����I�c���͢�S�|J��z� ��@Ƭ{f�
7�T��_�/.�u��!�R��Ūb7�S���������8�@vP�6�D���%s���7JH��!��v��ß�݉�Ĥ\�h�"G��+'�hҲ�Pu��:~ws�Y�|��2!�a�4V*L�*��,��쫚H&E�[E�\�f�ߜ:~sd�ė�����00�A-|,��u��bQ�Z�bO��d�Ff� 3��a� ��qED�˗Kn��L��`���M\MYK�V����W##��#��|�8��rl\w�<�ΗBs	�C �-�� �X{��C��V���uvq�9:�O�k����v��=YgYb��w�[��L�k�������mF�=�D;�gN��㑒��!��c�G�Ε�����_�?%b 1@���x#w�.����)���,����{�!���<�'1a[�;Yί�~ɴRpE%<�hPlcJ�����2�	�������E��wN|}�>E$�:t�'���'Q��L�!j��q[mf�ӤGIߥ��Eb�RDnTn�rl�CͿ�$��ĮVD��S!��9���$B�D䒤��vŮ�΅<"�L�܁C�1hI1�L��^l��PX~��H&�y�Ѓ��cӌa$� ��b'���o���#����J�2�Ui����J��� ඵW�������ϔ?qE�NO*�<NbD��F'�v#��ӣ/N���f�܅�!+ݜ���� �I;�"�q�u�i0��� Ք$�o��l�мl��~�!����$��C{�vZ��t�F�j_|������?�����P2�Ӕ�M?��3��µ�'&6�?��D�:����Y�����	BI���n��4]��ی�j>� :��DO.��CS��7�,/�i���洩H��e����*�S���˥����ZO>be�P�`�>��N�U���9�ue�G��MV0���d�9���_���@�dC��]|�$wc��_��)V���*��������(8���Q�:2j'R%��Jt��Ѭ4����?M��Os��H����\/�i�B�RN��||��Z�.��1��i�p��ڳ��V�L��sM��^�hG� Y3p�Pâ�}�����I�G��2 �>��� K��;�SB~�}	�6@��[x|B|5�W!@ӓj�=��O܌�)q��y����7��]>�@���������0���	��[��k
Q�p��=cm����bn����������}k��/�h\(���9�G�>�ү�8��{���w_�=�`:)͑9����%��!�s�`������}��#���Eg3�}F���ar!
�ޤS1M0>�+����<�����SWM��֙o1jܳ�Z���@-g��mk@j���MK��A���=GH�>8�b]����7	O�[�/������"�@G�⭺<2�a�Փ��x���Ǐh�����Nu�b��:���N���7�˸*OJ���7�����g9A�W�����0����,(|�ס��屆�<��d����:7�h�����F~ݱ,�Z�Zl_m��{��(��Z<͚8�}��� D�3�S��"_s��(�OZ�"��d�ޟ-��_`�myc"Fl-�(�`�������<��xQ���ַ6S�V���F�����O���K��^�g�>/`� y��j�?]R��2&@� �j�i�;���6&+��Z�T�7�Z��r�}��
w^n��S�ʟ!��]��?����K�F_�=�������U{��єf"�b�m ��zD����e��'�*+u�5.M�:x8�3�|�+,H�[;�ù��ʷ*�ӽ��P��$��)v�+��F�d?L�DLk�6H|��(���3��{�� b̈́����"��{�#D�.�o�a��T���%fH<�m�������EՊ�4?U�'���t��E$̲Li�ԄN�ӬF�����k+i:2e�@=3�oa]5�����K�N�c�����S���]�[t��Я�oEr�Ğ��M���9J�<oz0̵����y�d"�CMD��Jy�#����:�rn�������/��{��(hʢ�*m���M3�g�9�RP��_�h��cf<�oQ�Y��e��)�Ɇ����ݴ�.�8|#-��	J��G�E~u�=@�ܜ�?�"�����yEi1���?C����@�C�Y3�/D��?{���z������$ȸ`��f}46��H+�w>VF
�4����Λ�Y��<#�q�K����Ĝ'c�Y���rG�=C}ݔuH&�[��`�L$�1{bW�[D�'M�� n%/��S�AO���s?�B�&�%��zY� 9�R�-��Yw�[����Q0��V��
�|�X$�2�6��U��Q#h	��}/O�`�Q:w��'����Kp?��/���m3�t�;��%�	5=��;=:��x���1�*�>I�A��Jk���nb�i��^Ub�>}x	נ���q�Q6!�>��:���?~#�04��"Z_a0�y�z�=T��;�E��!g���)a�1ie��F+���>�)�c\�2�~~��)R��stLaխ^'kY�C�W��}sYc��k�QfjNRkejq�H>��|R���/R�4t��΅�n���������B�3��#I]��W���'�sA��A�h6��u�p\ϜֲP��0ˤ�����j�z���D���U5t��T~H
�1�u��$Ӡ�欱�q9YYd����\K�|&ce&]{Z��������iM�G�2M�A߾�@�7#�Ra�gn�����|�����۰e�T�l��sw��������sp��%ہ�,.�{X+�^9-��7U;`�J����e2�z��<[k�|KkV�{ڱ�u�q!_2��ɦԵ��ǃ�5����W�q��������+;�����T��i�RA�*lX'��K���^� wؕ���:{P�W��E�2�v�)>�\�G�~���k�3�� �l��J�A ��?9�J�� m-�5��0]�ka���s 0++*	)����3��O�r����#��M&�����t�X!҄Ǝ��ß�Hb�E�p�+�;\��C�Q!w�Rv%NN�؃��} ���3z  $4�a@���f���M>3��W
m�U'Z����1`���$XUƮd'�!*Nu�K�ݏ@��_)��mbE@�,,�������X�Ic�75�S���#l:��3 @�#�p�M��D8���D�ˏ	�XܸI��@M]2� )&�~8QY�	��]��L�]�g4P�vٯ{�W�18��ܲ)��LWU�ƛ2|׺1�tEG=���(Ww���{���`嫋�S��E����00��%�w���&��!�㠗#���:�ze�a��*��5w&
�r� ��ٺvʠ�h&�&�Y���3�&M�`�n^�ߕ_��t���ڶ���%�\tK�^½m8=�懶]��د+�:�'J������ٓ�I��m�Ũ0?&�~�݅�7O�iڙxo0����.�u�="0�z=zu�C����G_���RڀɆ��Ȋ\�G��^J��w Z����7%�K)�+?J�0���Pf�*+�7�t�����&��H�C��k����jS�d�A����pU�V��Mߩ�} &����U��u�-V&]�l����WL
{����m>�����Fjy��w�Y�������� ��5s�I"&��Mt��{��S�(n9�����>�;�j�U&y��z@"%�B��P~�|ۀ��e��
��N	��} �V�輩�(�U���Wf%�y��t�V�r���ء$;���Ӂ������
df�c����qp��E�u����c*[���ɸ*rE�0)�X}�]�?391J�&�Yx������@ 9A�A�K�����y�T��jx������=��%,��ݥx� �Q%�&�1в`;�x⾨�3 ��/MH%����6��*m|H���W=K$? ���	��5P}-kR2$3N�n#gt����+r�?�U�@i#8'ళ��H���#�$�� υ��N�=uFΙ& ��^_�G@�����A>=GZ��㙄W'(x�x<���l�\3��F-P��ә��P!b�s��$��j]#l2���?�=-z�)b/< �c��6�ۃn-���u/?2�T����^�7FT��X�{���дF�[��e����M齟`��n�i�	6��ݽ&�/v��~RB/=��������܂�@P��`Mt��+q��J�;�tô����6J�6o���~+!\LRMܜ����ߙQJz7��XO= �m���I�LP�����?ᒞ��&d��>9�+�vbϓ��̹J�q��gX|��:�	����Hm!th2�`�B�U�j��x?
��D"��z[ehG~_�\R��5�9>ܙ��U��g8��	�Z����v��! Fd�S�'���'���\%�IS��\ C $���p	:����}�bl��$ٽ.f|3��a�!�^��тBL�#!�m���%�5�ʙf�	_X�LM=7]��C��޾�y�h�B�N�8o��*�����b���9�<�c�E7l�!O$�S$��ã:!y?���K8�y�,(^JZFh�E )X���O�!�K���*h��A��; �^W��@&�������aÉt�L��D�&v�u6���er#o�:+�d�C:��(�l((r;���B��Ue�����+���^�{��� [�V�=Ġ�h�Kx1�y��`��հ~2���b�+a�X�Wy@����_3jA>��I�̸�#�����W�nI�{tyl�j֐�?�k����E���*h�!4j)o"���_�Q� >A�R��� ��5_��Jy�����@]�+�nxl�h�ޫ���v���c�l�U참1��Sg�ݲ�շ��J���J�AN�FP勃>�yJ�U.AW6�N�jA�<���:�y ;D%� ���[��>Ͽv��*���o=؛�w�um�z��e�~8qĚ�l�:�b�z�޾��4�o���³�D�Fɲ�_L}\�W�z^��b"3R�|��~���^9`/����P�C@���Oɔ}n����}A���v
���˭q�H��MxS �����������-ٶ)��Y�Vyo�7��yK��v�/�����P%�����r\�OZ��:��H�(�}�_y1�x{��w����65�^�Q)�+N�o>�_�WHư�P�*�^�ƃ�y0�19��a����ے0���{CG�����|�5����'̹�*�;5�<T�ϩ�WX)Ƅ�x�����!�Md���5�(��A�����U;B����ɦ����E�s>ª�9���4�VU
\@�E��V�f��z^dD�Y�����I�[8�X�Ib猾�� �QMd�Tc�*�u�!ufl���m�;�|���͎�pMU���]3�b´�?:��~�v'L�^�ۈw`8��1E�0��~��hY��yx�"�1�{�^0IKf8#{P��r�>b�aU����%oax�V�z˷�ɭ[g=	��{��q�����fs"�t�3�\L`!_6�T��1Z��9��0y���B�-}`��qd���D��B����ۙY�J�/U�g���6{�~2����Wװ�>z�Z�����Y��mDݶ��2]T�җ��C�~<�)5��*���n�V���i;ƨ�3�f�+��r� ߌO��U�"��N��:���Q6���ᄊ��7`.Ր�t����g��
]/0��$TLTի��~�o�]�[\�F�y���ME[KO���)�{�4OJ�As��F��<�Y��[b\ZNp^��LaP/)J9GY7��z@}�	�M��?q�1�V>G�G��_��P3᱇FS�`c������ �f��.��l0���9Sq@}�1MD�5D;��.���up�h9�|�#`�w�R;o%)	�C���At}�!5ׯ:�'� =<�N�,8���4�ٰ��������$:�6L��A���` ����H�y#��PA%Q������QJ����b���H�K�pm���@�A" N�~��C�b[g���=H��a[�$�:{*��j��z���3�*��S����8Y+���/0���:뀪��'�[�6��8�9//�pf/�P+�g��|�u�{��/����uë��&fU�2������}Gv��h�8r[ү	��mk�x䪡A偮��f�{��#�P�Q����0s|�v�n��]3:*��
�ln��t�f1k����S,��apM='�)��eQ�CP��;�c�������g�,燃��O(����H�X!M��j���x�K��ix޸x�����r�
	�+5�h��#$��m���B֋��#(/^��9zP+�Ī �<��K�(!�~�hE�#��ut9�I��M��g2���S��u�PȊ��f�!~5�����v�������n�G��%��I�8�|i5��ᘦ2�B2��[l+^����L�����%���{l�'��x�.��H��v�����2��rWK�A\�MTě�U��uPC�6N��2>u����/������E?~s-�cSݳ��!��qu��b�̣*�&Y���i��×\�,�)2Һg!k�E�Sq�%��rC���c�ۺ����=0%���yI��)���2�C�I��**�q�!Bf������S-n��_&��@'>?�w^�@�`��h0WgZ��WlY�]���+#,������83���H�h�M���Tr:U�4�9�*9.ؐ��'���t��7���3;�ku;h��t:�mēoY���a,eǗ�|��gVuș���_�b
<�Mk�˼��Y�S/�<����Du<Ks�yHt��O�a��Pf�yLB¬kO	�C��O�nr���eHtK-���PC~�z:fe�j'*��0a~-J9\�y��I��О���N�wk%�Mٳ�Z@�X�"���9uX`\�^e������A��lDD�7�b�v�����B�2��%ϵʔ��!|�8d�3�0׌]�+qޠ ����B�̙h�@�U�d�	��]@j�ɈGAf�Φ�0.`U����S�m(π�$\�	���a#;�;u�9|ϰ5f1E!�jTY;�U�u3O�F�$+�t�h^�fI�<z.�©(�v�j���T������E�����Z��+o�ް7"�U�NH0�X���A����~�Y|�X�n�x$KA�uA�'B1*e��1z�Q��Ү��`9n�0�·�'�A֥��3�:_e�����T�Q�[�lns��%7����kIQaj�t����|1�a��"i`�n:�$�¹<ax�g�����&uX߇���x�$"��wz�Hx�4 ]S^��А�`�H�) E��t��.�
�v"� p�� $�����!���Y�*f������q��u0�aQʙ�K.�3�h�����0�#OD�N'!j�@��yS����ܥ�A��ͼ�C(1��9��{�ytJZ�))����x�j����c7�|�Vf���ܘ(��}�< ��O��j�&��z�Y �0P"���"SBby�u	����!'�Pg}
�,�oO%�-�^��Q���P�w�r�:���y����(QO�����Y���O�}��b���?%�	��t�3�Z�wv�r)N6Ms�������0W�7��@���Yp�oK�y�k:�VW�c?���˔���zV����⒰/9cO�4��e��M�g��"2�"X�ZEܓ�4:�Tr�u�Wrd����#��%�E!+b">l*3ǧ/��^N/�6��M��N+jo���XT�ݺF���ήy�A��#���K2�� ��wMy;�����w�<�6�g��3�auX��%>��8����E�`�H.SAKz�͖̟��P�8����Y�=���q�.E_=����B\�雰���&�B�q�L����W���.�E_{s�'I$c1=�e�u���u��/I�
�Ir����/���PҋWΝ<��2zx�=�mZ�[r��w��1'�	�\�'F�*�.������犄�[21g����{�+��SӘ���j2]�(nG������
�~1k�*E���WuL=y�l'=㚴�{
jN>�?��I��v,�c30���%�sR�=P^��1��qF�a錚AGr��D�`��T���\�ǥ1���k��eA�h�Ii�'��4J�6�*w�9�nK/l+O��
4��ȭ-_t�+�;����L>���-)*��5W��Xˣ$)]��WVzj�h�������L���9w8�b��eeL]��	��LI7�:i,'�����K�Z�,ny�ym(@Q�o]1k��ͯ�⋪{�r��z�}aY�&�HD�:g_s_Ü�痕����_�vEp���h���lw�����wp�k0�k.�������L�Bn>?kI̶Cyr�	CX����ռ�V�_5H���bfl�'Q.0gB��������f֡�7�����h�/�ž�{�W�y��m�=c�I7�-�r�ڸ*u%��tݨi?{�1�m���^���a�Ip}x&#&c	��ʋ˔�7�OU���(}�YdM�rz��{y���yD�	cW�F��`�e�YBID�S\nog(?�b#�sU�o���+���L|.�aA�����}��h��s/_�чҠ�w��b�Q/���He���=�<^7|b��)�e�]�o}���N�k�(I@�3,�tA���QȤ~�_1f"u�۽Ŋ�&:İ�v��J�b�$��+�:v��`̅�8����a�%"��S�.��4�ڄ��_��P��G�2%<�aAk#���=�#���������Q��p�����7����Y���A/ͮk��
��c/������$kJ��ڞ�=(�{^}�;������b�U��0������i��yS���_�ocga���8�m�[�<܎�֒ ^��������k�+� ��GGk��$�S�/9�E_o���i2q�ᩜ��?��W��K�M���I�x���턜ӱ��?L��5�i��
03f��W�r8�C�	i��?QӕP�����+����m���E#���{��{s��F��x�hR"�+�ϭqBD�5�N$\��[�­�n�Z%vj~���|��'���p:`
Ӆ*G���
U(�_X���w.s�'�-�p� \�'��\�M�/��Z�AE�;q�,��
S��RQݎ�w�{�o{.�������J�0�x���k��O|��r�²�UT-	�f��b��9?�����!�Y-�J9����)AU�W��쐯�k]S�O�q6���ҏ��iu){�c�~wA���9[�*:��r����I���^��@oP����7�oIJC����jg��Z�"�#�ׇ��SQ�j�8�7>��P���K�����lp_�I=����u�WfZYȗ�y���'<|.��u:��h}T�ts]0�d��
�h��D's@Q-)�G@��6�#������#�s��%)�����d�e�$�_F�����|i��2���v��n�x���#�r֒�gS�I0يLdR|��>�>#�G�h�G�~D��8�)�]�(Z���� ��Z��?̢�*�!*�,�
����.������
�I�'ˑ>aN\	��}
~�	O��X\ua���[	F�k&��OEb����t��x��Ta�������!�5k2y����$4V�l`s�?�st�ܵ5?���5����ygWYY�5[j���#�N��;T�6� >��Q����C�|I�VV?XUtMY޺)-��v;.VK�`c�#?�=� �7��Gw��|���x�jGA����,�����;)���30O�x���عcv��w��V�7��^���ܠ�4|�=���hFi]��D�I:b�)om�)B'��ӱ{*C�H��+Ƞ��ޑ��)c�`C��	��1����&�`��$?c5?W�����wz�Gm��&�&�-�p�9�?|d/狖�oȐ-l<�����ΐ�j�[��{�-j�����p�>h�e 3�`?v��k�qГ,��6SӰ�2���\��|�Me�O��8P������;�D*^��t�ԗlB�yBup�!��ӌg��Ǥ�Sw���4ػӗD7x�	������ˀ��,�fz������p ��A�Y�]�af��Th�E�Ln�* ���#tj��L��G����]� Z(�S�fVT�� ����䴼 �vQ�G���"��Q�N.�k7�H/�C�F/"��z���{q��EYg��I>4l
9	��65���_�ЦP
Z�4~�����;��q�h��K�Jr�Y��3_]�㚮��r~���[H��g�7�]iٚ�
p���F�S��u|�r��{6�:���m�/eU�Y__4Xn|?�ד�Y
(8- ��Ѯ��Ԉ�F�[���f��-(J���{�Gҡ�s&*>���@Qq/2�7�K& �[x�l1r��{&�8�c��:��BۜSDFI��"�T�ҏ����w���$J\X~O������E���XΔ�(�e���=>�z��FFC8��bw\��y�,u�����%x���@]�m���I�il���r�s�#�L>~܄�~B�/�\vƷN��Sޑ�Ϥ���#q�����Ǐw�z<�X���D�a^(�ba��洁wH&��q�B�~k5 5�c��dF_���tg�����p/��[��̙n�Y���jX�Ɖxl�Z&�3�g�2��u�^T�>&�@��}ϻE�o����+��<QO:9ՙ�eF�X
�V�� �˜�*��p�\��]X�#{x[H�u�^�1��[��.f5���	�J1]�aPI����� T�[�Fn�q:t}BƘ��_���j=[��_�їc��O'N݄9�݋�Ce}�gc�}؏�|	�d���L���x�$�K�_�.�����$x�B�3����u�-t��6���������J��7b�� \��~v�iJ:��k���L�![��I?}�@in]��栓�1���W��5����'녅c/m�އ��|��C�Y߬�)`R�ΰZ�e����^�T���������o�cR���sY"'��k����=:�Ɋh'�H3�~��z�mdg�@1�h��)T�w=jj��`LT���F�'�9صGU�U&p�8Jêɐ�`�E�+��+�u�[�2k�x /R��LP� �LB�	��r����s������zn\� lh +�R� ��W,��6����G�H��:�F� 0�t�՝o��)u̹�����q��53wtDڧwu�y�b�a<~�n���X��갊���#��G�[�?�i88���!�9+�MZ5�MNukʖrm��{�%�٩/%�{�\����<4~"��غu�"ZZ"8H�I�8U'���%;dM��P׾Ჷ�߉��sWK�4�=v���Eq��H�^�N��N��hug('ў}OP%l��N� 0���X�K����R��90����Sg&�@Ei]M	������G7?'Gp��U��NW��pYԮ�;q�0	��f�nq1��N�������aC.�1��-q���*�넍�	���-���!f&sCJ��Hp.�g^D���l�(Ӈ>����=�ܝ�O�V�?�p��ZM(�!՝ 4��x�M:���&�h��Z�?���/X¹�c�������J"ߖӲ�A{װ��ب�oha�jlI߾O}�jJ�Y=�8<0 �������]�e�a7)!/�NԭjM@.���X4{��E����c7��B����6f�{l�����H��L��O�>x���/��=��\�''�-;3e�����R�ܱ��po�>S��a�̣����}S��S����.yl�[&�D�5�\�sz���������w�}l�!�Y����1�4b(1�_kI�W��x��gU�\�RW�%pE�Ӛ?� ��ЈP��A������0�h�@�r&!?^xe|���/]!�N/�lM�mV#��>�VUP����`��-��L�}R�4�CZ���?�M�P��6��IZ��f7�̴���6̓�#"�Q{i��<�cyi��Y��቎��������Ԯ�++!gp�.��t�G�P�d
-���K�@R?Q��P��ݐ��j�*H�=a�-��-�8�g9�
�Y�K�j|_h��ȼ#U^�BA������G�QOtHҨ�x
�z6+���v�L��$Q@�c]$�:�ª�퓂�';2/�H�>�hJ�3;IhGr��PUQ�4�j!I���j�FR�]=#y�]9�s[�����36Fʪ00Ɂ}�������P��n�n��"���w��HP"�2�04��~Ȓ0�?ņ����������
c��!���aѵ�c�?��2ˀ�U,UB�^�Kc`��:s67֢������J����Î$fĵ����+��珸��>s�N.�&k�	�d����#�z�~ ��3�ct4j�*w��ɗ _,5�)w��#a��%�az�-+�p��
 �w��r7�j�Z����Ht�#E  ;�ֹI(m��:��npIJ�}oK�4��
^Ҝ2}TC� �6G!h ��- ��L�Ǭ����}���axS���0����+�!!DU��0DyIo�k�Y~�v��-��iy C|*��
�e[靟07��	l"��_	�w�� 3wvq@������߰��f�!��CY@�Vo�u��$�B�r�$��0�!�+wC������ׄDl@�Vf�􅂏lW�M��2h��fW�u�.$�lk^G�Xz�E��0�V�h���������ʚ�S���5�٤F-��Y/k�?�U�4*D�F�STq.��e�8�J��;]0_������~ï�AxJA�GA+-U��y�8'"�yϚ����/��Yb��7�������\Rp�P�X�g�0��C�X��zi�>�PR��eӣ��p�.S`[i�>����~�WW'��w?�%�E/_ƨ�E��pU)%0�gy=����t�h�"������oj��=�/���tP�y�U���h܌%+{V�/��T�"�������I�d������u�r���S��h�IW K+hKx{C<�vI�7�h-�4��-�/�sC�9J�T�?�9'�΃ne�C�с�l�tAl !@�U�x�������Qc��A6v�7D���1T	��?���Vf�0��ŗ��K\������u���L�G�A�+��!�|"�~�$FzU���x�T��N�	�����a�wS�����wB��>V+2�]��Qs1�m�%��<���8��E*>Lpu�����?�9O�4��!�x��#�
-v�׍c�[M�Yq�������@'}�F�������Y�i�^��6?��	����ߘ1�� �W*��S?Nk�Dy��T�����_c_���>4���\C	���ڤ%��'���>0�o�WT�Sp���Ե֜ r�6o�*�r "ˎ���T���+݈�L?�l��8G��E��zvE���ߜ���z򧞶5I3a#�츱� c/c�Rϑs ��:>���#͉K7� y����"��\�Y/�O}k�/	�������_�󟕲��W�od����j@�XOo~�t_���`�'�rĦ1�GY���FaB���@����;�;ʱ�]g{��WXH+AƟ]6QB4r9�-�I�o����w`�|f|���5���S�A��*�4�EnA�A�	&�_{B�j&�ݽۊP��-����Hxܯ�8~_s�����u, vai$vM��%�f�v��7��,:g�jſ�# $��+\x���8���O�xl�G��Z}�QppY͖p����u�'%����&�
Z�!�	�U�t���g�<�H�ZX@�L~ޕzN�:������+	��e^�3���0E����>����Ơ�۞��o��c����Ð���?���tm��j�{��<�"��:eM��x���mz����]����fL��w
Y;���E���9H�8�K|p���7�!o_�L$X��P��!�RJ���~<z�G$�0��D=w(9�b�y@��C{�M�*۷xL^A���8��B�l"�E��0Ͳ]H!AR��:d<V<�и�Z��Nʆ\-mJ�@�Z�i�Fu~'�➖��#��¡v�ld�9��Q|z�}Гզo���K���T㖊)�����e��((O���?o��::��ة�8�����l�ˇ�\l'�|��k`jh�^��-���5���i0�%���"�J\��?�������M~s��ͼj�>q6wol�h�@���F�����&��*�7���;˿ޓ�k��ʌ���7`)�ۘV�΋+LV��4׉! �ōcL��:��� K��-%���g#Q.�D#tO�?�@K�YpCv���(�o�|{f�C�B��6��vKV��E���� KOd�$`8�!+�w�k���\
֗*]z>I�9�!�u����H�R2N��9W�{��I' -*�t���7��@ȼ�����g�C:vu�MH��^h�f��	�-�E��Pb`e���,�I@��W��,K�l�$٦�%�RN/��xb�,�'�X��^t2��x��h�3�|Y!ep�Q�6d(�������Z��{.d�Oϣ��E�uцW�K�+�7/ѕ�����ji�r�]GIL�������\�����x[���Ӊtp��K�s7�0� ��Y��&{�Pп�N�����XT�䭚"�pUNd��bPY�ym���GU�m_�΃Ġ6ά	7:#\p����KF���ख़�hM�JA�;*�	-���M.^��.h�&ܲ�w�+�{�7{GC̗>�an�M�`����%WlI�����u�-m��ȷp$y(�u^\j ��f���Tf�Z��e�I�J�!�3��\(J����w\T�x�\�����ҫ�������I�^����ν)�ţ���$4=�(����b����!����&+�،����S+��9~k���L��nGLT��rDC���d�����\��*����y�(�H!
bZTD�-K�ܥ��ٰs��-s	��hM�gs�3p��h0�� �����ϙ��*��'�2;}�X���!�-��x'�ke�.7L�D2��:�]�f�ʦ׳q�Xh=��V�����Mɵ�Mָ�O}��\I�������_�뵏 ���������<H�Ru�:x4M6zДg�]�����h��
0#���7)�b������w���{�^�L��ʹ,���7A�$�R����]�)���k�.���x��Za�霌�pU(���D�Y��s�o��!=�CFˇ���B��C�Shؔ�Am�N����aǇ����u+c:[LzH@�"�{�:��8C�@�b��u��%Dˋ�.�ͯ9R-ڞ���il��Fc�a-�s��yxFi	�K�[M��;�޷.��/�Rۦ��` D�y��lR)�;(
���dώI��Ŗ�ϒ����l%�<��,���lJs{Ԛ��x�9л����!��,�5�q�+�H<Z�d�$s�A-�ꁰ��/"�lE�_�a8 �三.;����SP�:��n-	I��JI�N+}$�q�:�S�J>t|���E���]��G�Vs��
��J]�SOM��~��}af
�/�ae��w,��B-�S���0 1@	g^�㼂2�FXg���A�<��ͷ:?K�H�O=W�٠~�j�$/��{�X�������[�+;�	�6��ix�{�(
X���Mj�N�zM���T�� ~���۠d%��
�B�.*����F��[ݰtV�"Ξ�J�]� ���B:�n���;��Y � 8�%i��P�g�!�ē�L�g���)�L�K�~^��{��`�����]~�"��Х�ҕx�eF�� �,˻�2�Fӥ�3+��
UW� ,)��?u��f��>��/���T�N����G�k��T��ö_��3cG�����V,#͢_^'ͳ�,�o|���A�UD=ݥю�^D����7r4@�ۤ
�*۬�p@�s�����XT� �g�(uB*�&�P٬��1�GrO[��}=S焨}�Y�!v��C�}�ޓ�Y��X�����֖�/�?�m�d)^�e��
"�N7**��~�D��Qn��6WT߁��Oڙ��� `�H���=u q>�xc�pB3y�&��ĸQ~
���$*�52��\����ތ�W�F�'x�(�z^��F>��`�1V|��BHW �~]/�R��Dr����X�߀Ct��b��)�R�'������b�TRO��!_�)Jڈ����)~��|Fd���<K���*�d��I�u�݉!X2�#�Y�3�5聓�z��t��8��K���u���_k���B��R\n����{��%�Q|ěb.�+�/�[-�&\?�!�>N?���^�A3��Z��V�ofp���/U��5��hxq�1�ɶ�h�`�P����tݞ3��Γ	�n+VGv����&�X��X,����Wa&-�������
k�#W���MF��<�%V�I�Db�rnoǗ �_S��?c�|`f���fP�J2JTUK��5���y��ҷ;���|���p'���H9�Z�i:�p3����ۚ֞寝�J=f�{.��o��P�h��}0�g�*qT�~)1�La�D�=���Z]�ȓ��[������c�Lb�n?���Ó����{�''�xw�n��@)4G����ƇӦ8���ʝ�{�ː�i��N� V���wğ�Fn�z�s1�	{�4��^�è�o��dg;Y�a)�:�T�/�3�*����w��I��/MJ�sL��aGx�o�biH��6�tg�2ưN�~3
��}��0�3��nbJ>���۩[��9s<��a>R ��;�c���s�5���vy3;�D��Q,�g�S��~��d)��:�\
��s�#3�m���&I�@7�y'�]�÷�B�W�Ҷ���`�M���Nm��Rc��z�y����J�>Ĝ��g=��G�IE`l�ү��=�B��2.�~g���萠<W��fl�_'�{�状q�Cͭ�������٦��*� ���~u
b���e�B�;٦S���`�~����F�J� �/��ڛ��U������mE���	��Wy<��%�;W͌n�0���&#Hx鹔l�8��O� 3�Ȼ�)C����>竺u�$wO���&�n��d���mm�*�$φ���Q�!n&����0��,݈Ĺ`�����q�,�w������nJ&��<�]�n�טt�&q:&�h|X&�D� �[��7���a���Gߟƽ
*p�%ѷ�>�MMU��?$�͊��{^M���Q�cH� ����%�����$����w�C��R(�=z&�����\�1R��I��5w�~�36u�W�Ig��y\J�YA��Nq�����R���x%V��?L�S���@'e�鵝k�z�F�_�{fP�S��kRI��4͙lVP ���獡�<Hę�` Y~"Msɩ��f�����S��