��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���N��`�G�?��Ɉ8A���*{���D�H%f��p$��^���N̡ϵؚ~�X�jTǞ�����r�_�)�.H=�I�]}U����U|zw�-�K���4�����[J�hK��;Er�4EM6󵡣���n��w��fLd�b�hx��-5kwH�Y��+��W��3؉6H�o�$�}�}*m��;Rg�>��x�~���g�UF�A&)Q��xGM'�5hG����p�L�����'H�B����Cu��N��Ñ�>aM��	�[�xp���8�!a�U�7C�;�$��댞8����im�K�ĵ��g*]K�j��H���riT���s�)u��lw���a�Z+�z1�t�K��=��|�	W�~��m���kP�\�'���iF5�w��=��Y�vPl���)cV�b���"��,��q��m���]k�(q~��@�~���(���`�`�T;-���M�u���J�ϭ�l�YD��ƫ��d��EL�r��R�5ՃT�f�-���=��º9����[���̡�м��tC��Dª#	hK�� _;EZ��P&F"CTeK�T��˖1��Ao�B��*��	*�T��jV�Bu��\�y[N�2��4�D��L���0p��[�J�/R7C��TT�E6�^��Vs�8ly�5Fp�;�۟{���i���)[xr��R��>rax���9p�t�r
)��\1���\�{���,����x�]�rv�S��@�dF�6�e���Js�g����W������v<u�������n�&�H,����O�.2�F�[�e���f����3d�����Ij�NPu�q�0��yT6`S������a`��ФBv50L�hy���%j8h����aG����!��O,�D	��xm�A��� �J%����D�oW�r�lf��o8h�*�o����e'<���g�|��?#7�K�%�<�:~377�N�R����`�|ю,���a�^a��\fnD���+-#�.3y<�2>�R�tBckOj=w�[��T��3�o
f��3�r�_p���ώ��ԥ\���IL��c����M���*+�E���%�Z�B�gF;1�ǒr���J'���
�������n0(J"��צ�
W��K_����[����~X҇����h`v��p�}�����VW���#�Ak�����4���=�4��d�GN��G`G.mr��~�:Ì�@,S�� �,����[���JS�@���/#��U
˗���~�m`ě1Ћ��R��
b<}�6����B
�	�Sv9]QW̦�4��a9�z�9��̲��0�qw+¦V��趞؁���D��V�\N��,�Z+[Cb"]���hVa���s��L�a:U�7i�\���O�+��O���b2gC{B�r1�ʋC򫢡si̞"͈x�]�j&S&Lؚٸ3�S����F�6����`�����&k��]���Οa=F� �q<�]��^�Ԕ�rT>03��Nɻ��*pF7��v����S�	K�JU�u�"���E�,���'{9�1�uS�v���.3�ZB� ��V,]���>�Z\!7�|�9+��s�%j1_���S��n�P'u���F�EH(���FV09ʛ���3�1�dR�:b<�K��?K��A��'�+|#�%9T�!`�̍ڒnݯ��У>�JZW����v�S�0P'��������mQ���&��'�T*�n�݈6OL��PQ�,��p4�m� � �I�*���'\�P__+��iV�B�&r����g�.������+�:0������աA����G���I͢
�6�����6�'��W�L>���9��k���@�A�K%��}�1�ç	����a%������?�����<4:����:�����_�r0D�Ι[x�0G׸N�<)ԝ�fK� ��r&�>'B�G9n��Q�����Nh^	Ea,�m��L%�g���zw�P��z�)4zczri�F�9��w�Is+�V*LJ<5�����s��Z��[4:t��D6�>��W�x���ˆ�J�i�wW�Ә�,��i*�>�m)�a��Э
�n
$l��MX0^�,���Pm����ǿb�(nO�Z|N��� �Hg�_��R��F�\#��I�v&��
�b�h} sbPy*�<Q������{YJ'�Fյ9�(�YMYc �����W\4�X'��#����%���Hᩊ�!od���,����D@���Tz�mN�})T`���K~���N|#{%��������%¨�d�tŭ�K��+I\f�L�w�}0��c�R��1�K6`[�h�w�]�_PJb온ihu�b���wb�l釉���SZz���{�� $ħ��}���.��<�,Y���#R��l冴*�B-����-j�@��K��қ��jl��Ã��[Gk���g�Hc�7�Q5_�T��«�
!�[0���3�A�|��ҝ��Ba�H��:�i�{�1�L�Ur��,!G
=�2;�)��>����Yk%7Tt����ar�36��%]��<���+�Cfj5�9�,Z"�9^���A��sw�^���Y�G�V�m����}kf��(᷋���ܬ9Lu�ʬ|��'��瑉��(�Zp���ۨe3BK�r�?��L#W��" ��J�v�
"�6�u��TX������^G��w��U!(
;���baI�`��\U���`h��ɔC^x���rp���汮���o�֋��u[�Ǝ���7���Iz9L�T_�&��Gn�$JO4��@�/�:��߉�O_���C__,dy�]X�W�\�tl��ѹ�~��6Y�64c$IU�`����MV	B����`D��IOHW��(1�s#'C�|���c����@�Nڰ��5�l�/^�3��.���Q������w�{c���G���FT�tl�vg��ֆ�J/�ʄ(5���B�Ջc#޷��M�V�3�!?�%��̂V��V��A��V��J��b`\��|s(?���
�8�'ծ�⊺Uu�sXKw����z�p�y�r�Q��dVJz��ٱGt���Di��>r;Y�Id4���+�V�\e�|��+M��5q��M�� w���Wn>�~��,w�Z=YF�'��QR�2�����W�T@���G�XGp1���Sh��d�	d�˫��ܦG 8���fa��k�{q����k�t��udx[
&)ۧV��B�����?W�_�:.x��<`'�s7�\��@Xކ9���le����%�mE�j�@D�m��!��[���W^DcBm[�~�����4�"<e�2�Gk�t��,#�2ʬ��q��<���Ke��F���n��p�D��N�K�!�rk�2�.A�
�l~���`��<��BL��j{��"�B��w��.-j�S��Q���?W�qz��y�?���EĤ�ބ(=�ݒ����HReu�~V�@��]��t�Rl�*�����2ٚ<E³%�XpAU�1] �k��\y���~��P��ώ��y��P���c���E& ԝ��$����j�z�V1���[�g���qF}��3�-�#B{��D���0W��z�T��Ʀ�h���1�i����+�W}:w���~�!,=�*�����}��hky����;��M}��}��~mC�qx�E�����~Ԣ�2,9��<��t`�iid��[����3�}��q!�+�藛ɬ@ȠVm���p)T< �q�橗���n/�U��(س�����C���ɜ9�E�|HJ��W޻趔9�Xj䐚��VE���n�0�f�T;S�6mi8cѲb�5C_f|�u���}��U�w�������c)�.�)�=B�P-����-��o� bo��:�X�Cyw�����?/[�#vrA�!�k�w2��״�wxF蓯���&�e������.wr/m�vs���x��-E=Sd��V
�����1��^�`����V�\o�F'�N;Ǐ�6[~K���6r��s�$�Ae������I���0��C�ؕ[�ڃ[��ǡ� ���MH�0�����	�DC6�3M�ӥ��Ihu��O�����!P��m���[&�/�Z�85F������lY�ct?z.�����w���M,覆
������M8X�֪/\t�	x�r�v��!�����MӸ"_ ��h�P
�e4a�JxX��A-gf��^[�X��r��v����I�mH�8W��DU������BȈ��K�i#��ѷČϢ�W��γ=���R�!&�Y���[62LxkT�����3 |���{D�CYJ
ޫd��4P��3�Ybw�+:���N"�dm��ʂEq��+R�2ʪo5�DW�b�fׁ�̾�������/7�]�fG
�(�(�:��'�m�j������@�n�E��P�9#ؒΊ�*VC�1P�~��q�k�d�cs#�j!+��*��[�w4��z�#1��u?�|�_x�*7��Y1�i95�:�<��@���Ax ��!￿+�сy���ц-�l���>zcs�'A��N�+.��v�xV?v�A�����w�)}��؉��U��h�濏QΒ�=(YA[9hNMPc5t�Q'�+4����*�J��Y�\[���ŌI�d�Z1�hY>����!�$��ݜ���$��#\�G�tU���F��FE��(�ǯ.}����n�܀=�$�K�HH��TM�����r����+��p}���X�%�_SF���%��*�3AK��M�v��&��R��T�/H��V��V��y�/=rL����k�u�����=[�Cy8�
���1)� �*�8������T�+����w<���ə���(�/P�L�º�<RV?�ǚʜ�(��f��d��+2"K��iv|���98�U�H�_��*��ĵJ[=a�:��1��]��U����.A�* �+[��\�p�~c4Q�a�� �O�Ty$W����Ҋ�ܐ)�Bm���&%	 ���W
Tm�׬U�1ߊc�v4hz�oq���	]��C!�eQgsSAo{b���k��3��"����v[���eq�����ɸ�cu�Q����Iǁ���Bp�>K@"������h66!$�%e5�txm|Q)a�;kon���H�� c��s�������o��c	��n�\ۡ��#�YH�A�Klۍ��/ �7�H7����y�/w�\�����F?V�)H�w���KTLF�R:־��>5D�H�}�'r�澶 ��i��(�Z���~fH�8�Cc��0m��J-�:�?��?+��.����� �b;��ZdvkP V�$�f52�a�3,Q�~��9�SX�5Q�Q2�rؖ��n9v|a�c_I��аҀ�E��HH�ya����h�|��Z�n���a�P�)��1��y3P��K��<Kf�䚀���W�\��z,��A<��JW�n�"{g6��©M�r�F� ��yF÷w����~ݙ7��.*��I��� �o�YR3��֚�ZF"�"��@|�E�m��$�α��%)�_ָ�mH�@��������"��$ft�	՜!&����b��>�џ���*�%�}{�`�3:�0\G�:�������S\~�S�
�*O�=u�F��K���Ȇ���wgO�#ߙ�sг��+�pS������ݵ�cOۍ{���Pc9������M[9������6#�(>�Y�ý���֌����e�>?u�A{+�[��~G�3ό�6�2aCf��B2��d}q�8��S@f���7���B	Mt��U��8!lx���;Ɖ�&�ƈ���a�v�)��f�-g�Ţ(<m���L��\o󎒫._�tʽ���*o��K՗��؃�U���Є��D z��uF�A��]X�������G�Y��GM�m߲���)!��ϩPdқN|����Zzf����z���ޓ6Q�אs��4+�v6�蓠3�b�S@���?fuި"�!����>ڋ�XBi=VU���Q3ߵ;Y��3����h��[��rW��ړ�qIX�/{N�M	^��'�Q��|����A�m̕Z(�1]�����9ǿ�L�-�zU'{y�OS�}7��jEw;Z�h:�[ ����2N�>����sp45H��)����Ɖ�d��s�9^U]\`k�����l������(g���2�W݌B��u�ʗTa��2�6��-�#޳ss�����!��~����?<t�A""�M[���郮x��+��5�{��nHp�1�|
���V���FoQ��o�H�[���RԞt2�D�����},�}�&��3�V�o���J3~W�\�@;�g�Ò#D�K�GR�;��o��}ې�lK�|��<��s�{>}��pH�6jC�0J�mqZZN|�X	�[�|��W+�z��m�`ӊ�SU삮]���a�?���xlK�l�<?}.��V��T��ܷO"ԥz	�����sk@/&�GН�$JЎp��o�;]F&��O��P�a���q�I����G��^��
�y�_,H�U�� |n^��'����W�(gA��7ę(�ĝk2]No�@ӵ�^1
uOڧ����x����	�טA������dA?))|�!��i�p�m����@$��fѽ.�q�	�H��(�u��/�;YC̱�Z�Je�qU\ ��"�D�����~�;)��{SZ1�&�ޟ�W/󠍖��h��E�7�	�p����"�W(��yة�d�ٖ�"j�7]�l��*~;)�KxHr*��'�jD�dJo�q���r��#���ɼ��t��ݪ��?(n�qi˜Sb?�s֩BsB�$eχ�������k�7N���F�kS�0����2>5�F�w�#�����w�t�L���:5��i�Z]q���`�ydަ]�qk?"ԍ�~,1/��6z ��>*y=����|ߡ�癵Ҋc�P!��n\�eߺ*b�A�/�1%��&+}K��J� Q���L�hU/0E��Z�V�f�g�2�3� ŷ�IZ�}�MR��bY�F�;�Mf���p�y]��br�y����~:��ZH(�mxr��Z��#�$O � ��6� V"�E���[G&iz+�iˣA[����z��ΏTo�Y0�L�2ɫU8��d���z_�`�7��'��#��R_���%����gĐ?�.�I*E�|����)�`��U�5�v�	�5�%��!q�R
p�83�B�%�TT+�����Rd���N0׶�����@ɽ4lӲN�9ќ��A�ȶ�|���SΔ�2�a��?8gӿ����!���_$25e�7��uSH<�S��(�I�#��C���c�$��Di���i#�te����_��k"Ӌ������^������w�����c���������5k��׵���%�� E
��7f��*W7���\�j*���� � �ꩢ	V�s��Xƶ��7�� }I
�2���)���E4dAN�=|j�?��m�i2$,I+^`;���9�V��y8�T��-�$�$_9r�@�O��۳T�G�E��v؜q����=5���_p��}&J&�z���&�5�-���/��嬪'bV`��gi�`�͉f�l�f�c���A�=������l\�K�
?^�X����Æ����X��N�����P��0�6W3(�w
+�����CNW�u�Op�f���,�^

[&�&'υ%PT��*�Li��^x�Ne\��
N<V�'�|_�x ����dHFC�&R���Y�>k��d@�4�T�3�"'��d7�x'<��Oǋ�y^��A�wPi�Čs�����sw�<���0��X86�Q��Mn]gW���s�yD_��`�]����\΋�7.a�F'ͫ�J�H�"��!�/���[?��i�\���t�'n����˅��I�W��B�	-���O'�/��0��L��p�b��-wZ�*�xv��l�S���"n$5����Z}���º̫��l<#�)�+V�m*ٕ��^J&�M䤠;u�ð�q�w%R �pS!I=$4�wd~W�<����[h��%Uԋd���:��<��3�O2�����u�-�ٌC홷 *��#9b�.����"6X�S~*�%��vB��� <�j�t� ��)�+Gv]�cF?�.�;h�/�퇃�c=߁���`e�:�@�lHx_���9��:5� l��ĖA2G�:D�h���f�p����2����Ҭ��5ٲ�u��H2�{�s<�j��cF��ȣ[:-g����4���R
P�^zU�k�[s�C�r.��T1b<=@��2$�v���n!�e(�u[�1���v����B�m����.���DǛ4���z~�3���T�.^�Tj��	|��M�I��S0���nؿ���p���*���aA��~C�[l�L&k*�%NF��L�����:=	�����Rcr0���|�rWD�	����IoI�<i�,Ğ��ؖ���#��Υz��w���z�u��I��@�ʶM���VO�xD���K�GogLj�M;K�-��B������2ɖP��6{��Nî�a�͐���q?V`3Ȝ1�����ʧ��\d7��z��P���C�Ύ��&�_�a�Y�o��hDS7A7���U<�� 9�EK�ӠÎ2�	�(�HG	Sמ� Ng�rmnS#���C�j��x�:\�T�L���������?٣ܘ�Y=V:����)T?����
\߄��w)N���JԌ���ܰ����U�D��(%qS�!4}A�Ĕ�bp�T13�R:�^ЯV�b�F����/�utg�$
4����(���\�_�܇��z��ܣ0����%����?��.�Cw3	�4��`A +ܚ�:r�Sg7��hgKr���PQ14!��ֲ3��������6`�[�;�F*C��7-'���M�P7���A�f^yT���(�x���Q'%�aC���z�]�NU��s���M!�7nx�=9�A�˟X�#�8\{���l�e�4�.$�j��ݏ���5� ���[��ecS�S��!&Y#5�V�n>E�:o�&�XlEa���@
�sI�4=M�B��!�<ZOر@[��gf���I���OIg�m���2����},�M�-��7�ւb�������~/"�˛<I#���E�j�5ÿ�M��6�a8��	1�7�2�BP\��D�M�g⁥ ����D��u���`���|ļ{�P���Os�tp���8u;bˤB�Vyn�F�I����K�q�iu* T��7mD����Q[�ݞ
�۞!ׁI�/@�V�<��:I[K��<��Q}�?���9� {d-����J���8��{ �����a_B�ۼ��}�2PU��:S��Z���g�h���Ů2����-�n��ܹ�Á���SK�} "�*��lm
�G޷���%?�2���"��g�C�S�L�Lnмh�W��GDqkn<�x[ON�{��Z�|�J-�:dBL��kzĬ_��J�5Ѧ�z=K���5z����4��Q���w6�d}��o�d�(�O>|ne��]E��~�.B�Bq˳e��G��U��;��WϽ��Ig��Ir����f�zm|������\�lhi��$+^2E|a�	M������y3��Ԛ���kn�K��x�\ql���`,��ma.b�%aW��C���ۻOՙ�L�e0�N���!��cF��b����kGVd��6TZw�n��t�J�}A�-�Q+~~�t�ƥA����rD�,��=ƾ�9l˲�ַ�>�-�/����U�����-s�6.�^Jl$�@��P�W^^���!�����~���|��ƈ��Y�O"^YW��:��'��u? z�UB4s�У��x�>:p=P
��L�٪{U%��Oh� �u�|P��>�D5	��(Q��]�:�`��z϶"'�%b	y夎x��N�$o����O����7�\�홦K�O^���esU��hU}٭���ۏa�J,��v?�HsI@�|��ҝ_�ɼ��|�xڭU2,H!�=Xi�>����OA\�0�d�8��Ohe��]�˾�[��j���]>��k��ϙ�9QFH�V˕M^7������]@��
�^�F  ��k�]�� ��?] ��-S�L�����V��6��=$]"vn�~áI�j�@�ߢ�WV��No��`3�QaI�Lަͩ�N��BbJ�\n������y����s\ﺮ^{O���K�ԑ�s��`Nz�w|=�t�}U9�����4�z�X�$��@R�d��p���F�W'�Q@9�m���y.O�c�ɣ?Kq]8�(cZ%.���3�S"����[N�Z��cfV2�t������
`�Vg�t˟����Z�{(���cՐ^vؠ�ܒ���r]��Q]@�Ӆ`3J��$�{�SL�^�W��p����Ӿ{�ig��O5�a���+ϻ�ϲ8V�)�تXR<�PBQ�`�.ll�����#�{xk_%a��:�'�
P�Գ�<>`�R�u��5���v�?J�_%E TfTX_�uB�,��]�
o�6�q^���w�١�О�^�54\P�5��Ir�$��7��!!Ѣ�͢LG}��A���)h�Ͷ��&�uNB)s0��	*̩����S4a:�����j�%���'�z�2�\핉�]���B&/c��.�݋�w��)� *�@�R��8u��%�HM�UE�dJM�jq��tF�E����C*�*`%LX�й�^1�E���Ub���qgȡ����~��+���z� }bR[>����E>7�`�@� V\��Ъ[34�$�M�4JF!�C�������+ቌ�MD,�U�_a-��������{_�X��]>+���~{��No�7�rr��z��U`��2��6��l�6h��M�tn��Qe�Kt�����	�4����6ۿ�x�6%�5�t���༌��~2��?)ƒoxEvIa���iqYԬq�ſ
��������S�	UL�c�V[G~dX�3Q=�1i{�<����4^��G:6
D�.嵊�ܝO�l�"g�7��ݘ�+2��p�c���]�|�8D9=F}��y���n�e��}�L�#5;���
��O@1U���B�,ҒI�[f;G�8[J�<�h�M����c���F�7�����{��Cyz�\)p�,v���?��SGX�Ֆ#3��ָ������Q�=�BֆQ�4� Y|�d=$p���0���^�
�d��h�$YY�Gĕ�Nk�Z��ĵ?�x(����Z*}��EON�?/�[J�za�r����&���?t�K[w�|^s��PY�b�-�������Tנ���?�Δ��f�ѐ9�X��7��Ef�X�"�%�Vb�~C/�?�2Ln��w�M�T�0�;C2 iyo���O��%6������^�Y���-�T����]}�"��lA)�$i7ҌD��	0p��K��7X���`�;Wi�1��-�"� �"�k�7#���k��K'v�QA���~��L��x8bs�+XP���$� �t��%/��c�{�dk�M��j�C�$��:l����� ���a^��a_�����݊��vC�z�v�����Ԕ#��Q(���ۓ��h�ƖŦ8}�O?��)j9���*?j��}y�/�_� wg@1KA�E0bR^�T\	QU-JAd�pE��φ�@���as��8�E�c}@��W
��p���f�G����do��S�?�3?�b�2�ګE}y��1V�]R�o��N(|���;�>m*�F�1�{MYt삾)QV��FRx>�x�'tKm�p�%{���>�<�K��h�~�|�07���7)��(��z�^�yq�s���d3�����d(}	j��Z�X�^�����7))i%�Uc橮�}}?	Qڶ��#F<�������s�����N6Mj�W�	=����E�#���5d�J&�kN�?c��Lf�DR�Iz�{s�j��Ƹ��+�3ױ��g�^Ԥ��rql��˜��#=ԃM�h�e�0&B�"�hz��ٷ.}��t���J�H9#l#;��ҀZF�ˬ�O��֪��3�Q��
ָeձ�y�
��z�5J�~��jзH�:� ��h��m�K����c�i���҅[X���v��y��Q_l�-�kI:y<�6�rx]6��H���j�����!��@�2��:r�T��ՇqAJa($θ�JyE\�yAQ�M�^�~�/��X7m�)� 
��ĵ���g�'�#��O^?��Tc�q`p)�����O?�qΊ�pP���X��cg����0�L����B�O�4�6�. V���_��Ő;����&�j���a�X��wv`�Cq+��#�O!3WO�}	��_j=�?�*�ո��oB����K�qnpɏ�0�"n��⨭�i��fq|��G�L�c�_��/��J�7^&4J�$8���˾��s��sUw�G(=�]�5��'��h8	ɋ��?%*ee���d!�:��
�9�;AԀs�/�XlLgǋs�ȃ��R��ES����G���Rӊ@�J
��~���,���k*�0�/���ܯ��Z_d�V2��zEj���?�1\v%����f�]ۧu��M��}����qH(���l�&����	���1���e[�$cë���왫&j�IwLNRр��%��ݩ98�\Az�#�yy��k���;[&� /��/���9V��E��zG߳�5C�P����8���A�Y�����WU�x����!�u^����Ѧ�X;��CՍ�]�e����ʞ�'&�:�+W�c�aNWm��[�:����Z�_�3Y��� �w�\Cp�����Ԙ�6X�t<{��Y[��ˑ���ӻ�r脞.1s�P�L	l.\H�zbJ�o�(��S7���
�Cw�T{�a�T;y�:0��7��4�(= �T���tRT �M�~k}9�[������Bٜ�U�ȋ~m'V�8��hG�=�M�-֥��9�	��e�>��%�Ja, ����R��(~����QNs�]�I����E~t'�g����8��q�zBт݁!&򹥭��>�N��`���*���!%4�EE@=�O�}V�qܕ��ʸ�d�+Z��$<��ܔ���3ѠRN��1BH�v1��/�)�G��рg�B'b�Xk;�����}hr�~,���� pJ����*m.|"՜ �$��7ɷ8e74���p������&���}��'�mf_��h�ߨ�Z&6Y���� @s�>�7�p[ӒQ�R���yz�<�	/ska����@�zFZ�?�}3s�*Ł,&�(lM�W!��d�\N��� W��SZ������Ii�V��N����NNr.�����}�pN�)�7-�I���lR�嚥�	D�up��ؐ���ӥ �|9�л�%�����Q��LE*�jq�7��!�j�?��}�+��cs
p��N��o�dA}�d���_��q�g5�V >���+�X�N�z:_�e���V波�����P�|[��`ZW���V�<=�]"*��� g�v�3	�C\�j� ��'�E�?���∗	���'N|��_D�5�����5�e�#%e*0��mM�0J"gy�:Uƚ�j�ƿ������L��Q�zˀN�N+��2��;,�S�k<ӿ�w��hnD��������A�@6ƴ�[����s���
d�*oZ~U8���N���E�W15p��O��	�I�ƃr�
os��W��~g@#��ۻ��xgL�q��#���{�v�z��:IE�t� ��Q���7o3qY����%��O!&aR�"��p�DG��!Mrx���g�R�+���*�f������T?�]c�j�@���.ݷg`秏}��o� >�6�TEq��� ���Y=�!:`yĳp�9v��=I�xBP�~B�<E.&�S���>�@�<�Ĵx�gs�8�R�4e���	��B#�[f+���r��)c�z�J����s1?�\��m� `�����+XL���^�1��*y����{<�ו�R B>I�%�/��8���1�o�%�&Z�y6��{I��,8�g��}�h� +�1o[ʴ� �,,T�;ͅ��Vty~%Tuɽfw+�,R�޸#�]�L�I�N"_�'�����ި�D3���_I�����F6�ŹV���Z(Ά�b�bau�vB�	�JD�!��X�*��~(��!*����Wa�lQ�v7GY�{A�^�բC�1P�`���A�L��Uxy��O�^�O�e��!��,���P� ����$���F�؈�j�0E��������a�ۻ+r�&vDmI�9�?dԇ�
-v>QU&��A��} ��e�jZ��V����}�w���8�9ǡK�����s����X�s�e���d�F�� �+����]m� �܌��cې��؎L9:�=�����t�gR ��}�Z�}�t�$�EMO���3�X��yQ.��$ib��Yv�L3�{�Ƹ�O��w�=����:���c+�GY1@�,C����]V\PjE�ҷ
�)l*D����;g�m�'��}�څ?Q3[X4�Y mE�E��R����$L$c�"c\���@|��+ԫ؏�z=��CWH�7� b��C5��m�D�ӭպz��~��9��P�1��-�����;�9d��ofQ����rOv�z���X�F�ggW�BpX?���ә^��5�w��������!�r��s?���5
c�������-��= "羺�n��2����-����e�
z�o���ȐQv���M0��4y ��3Dq�Ϥ�{�'T=�z�b8��`D����~��L�Jk�#l����u�]�T���e'�ú���$b���:d�� �`W����𖽽���=���=��I�1���Z�@�]���wA����V����Tu�s��i�}k���j������aG�|)���K�S��? Ϙ�5R�
|�D�#��Z	����@1�7s��TMK���7j\�R�?L�i�g^���HA��&�I;�ȗ�b�(iЖ��C�Ş�ǋDu��R�	y�%��޸��6@��[�;�(�_g��O�,;�#@�� Y�/l�ތ�5:n# ��I���އԢ�D`��}	�{	�'�� �������+�9�s;�2t�M\ޔ��JA��!4��Ju<ݨ��墌y�{�6���������e!�U䑞L��Ma�Cg� �G� [l��)�ԭJ�k�Z��z�f��tS�<�!L��̙�M>��������-�#)/�ݏz\E9���7�+�-S51�����a���E qY륿S�
�c����pQtTD�d�{�Q�]�ߕ��a�E�(��S㋰{0a�so�
PX$���w���唧h��E�s�_u���?k�npfTWpl��P�;�z�(����7G�{�?�6��|�l��R<�q���Y����&�>�F?_F�; � }Z�T,��#���tG�GU&�t���?��j��)����TK���X�J�eI1�(�맱r��C���4���Lp��p4����L/�7�ç��>h�8?}�)�9�'.�\��S&�NGRL~`�_�햂Q�jP^��+������܇��]���뫐E��[NqU��e4Fc�2�x�k�?C�׺a�b�k|�##����"��-�YU3x�l�r��Qg?��}�$2�p�eP�d�"[h�*�m|z�?�)���P���F�6��2���!=��{Dj*�P�ty�=�Cu�"��:��GaXM�d�jJ���<��w���la�41o��w���&ڎ�TV�@!����?,�����.��,ڧKqѻ%e.��w��C��v�D2yQ�`?�;��1��:�-��H�8���B��Cdq���$�3岟��O%�v_����)^�9�ּŻ�h&ܖ���0��R��$��UW)��=�h���2@�5�d����c��
�X�|�i'~z0��,l�������0i�Y�:B��#�b82
��j�3���\J�.�C�XiK1���5���Q���v�oDu�A���s��Shbl��cr�I�ht�j��\{41���NmWV�Vd�^�Y�NȊ�.1�m��$���v�F��Zi%{f�t�[Ŭ�y�yL�Nq?�����ć���у�}d�o}�u��Mv��54a�#|����-�7�7Q��`�no��9�r��������\��Dp(��#x8�ɰ�Hw��Sw�Mt7�j0;$�»���գ"���������Y�6DJ�ym�@;����	-�~�N��F������S�zSg�(��ѿ)��:��PfrD�}�[��7�.l�U~L0vq����-΋����Ċ6��qvn�"��g9l�#.���U��Ȳ���:���h�R��P�����$[,A��O��W�2��賨�AD�Mɧ���<5��; �)��8j��Q���?����n�J#�d���`�1q�w���,1\��K����f%�k���SJ�Ug��Ԟ���L+�v{z�P2<��c0��i����1��&byݬ[ќ_��;�9�i���҂�˛G���0�JQCf��\G�Է������4�u{Kp�f2d���|�'`�����@�ɨ�u%���H�:���� ��HA�n=5��O���`w�M(p ;*�A�{xQa��z���"�J����f�H�U��=�	�m����d[ːp�Q��h��.�G�)>)�s� sMK����ZW�	��!��(I�ZI��,�E�I��L�"{?�������0����� ��b� ��&�ǡ��^ı���*��/�:?��}氅[Y`䉴i��璘��]�$�[�(�Ԑ�y��I��	��x�5�04�}fP0�/��V	�-�Y>XU���H�'�\���>"��Ć�vr��a��wO#��e�R5��@cݵ�`Uʫ�o�<D�%d��ei��Ѓ��C J?� ��p>��P+�̃�"���,�i�O1�������0�Ļ�a�>,:6f=$L��2»=6/����!n�t�����"��|񷯻��H�F�q�^�vp�����h컀�ء��O*����O =G|pj�ɯ(���d�a>N��0^Yх�Ö�C�B��� �A��߇a'JS�[ rಥ��x�V���X��&3�z
��O	<� K El��d��tu�+��/>*y�i����b�>A��?tΫA�J�	���~ ;�X�
5���/ �ڭO���TD��r�N�����*�u��r���Ԡ�~ߌ� t�$�˓	�o�9�V�Ȅ�:�bm�J�yoTO� ��J��v���梨Ucǅ>������=�"[��A;�G~�n��q�>U[{\��v��-�5�:d���)�J3!<'9��[�;$��,t�0�I,Ph	��L�+����m.	�9�8��TB����:��́P��NZ��g?���G��Q��UpЎ�̧^E
�)�:��~
转�]YD!ti�''&a<�4g��x\GC�ۆ�}�iJ�Ȍ��A�F~��}���c�mV��/�Sa�D�����D�]����m1��H��<�Y��n����M��z�ɓ����*+vC����`)AL
H	� \��WB:f[	{��T��� `Ea���1O�}�
~k48��(#�:i8���BE�,|��rD��T�X��
�e��z{�꾆�������7�x���nk�����=X�!����%'0]�)�S=�\6�'���ZT9D��!��X�*/m
������רT�dbm@=������t�D�h� �P�*r���R
��-��G��j�ͺ!��9�)X(i�)P(^�_�pN���*��l�G�s��E_���a�ph����I�&�:dE����O��iB�l>·�,�:�[���X�m�f�襲W�@;���=�%��ͣ���ݣ��q>�C�]G��aĚ�!Y2;�	TH��L��/�
S6|�ԝP�S˳Z��4�џ�Ƕ�;��?@F7��v���p0��M�;@*�8��h��ہ �;�e�PJA��E2o�1� z��ە�8�Б�W^����M6�e��/��f�ҨJ�C�,o�l��Q�S�l����Jf��6G�
4�.;��Y�K�S�MqwOx����6��ʮ��So1W�(5-�(�ߩ���P��5��@~}�����h�������Ei��/A$w���rp�r��&m&�r{�20rxo� F�!�Aj�B�~ٕ��|#N���vKee�-w�d, gy��o�t�9�^kڪ=��aO>�(�g�DH�2�3 :���m�dmp�[뺧�����8? ;o��\MT�x�>~�Qc�t��jUN�O�'2[�Ú�>"3�y	Y��%�ns����S���5�˘}��C O�x<ϰ7�$����+���.R��KC�M���T��F������lY\Xϥ��G�^�G�ncH\}�����&Z�-�l��A�/vj�"��3%Or�l��`��]�ʎ��7+�w�bFc'j+2�[�;.V���j&6����+MSS��I��d��L���g�1�8�Yk��e���R�d������α����4�u�ǽ�A[���V;2��0<:X����ܭ��	�X�����q7�����@	U�rVO�%Oj�p����OC��l*3{�I�7��S /�.�n�wj.�x�q|�Dx-r0��kxz�2\���q?�A�T�W��L���-�9��덷�:�7�θ�*Uk�V^ Ҫ�ps<�-��K�/j�J�"��`P�;��֫6"4'jSL3�=R�U&לY�7���I�2���̉"-C=�RL?7�4�ݥ�Fi�F[�)Sޞ��;���05r(���!0��}���z}�4�`3�|z��4������
Ak�T��w+�ya�C�K,�s���K[oA�ɮ�����f[�U�rW���(K��6��Q�ě��_$��z���Znȹa�j��:�1��A�J���_c�U�:.\��՘dv0��0==t���ʤ�[Z��0؅`�d�DY��G�^�5�Jl� �X��7��j�GJ<n�wo��(S�i(�wm���^��,�~1���L\���H19JAĪ�4��V�sF�h�p� m�_¿��c�,�������m�Kk��[7���(HHA�+���ԑy����7�sf�L͗(�k�5��e���T����:xc'Px��Z80-�������`z?;�$�[7l+`�Bm����!�GU�S��ZN2	y�T� �\�ƁPў�:�w���7
	�&���WEɧ��Nm�RN"�C��ڼ*��gYs���	&�:R�M����e��S�N�!5�qӲ|������<M}qh>�3<r���V?���imP�X�q�F�ڱ���]k���`(/�3�j	AM��-$��f`dM���$$�L<j�����?Y;��8�Ŏu	�V#�U ax�J%����+*��'��K�d���G�b�RƖ.#u��/(�S����f��Ի��qu���i�O���js�,�"Qpc�)��kQH� ^Yg�Ӑ���)Q�Q�5���|+����?���i]gۈV◒�.���E�,�L�ָ�7��Խ�pK��ڨ��UY��9�9Oa�'���f�o��a�k�ٶ ��s�hQSNv�J%��iq))�gL$�rWP\���3J�6!�� 0��F�]��<ovT�����덲�B�moL������T����]��r��l(�[R��E�մR���KQ�H����;0�]�������5F������i�2�A�����]uS�]dN�P����o 6׀ oεQA��m�w�c���e�S-c/���nC'u ������+x�B8[�b��i����$j9FO��c3�1�s��;&d��n,�:,��\>���
?�R��=�h#�A�Cq*|�i-e���R��-(�w�)*��3�i��Ah���7�ڦ��[�$�7:Vm���r�%]���Z/�2��ߠ�/O�V�?�Zye�0:a�;��&���Fep0�'�	]Q|(�<M��{���s�!��t�D����J��ʤ��y�
I�x�=��a6oT*�Х�Wb����	Hքi�j/^���`���)z����@�Oh��
�J5(�j����T!G9r��⟬��rS�;ah�4}1��x�3W8(_�y��.<��V��y��oJ�B����z��*� �շ���/�9�����ר�@��7��m���%q�O<m�W-�{3fݭ
�;6B��3C�79\��j���A�h#�0�,bd��5U���w}t��$R(���:_A�2ט?EzД�¶2�v�F��M%�m��f^����#Q�<���� 7	�`^�y��R?K��E|�ύ�--O�\W�7��v��y�W�<5��}x�`���GbJ��1�k��3��~�n�)-�:�@<}�K�_U���ϕg{3�=��/k��@�P�I���ӑ��� ��}���lӢ��� >�� �CwV$Xw����tM�\��yWm�G�̋�6�/��6������2��gmŅ�0�샄�Mt_��ͦG�4�t��0\ٕ��43������r�$�o��e�L�#�0�XI�'����XoOI�a'��l�z��}��sSw�N���y�.�i��Y� �3������P���ߎ�2�%J�S���zA�~O|����ў!�{Bk�s�����:�LW,ש���Q��d!a��b�X�4����<�A9w�]��3��.��wG@�U��8�P ��n~�R���\��Vu@e'�- h��I�J �6���ե~�A�����K2� �� 8��8G��@��x�rP������ۇ����d]�OOD'U&|hp�B���Bx�_�r�3��9~<D��@^���^���O*f!˴��ů��,��P��q�/��?y#7���a�Q�Ņ�g��<��wI��&몏4g�[e]���ڠG�=DȲT!�dI0�+u�� ��眮�RQ���21�G"�/T�.LJ_���{v`���T�vc���n;:=eK����=0CD�� X��O>7*�����9C�X6��0>E�ާ.�
|�i�� �Ȏ��k��t��aב�s��x �^�{��	�]N>0��Q���Z�Ի�Ӻ��r	h�ګQ{\�
V?���9����w�f%��%fHI4���/��zU���R��.��hp-��]�����ӽ�W�6����K�8	�S�� �!�01�����j��$�?�v}k��d$E�4�% 47�j�R�c�zw���[ U!�h�����h����LrE��h2��ylM=b��WI����1���uh`R�熗���&x/l)8���p�o��15P�6�9�"��E��6����<��FFS'�*��A��(RR�|Q,�;LP�k�vx���e��ƌ�$Vc\�E^�"�+���{�J�����f�P�:q�~�[�=N����Ǧiq2�Zm�G[7,����1A�(	�	���yE����C�� ��:��z��'F����Е�������J����H�55|���!o��
mσ���U�7[s������g<��ٚ����5��eDπ���q��%8��%�����ͷ��.�;Àb���Ly�m��#Ir.���w������yVv(�҅ҭ���AI��uuk.p�2��sБ�1
�J�8҇��&��w=���W��[t�TSom>�KL�pOB��^|�^���y3Ad-�mRk�-�!����2�-���H��\d�[ħF�n�����hv5��Ɋ�$ˆ5��T��;�e>o�Py*P��b�'<��0�J7H�-��#B^U�|�L�\w�����}qO��]�����tR�8R���^�fd�
���T廢b`��NH�|���ܜS4r5�|J�بu����0�B����w
v3X�!�n'�[u2��/�-+��tI�`O**�F��	V���} ���a��Ԁ|���x�jˬ���Au�i�����%�Yaf����#J�"�p�G�N$��#����=$T������"�Riƕ> g(��[Ǟ#��'�"�ù���)�dj��@t�&�:�ب�$�4��n���5��nyL��L�x���BpM���@4\�����}�;�$p�o �eD�[4��)�p��)L�-�V�UH��u�My��%J���p����>��{��<�T��Eh�[�u.:�|�B�vF��D�$��+� a�_��;��(+����-�;%����s�t[C�D���2&W��]� ���)p� !����͝����j����ktj�(��`�L��eoDj��sͲ0SMfEdu|8�Tf��G�� �T�(���u�0�LꔶX�=�&u1�;�r�K�X��/OS�,��"O����nL6pY�ט�"Tv��%	�w��À�N*�� '��i��&�W9,h'�1�E��Tk�F�8�c
�^��g��{�3S�v:�B��M4 G)�ߠ6 wf	��	9��n��]�9�L�&d�I��h˳�4N�3e!0��YMw3��Ћ��F�K_�n��$攊�,��zGl���,c��A1b;��߾pbsh��=(^2���Z�]F�q�;�;��Ԛ�	X�w/����)�.�5>pn,dk�>�irS��A��j�@ߜ=�]X��/#���yyEJo �b����o��Lx",u�S1�^��"�s�*W+��Ň�DT��%����`�1�F���2	2��������t�!2R\��eP�O��G鮸��Ä3�H�1�nd䳔%8��m���t��Jf�z	��hp��|c���y�	弢Ç�n�c���5���BT�L[������?���� ��Xia�;��0�@����	�j!��u�U!��5��X׮��]�AΈũV}�p@������{"U����^_�[�נ���I�F�P�)/S�ؘټ-4�;�f�\�T@�uS	�N ^c���^�q���:��u�B+Mb�i��IV�ul��XR#gv����`w���:���Z=�2٭�Ud:�[>�d�Ѹ=��Pv�h0%�<zӓ��W���_�>fI$�Uˇ&�D���¨ j���i-�����lt�
G�F!`H��}������<TX���̐ sf	y��!�Z��ᩇ�B��8
��.���7�t�F�~�(qT�|����P��P&���M̒�^6��iH"#�~a��XĠ+I���g��'.��t<8a9��S
�#���s�MF�N�i���b ��I��&.�n��T��N[��n\κ롐Y,��0-~?z+�Y�9��L�Jg�9�ל;F�8q�3���d��.�)Q��E���N�/�*}�X������w�y��Od�Д�<�a"=�����T�$W�0T;*)΅fG~�M�9c�?ըKi�/���yҙ"\_�m��n����`�J��#�6P�~�E�l{�����%���NN�c����-������	C5c��f��ٻ��5EG�YsVM5J�}6�T� �0AV�3��s��݀�)�Ft��]q��9"5X��2%jDp��L$�|/k6Qe��Ӭ[�����1�b�f*�I����>y/�G���.��<�Y��e��2�q�x��w^Ū3f�0+KFVd�^ed/r3G:P��\n��L|�~�ؔ	��*��Jj,�1�Z�%�r|<{�f�.2���~�)����i&�.�׷�ff1fQI.^$����A�ug��~>�	��i�oN� ~1
X}�!賔ڵ�S�}�E�[����2h����j����{�^�c_,��mtxO]Al�'�/͚c<X��J���@�n�[�M@�䄳ǪӼ�� �>�u&4� �?�3=�	l��My��+���bL=���	5�+l�}8��0!��
��ʛ���R)�2�+��3=�-"�~�%f޲	��������w��ڿ�P��	8�*���t�to�yR/I������eJUͥ䆼�$�} �sUhq�DX���0@��ryӫ�a�T�U�4c�8��qט0��_D����DXQ	���{��W���+�gc�V$M�J�NZ`��gwy�^��W?h���m�)e����VpxOtx�L����#�-��v��� ��q'Q��GO��ڟkW��Y�6�K�k�H���`UÕ��w;���o��ioۈ,6aV�	�E��&�M$���~<{�zr�IZ^Q�ފP��a`N�Y�f�l�B�c���-E�C�h;�Զ4���2��"i)��<ڿ��{6�e�,�R�F&Җ�Z	ذ;��Ɏr�P������Y��"���~̹��7�$�e������y��
�R��R��A�}[����]�Ȭ���r����w,�#�?��7C�A��r�A(i"01֧��Rā�2jb���Ψ� d뉂�њ��QEU�[9a!�/���Fʲ����LL�$�y��71����g�ŝ��+G� �z�O]��$-�@�a����S�z����qx�٧�\ȻʹY�@Qa�Y�������1�K�/���֛�.� ����=V���V ֣�bl8���V�w�k0o�t���Ydyg0�I�ϰ��$��_Orf&Cx �:��1%�� ��>6q��J��N;�y�_J��W���7B�K6�jL�Ꮏ{k�axB��g:k��/_�-�%�bi�q"���`�E-=�O�DW`(��j�A|�ek��w\�n0	�0�N�I����k��e�0_#h@G�h�FF����|
WV,�;�3/�v"���'�S����O/fu1O=�&{�>b�T7�_�b����ϭ#V`�]�f4�e�K��G��@��������Pu! ��L�|&\�����i�}�ޏ��d�W��P�֯*�խ!��f��4p��X�M�=K�$��v���hSo�;����RCl���4�3�H�E��E!�����%uQ���L�T�����FM`��˵��A���XZ��Ѿ�� �t�-�}���fi���Cʅ���ߍ۫���.G�1W�Ҳ:`�ʛ��z����Z%�?��zT`|�&�#x�K����Q�qzO�zD�6���_�wQ*i��v&�'���\K�Ͷ�N�4��j��gc�<q��9�R�[D�nYL�]ț
���z��*t�������f��I��4�׶pmp�\d������� �zW�ѷ���=�dp1_{Kapg��U'e�]r�I8o��C��ܡ�����q�aPR&[��~x#�g���\"5�wLqPB�S\�?�t�ݺ���H2j��d��}X����̳�S�o�yx¼�25�þ����(q�{��$�؅��mϹ����nX��:�5�)���,8����C�]2��1�\�wgŪj�����"[7�r�X.M^���/L�\��yQ5��7!V+�%	.�4{�w�Fs�%����6|Y�V��2ePbO�w����PNKC��sb[l,X�J4�W*�;�2
(���H� 7��ٜ��n�t-2�O[2�Z=��hWYH�rXY�s�%��n���^���|z���%E�����\Jd\���7�=�v�h91cp�����撢�H��)�^�����cK�D����M_OD��-�	�(�,��ņp�[@<A�X ?ݧ�):W�A���>�=�X#	,�v��S��8�t�^͹V�nG�5��u�n����Q�����v,z�  �D}�}I����2���B���+��Z�1�xܑ��N����r4�`�����M�ԳE�E?9g����,���sZ& >
��8%���N�.���8�VG\��&[��S�s(�q���u��S�0�2���ٌ�uv�z���/Q�	<;GC�$�
����'�t�5T��w]U��"���bg���_�w��V�-��|M�Orв:��}��01-��&<\�Ű�"����ne���\�e�ȴ߄���ԫ�Y���;��>8��͜�d��4�v0�Ѭp�/Tm}o#I�1df@��]��u�ز�)榲6���PJb�n�x⣮�UNi$'3%�������\-Q.���2�{L��Z$cU�i
u���d��Ȅ��=��>O�RJ����M+_���H��BB*9��8�(B�c(:7?�H��}GF�]�1�;�!0�*��'�O`��j�����B�6����O~�I�/d�V�^Y�? �6�8��=v`�W:��*dH��=i4O�x�q��8�&V:{�߻0w�鰞�k�������˟�}�R[Ȏ�;��xxO��H�uRBT�+5'��lL9z�"���-}�r��������\���狿`����8��|-3%���v���u
�I���,t=E-����KBf}s�603���r��^��;#A%)��&��g������5��XO]dD��ء˷�F������s�Zn9�`�[3M��.�L����o�W��>��u��-���5s�~�b*�]�������Dħ�)lJ�H� �U7�����#��@�$f�������J�\V��خ�߽���r�������dU�#���بz�)ݵ*صH,��V��P��K��޼�U���񭇣�f��4����EJ X�W���������Q��1k9�� ����\ʡ�X _�p��A���y/l���j�ޣ&���_ht�L
 ��F�&J�츲�k��<ID���E��E���P�d~�^}�����vh�f�lM���Lʵ�Y3^�\���Z�:Y�;{FKlD{��Q�-�O[K���YӨ-F�/��:�J9t�"��άQ�F�G$8�pb�����]���Q�ۻ|Ꭳ��\�b#!�d*�Qe�'��W�~<�@6B�W�Ӕ�MmzK����������Sz~��'{Y09�j�[&=��y~�'��$���1�񦌰`:7�/�Tv���d�[�fA�$9N�?P%�1�&웸��P$Xǎ�02��yݨ�&!�5'w���H����Ǉ�x�Ƹ���Sd%�a!C�O����k�E�{���y�����lz�t6JJ�b��D��g
OkbD���9��mzO�����"EceG�|j�j�S�9S�R�����"�$����E�o�����\u?4�dk`>v�g +:��*�V�yX@'ʱ�:*���C"Z�������s�%�l5?I۹t����cyWG3��S��� Dv9_C~��>Ĥ^8wx�= �X��xh-7' ��:��9җ�	�[����#?m��M�Oqs��Y����xx�ē���s�5��,5�yX��B�j�6♉2��ﱊ��~ 2��1Pw![�?�� (��$�0�e�=�L�lXS5�?(����І�:��N�D��I���f�xp�+^m�Ya����`����ُG�pDSf���B�9Ƙ��*/ԏq҃,'�-Z���Ȕ����6�~��D�P}#P�D�o�7��H/��W��DpD7+���QW&G�M`�����ܩ�H�早AƸ^EA����Q��ă���`��Ȟ.�4��p1���^�+�1r�ò[�re�uL��|{�>�	G#D�aD�&֖��d���/i�4q�)^a�^���̙���`��4�E�� -��L�uq�m���,�*�O��r-�+OE)��#�/�V���P�pøp���b�4[�0�1�Ll����m)8�w����tt`�ԣ
+MY�D�h�Ge�e´1���N%Cզl���<�a���ds� ��1vk��!���:�8o�jٟkzÙ!��_��N�=X��<����-���h*fo8.����'?� )�\�4�����@�ǰ��k������a>�r� 9�:0����M
hg��3�f4�'�M��,彿!q�p��٤��\���C�m��~1n6���5����ԩ�1]S� ���0���H����'��=!���BG3ɾ#
�
ؙf}��<�!� }�(�:ʣ&z|���)��:����ĪǓ���a�!�#>�3=D�-*���8W�C�~� �Z������v��5��c�&WM��?��^��4�(�C��Ľ8�*��s�m$߲r�,��!�Wg,�}Ը���ko��oƌ�ͯ��B�wdfђ*�~��ڔ6uX���.���ۮGXGQ��l��"⢏�c�x�ϡ�]�L�'�-Ʉ��������tV3����O�CCX7T�y5I�Q����]��� �%O�P(��e��͌1|6�^άF�t����/ҢH%���)�vV�Oh���G���\����,*�r�z��9Cw�.��O�1�zzZ�lg)jR�W+���O�H�n�}%&�%��`M�7U�v1L����ˑ�w��;n������;�&r!�,�ZƟ�-�P��ՠh~K�W���(jxg;عR��hp�f^6�s���NnPHAs���c?U���4���ׂ�	TZs�P~)�O	�;���wFr*ǒ�F���(��r+�1H,��np��D�D��*��J���MX*a"�	f?-,N��@�"�l(�]²�J��������x�q���Y	&w�<�k��/�I��r�/�@���B㢵hT��ж��ӣ`Ӑ�/�	H ��`���zǡ �:�*�3�턉������痁����y��)!�L�4$�Dj*�a�d-��$��	>��޺D�|df�b.��g��ҥWR�µ�mW�Bz�<�Q�Ԃ�)�đ��zzq�b���e0~��(���b4R�lQ���N��b���1W"�\+�����3������.�^-x���&�T�0/)�5s�k��^(�Uί�Ź�����b>'y|��Oa�I:8�㏡���jًٗ!�ki@�!#�� ���ƹ��5���<F�ٕt�۔y�g
�ܷ���l3Vw(��hg�͒�f�M<�y�3�ζ��ۛ`�b��j�����gX����˄$|�0� Ox�9�:���eiM�dҲ��<�		@=@^�(s��h��8������Zu��?�����X��O8�q"ҕ^h�Q�(L'�{%�a�5�S4�f���$����I��!\�%Z�+��� G�$�R$�X>����n��)�������'���S����K�n������)u��׾�&�m>BS�V�䡤�Ԇ &jI2�(�X,<� /l&-VV��K�t�nʈ&�R�?X@V��K�I�'�r[�������G����@���پ������D5`��nF���dNm_��AW�rar�+�B$B�O֓~G�"z��9����ߌ������5Z;�Bh��S�L]je���rwb����K6��?��u������i�ؑ(�N�_�K¾�����OD�;px���!����KMAۗ#8(�S��E�$��D�*h�(E�3/�[��Hy�?�}U�s���A,�����*8��=�N� ��h����E����n�ւ�&�-v<T��T� �+kZC���`O�l�I��';���~<�~�Q��G2��eN[r(h�Z����VH���(�,T_klp"�����W�]�8����)��ޏ��N���i��k����To�Q�@�n- 9놭��5�?;���ڔ�`����9?�i@�B;���nƃB&�~x�'F;vf��b&�^�y�������3y�H�Hqz���Zk��gO䵈�{��D�~�5�Ĳ�#;0��e����`���K���_y�t�ń�/�mt>�v�sdH�������7|:2����2[�]{Ĺ;i�Bʦ����*�OR�j�js�ɰW//��"+؅L;0��yf����"|z疔�7m�Y�"�M�{��oWA�q�5'��2x�	k7q� J���E{��ȻNbd|�(a�L�0� {!-uU6����y��S+��LՓc2�J;����<�F��éW�����=9/����_#����;"�B���E��k{v�淍QT��9��)|z7�h}�ɯ��vg'�v��A���+��S
y⮢T�JMt�U���P!Z��T���`�D�>�%��c�͌�D��_�bWM����2��+��zf$�f��W��5S]g����4xW�߽����1ߦgm�����������#H�n����H���&���4z�Ti��l�{�k�;p�*��5`z%�A�ZS�ye��Ξ/��2�ӕ9�8�r%"��SP1^i������L���i��ȳd~+.SZ�0���h)7��o)�2��u�:�X��vj���l����t��^����r��h�+�`�J��<Iy+h�A�x��l�����;����	������&�]E9�ƫOn�E��5�P�� Y��R�,�ʆ��_5p�Juf�g�g���\��^�}��ߊ��3�QYԚ�W������Os=�|~����1�0#]�64v6�"�{�����S.���W�]��hR�u��b��!��"QijPQv�i��5�P_�9+��2C��Mzl  Jս���dM+��$Lb�`J���Z�S�j)��H�;C=8��,ˬ$V��E�������2���ę/���G^�oE	��#m6�1%�ю��]1��Ey�i�HiqX��:t7�!^�X�C������*/�����ȲҾp���Q�斓�f� ��_��v�<Ծ4�Bż��ͱ�%k/�e�w�y�`�`����L�"��ݚ{:�Ţ�IЏ����+s=���I����/Y����W����!v,iM��䓁qm�.���Q�@!�R��_�J 0�w:��<�:w���1O���U�[ ڏ��Lt���x�fF]�)�;V[Z�̳}��q�1����;�K��(�z��O����}ڥ��d�F`7؁��7��&�:8��a�t��pͣ�Y�1���݇߆�ҵݹKd�A�?��+z�t9�vc賛1g�_�Ա6�(ɫ{P<�
���) ��6()p��V��,��q�����	�'�P�Žt��b�iQ���s�b��p'�vo�(���T������%����I�=��یUVV�x9�9��J���W�{ՠ@%��G_�h"e±�^�ƚ���@,HŘk��*<�&�Oo����#��E�i.�������֛��2���H�#jA��*�7Ӓ-�f�K��E䒤|Yl��p ��W�Åw�P��@=�3"T^Z<��FZ�ݠ�F����U{�c�@��>q�u����tA]�^�ibsZ��3�����sw)	���7U7g��>W�[�万�V//x]q��OՒ��E'�\1��I� �A���ʕF8��;vw�2���p�v�g˦��9��¾�����y�>[8�����%�@�V����&�/߰&Um2�V
���R��=������{�y�^c�%�p�R-��6����3fN_x��Sz�d꽆�oi5l�n���p��i��Y�������*݁�ک�v����	*�~�A*�i��2���λn�aC~p|�<H3s�����^!�q?0v"<��PH����2�J R��V�k<a��/�F�'��?�������[	zʞ����W��Nχ�׋����v�"?��&0�?���X�v9�;?�J�:(����x�q���Z�Q�)��g�M�>ӫ oT=�ї.�M�Y���%�[��2��/�&��I��}�Ǐ��W;ڡ:���t�ɳ=l����>�|��ѯ ʴ����	����@��Q�[��w(�f�q3	�!
�������1bY�	�
���j�K�ΤBcQ��\i&����ivݸY�h�*��	LO�-I�b����}!t	~�r���f��R�%�������`Y�/+}��T��L*�-fC<�WV~gq���e�|@!�E"/�u �朣���L�ͱ�v����ӿ4nǫIʤM�;j���v������:�y*���)9��8�J��k憎�M�i�&��vԂ�4冭��ʎ�G�1�^���/���@���1A��}\R��٪ �E���(I�>Zm�Ax��]�~n�����Q��xg������Sd�,gt'��p���هf�)�����I3����d��E4t��aY�v����׳�O�ޔj�V�����y�\Ӛ�B)�cV�SiV5=l4'+S���C��.:>����S�������<�"s�M_�ٝ���b͆i�J5�&zp5����B"���P�A������jx���ɖ���K��D �k�ٱ�E����k�P�b���h�*��R�G
y��jBtd�3��R�'ޱO�k#�N;A����"8�A8)�V���u�PH\e�U�"���K2Pp+�l^i~�8V��9���z������"�w�q�(xݘ�Q�ZB��;�������d7�uK0�P�-��Ϲ�v�5+z�*�@�b��H\L�z�D� ^[I`O���ܖ�[�������z��^�ejF[`üI����o-!�JbV��܆)Ï��q$&�KNKi�X3�٬�C������S+�02���C�� =��L4�v��F�@����IM�[b���ߝ���?��<�[��l�ufa��������ݚ.k���I7��z���Ru@{��,�cD�����GP*t��׆�w����� {����Gܹ?&X����-�Uk���	���%�m�d�^c:QHu����߁H�M8���!�Q�COpo��bf�.�$�0h� .! *)�:����4�d�ѥ�MKF�p}��������Zӂ+<?=ݲ���N���Ꭵ�~��k�F�'�w�:6�a4���/`���.��0�HUu >���3�*��=õdD5��@�Wz�!+��í����f��6���H糗(~5�:�
C@�X"h���d_�8G�n��>��b��D����j6��
poƖxWW����Ǹ�)�i�ɴ�'��+1�x~��Q,�D���d6�r^����@ւ�y?Ps�&{Tm�%�s�BEU��=.�6�";�� �D��r�0��>�~��62����Q0�r3ڋ��>ԥ�����ߚ
����vZFNq|���z�hȜ�5�g�ae�0����|y��ΔMl�6�CE��ۣh��m%��+�)��x���]�~5��n��Fv:����^���!��&�9j-M������1k2Ȼȫ�F/(/G$����%���>�f���A��YV!~*+F�:������J��;��B���C��Z��j:��~�bi1 $!���Dn�u�2�}M,Q�9g���7U�w��S��wFZ�r8�p�]_��Jf�[��jc��!K�I��2ǡ/8M���$��%`�JC&+Ř6�h�WշC5�1���Y����S@vƠu{x���Ǻ�GıS��&��rX�uE0��)�0wD�����c�,�q������M�t��M�c�G~;x�B��#�N'>���l�/�p=.�� ZO���~z��<R�=%~?[�N��,�r�%�ŕ�l|d ���=:OY��!&Z	[���wK�������>�'�Aټ�$���+է��G'�����͝B-U�:��AѨL���:�̫���i��v��=_��"�	�b!��i0�C3�"����EG�?��b̊4�1^�u��o8 kY�׺_�i0��*�S�� �`�\`{����<��mz�v��!/�#p�d1s��\� �O!m��a��/xi۾��o��B��>���0�����MP��奖Rc�=Q���mX��xaj��-�q!7v�?�O����bG�E��y��� P�Un,�f1oK]���:�i�X�V��b����K�+���<fMt�+�9H�?�i�*�P������9�X0%P4�Tcj�6SM�:�M9H�8
�*n��W�!�7C��V��N�x��\��[	r�4I@Ü��n��o��qX���쌣�1���;���n����cIX�2)$�+{l�.�u��\uϰ(�u@sϰ|��*QZ:s?(Ĵ����_1�rb����>��X�}�_��
�\y;�_�)(�X��l��́ŻO�UBs�c0U��R�U���hJ!�s���Hn�t�@>�W���0�ߐf�����\��L�~	�h��X^���<�e�#ٞQ��AEiWV�~��[�<��UP ܄��7z�����Z����܏��,��d�ɸ��H)�ՕT���Գ�{���|��Ҫ=�\]O�e;˖��]P,�5�B9'3�s�<�gTݑ�)�j�i+�+j�k���c5���QЖ�P���o�0�%��d(��󞏨��+��1�<�C����^r�ǌ��vI�lCvއ�ͧw/N'n�ęFȠ ��xoO���5�8��КhR��R ��_��r��o�bZ2[Ҫ�pܘs�f��z�J�	"��!���^!	!���?����9���i�̐��<����\nW�����2�UnJ[<���-N� ���]�Ӭ�m��?z'�?ժ�����ڟ����ig<�l�-`�������}n�6�4�g� �
:1>��4���MCzgx��4@�)��8,h4���I/���z��|vx�7���6ӠL�ST�rh��bk��;�鐣�#`�%�AB���ڻ/jC��Wk^݋����탠f���TPZ�v��J~�w����J�� g`e&�ϘĒ?��ݐ���
��M��ȟ��9��9�v��b)f�&���A�D���qǢA�^N�}�0t6�$@uU�E�(�Φ�f�POW�xlq0�q^�nZ����q`�+~�۰ҟ̓�-���/���C~�5<$Q����ߊ E�:gE�*�]�����Xy�)�mr���؋p^N���O�"���E 8�=ȹ���o�Tn�dV��[�}J��V���Z�Td�7�Mi2��,��mp���Ok5����\kk�'���5-�0��\=��;�x6�y��j��=��L�=�d�]�uN������t���	�4�&z_zv���Id)uS�B�p=�U�ļ�I����7T��m,#IS�@������WV���fۀ�����/D`���<��Y颢�Od�¯�E�1g䀕�c�0�C �Ё��G#�pg(�@�r&G�\��M�̿�ޢoX42��������-�U����V�������-E;�� XC�`������7�C{��se�T!o�<C�dZ-�5����I�U٣U����>�8w2I�J3��8'�o�_˒�4�'bD����I�.ո�s�r��0�s�'̪S]����/���o�ʸ=&ß&�\z�6��Zb�RArc��і7�x�J�� ����d�^�X�3%�Bta��s���D~�ZIm��+֯-QBx�\�b�di�>,E��7���k�M.Rcal�Q�Dݖ�[E��"�A��%�����K�S�����t��Y�~�6ƙ@�k��,f�ڒ�fL�x���(��ڛ��i�HO�����i�1/S�5�q�>��|]���%Ǝ��Gor�dˊko93�5bX�%~R�k�L������]^G�?b����y}�0V�`����yW��I��~2��J&;�}	%d%�2_m��#�3�S	W.� �Η���e�x�ը�f��,^�#� �pV(����`c�B��bp�Ԃ��>酅�c�|l�g�"���}#��H>�$XQ��d���g#����B��	�Q���k��r��E�xA��y
�-���en2o��>C�.��&�p��W'= ��|j%��ܔDz��U#C�2!�x� ?M��ji_����s,چ;��DK�e�t�`��F�b �x��d���t��ݳc�?
'c`��(J�G�b���_����bռj<�z%]�-���lO�x24�%����h�,�|h���Lq=��^�>)Һxt:d]��c�������؊>�����;��'�)���'��{p}�S�څ�j�D,�����;�bI��8��iyJ�e �BelL�_Ь(�C�QP���V��y�{Ј���^��V�#�u�I������I��30	!:��CI�H�HΝ���61� ����!��s���mȂض���}1�T]B GтbD>��i>t�N�V��|�=U���J.���GA]�Cle@i��!���H���N�Xѳ�j��Y����q��#�G�>�Z�汀y�S1����(��[x�v�;�.�6�,����9�;��t��sYv�C�:�q���
\co�@:SS�UG�p��v���e���I�T6�L��/�c!?��W�<4�)�(-�9P�v���-5ip�o��C3���(f+� ���~�(��n�6�X��f�b�^ƨĵb#�/�x�������cp�
�:���Al~任�L��g���ʏ����QW��_"{rc\��V)��؜q��B��У�y����'�%���QP�<�꾔.�F_��r�6t��'���㧟�v�O)�u|�v��hc�&�9�N6�~&Wd�:O�6��q1^vD�؝C��w��mڤ1��F�3����\�m��w�$�t5J76���`r��$u�9oN��bA�j�cK˫�<�f���|'܌Q+۸�����o�����R�&T,�(��p᥻�3��a���<����B��b,���'fW���1D���H�V� O	(ͷY�s�wI	��%�ջ�3��
r��EВ��X�s�<Q�nlk�s��%�^�`����̗�R�������@��r�[8�����S2�8N��a�7�;��Y�	���(˓��(;�7J�ntS��]�/z�Ź<g�O!��oJѧ�-�0���t������idG"�?9���bG��UP0 �Ɯ��㣦�ч�l&�)m�_��b�@�y�_�R��29 e���&�%&QP����X��f�Ls>�M�Mm4��$I���F�ya�"џF��V������Gd�r|���g�3*�h�v�L>��߭2x&����ɶ�a3a���������k��?�{�U��WD��B?�e���sU��_������Zq��McS��	m���+�R����j}g���D0wz��o�\����p�MFS�)}i�U�i�!n��ͽh�A�SL���dN�nBy��#�c��jx��U��x���4�5�0Wq8�@t���Ƙ�,����>�t�$mҝ�q�o0mx�.LB>��.5�r{�?��� ��h���7 ��Q>�g�n�[�NX�)o��L8���=s+-ti+���dLS7��x��;:�`f�:~��2u|](�����	�k���9_l�5��<7}�X`sI\)��T��X��hzw8�= Pk]��
�;���*U��!��q13>�)��AH�S+������zŉ��@���cc�YY�n�
��������oթ��*����2;�Cn�^K�!�Hurk��/��`_�J�<�Rh[#s�x,V�����9�1w��W���u[.����#Z����k�/�~�gHDY*�s���}�&W�P�C����n忙hIn�9��#S�7����~P���U���m�S�AV�b2"����M��1(��%|�	�W�ڒ�Sx�K5q�]�g?�uaH�蕄˙��f����4�o,?y��
u?Etٰ�s�A�Ƞ#����O�K@-.a���`�~�Yr��,��ێ꣘:�CAI����3'R7	���]�y��I`H}���廻����*�w˥M�0�@8������MfʭF�ΊIs4���[v��)fb�0�ep�������`��n艠]N��"�WW�n]�쯣c�ӎ4���[K��\H�B�wJ�Y1c��� ����~���s|E�Ǳh��َ��>qp�	7ܳQ*|��B5�.��B�?�#�Y�.>k��W��r�RWL$�������F�J�Y2s��ӡ��Ӆ���H���>"1��9��$
���Ꞑ��q�8���}f��1y2�''�I��s {��Xb|�0�q�,�[^N�2ug'(fr�qeV��S���<�XKO*h�\��wN�n�-E�������M�x�)���=�Z+��1a�o�Sl%�Z=�5�R�{F����y)�M!V����L�����L}&�Yq��i�\��Rę�zݰ����i�6&i�#�s�	�!j���gCse}3\4�La�V���Dµ��Jb���y7�J`#�(%Z�1��ח�NXnPX�4PN-��9I�(�>��&�&
��� �?�u�������HW�)��
��������T��9Zs��������Nb@T�?ة��\{�A@Gy�<��ld�ʔi}%PR
�t�|J2�b!d� c�p0��5"튄|$sh�Ya�Ս
�Ӎ-�!h���3�&�9122����*7��$;�����c�~ �b���
�����/���\�@�%�{�bO@���SH�j%\��e3jdJ�s�,�	�z�X���V�"b�P�$HkoM��Im�!��N�3����f��!D�ts��V�yݣ:�u�3x�O@�h��	�݃���eOs�W���}��XC���D��Bl3�C7�j
�h	B+�y8��Fc�&�NsqɃ'>���R��֕PV(&��%m�׽���{G�c1�!^|�����ŀM�P4�B�;���Fx�)bQ�Ѿ�����X�g��}�!��V"oϲl�{?|Q|��>�]��JH-Q�I����~,���|���a?�H����o���Oֻ��Z���������q���۪�CA���}(?���>�g�W��>D�=U��KO�NW��Pմ����}��^��m�l��/+'D���ǿF���0�N�,��IԿQDX�.O���a%P���Y�wC0{P��^���Ծj�h��� geX��
����'\�ǭV����r���B�>.����$�u��E���́�E;N�1}������]`�s��3�3G�g~�*?#��6ǁ�2�6v����b����J���}q�B����)�Nw�giϚ>G!�O (8l׵���_ݘ< `�	7���<w�>�wྡྷ�����}�m�^&fߥm��a\z)����CA����2xnp�M��#��l�ң��h��T.�r��"���HɁ}�#B�bl��"<�4>H:+���MKU����'v[Ȉ~2��)�ժ��M��0�H�|��]�,�}�{�EH�yY��yP/����������GC6<�*:��A��%V1�
��/#�hA]d^q-vE>�_߰G����c�Q\|� ����i���/�.s����J[�KL�x԰�thՇU����٣%<��^�s������ݴ�:z�lc�$�F��h����h�w�����0+�}����Hj�K��)黋�9�2���&�q"ﰌ>�7̃�\�~�ĦE�-�]���?�Q1i�_#�Gt�!�S:/�26h[�	��(�X�
���E�nD�d��aCeLǠ!�o�fK?�@�m�1��y+���	n����SA!D���cǼ�2/�&����L1W�Y��D��]�W�d�(	�@�(@�ߵ���(ɤr�5G�FC�Y���Z���>71�~ߖT�=���{�ezg�l1�w[*?D������Q���0��������Ym���{K����"_b�61{/I~��\^=s�YimoRA�|�K�����Oz֥^#��Dpl�w��K�<�����!pG���:F���H{,?3�{��,8-��X=���L��XU�LJ�)�x�,�r-�dɬz$�#S�g���pk��h�aFb�ɇB�ުt�;����-k��L�m2�8�R廽RfH�Č�>i�iF��/�3�:Kp����6`��Qu3K�+ߛO>�X�xs;u��*f��Ɯ�HQ��f�B�E�|���G�6�*��S�%��-2��P�)���[��oE3�H�j�n�Z>�nĝ�~AH,���Ch�����!�����y�(��� V���:D�3��~��!����*FE��1���@)��sjS�z
��Wrxz�日�#=f^���N4p� +D�a�wi��EܟF���Mv�;�~���Ic%����E�(��))����n"tX���ÇMR���B㬏~��D��� mDQ&0�d0T����i�SK� MJel��&�����.)�Y���Vm��p��S�A`)�"l�nz���A3�Z�Y��Ff���|�in?��.�2���@0���V�/�=Mc���6Z�&	��0�h_˳��A�5oH�Q�,�\#�dtX�4TZ{Gɬ���W#S��+X�q�$*'�FwL�/ѵM�Z�6Y�p�Av0,�Z�B9���D��0L�\�Gg$����N�����s���q���Y�$V���7^I1�	t�4r�ߧk��L|@hp�uv`���-;&W6�ߪ�����M�ȬU$��>�R�Ԫm�����	1���(f��l���{N��G%�4��-9�j���`R�*0=g{�G؄�F�F=��9�:j;"����o�� �6�����'�7ɓ��uK�ĉ=6C��U�]��;��,#K}���q�-q7�N����:��
�������P�A���.k#GB_&(��ɋSnqT�V��C��F$2oo�f ��� �(��Ql� ���Lը]<[U~�B��@��bz�*j�N��BD�_96װ�2��q���=��C����ZV���ݻ�� 5����N�p۷��Fc�H�/�\���o��������nGѧ��o�q�5ǩ�o���0^�_*�O�s��cvxՀ�^�  ��q�$�ã��?e�F2����������
��f�U���I�ۙS5XvP�)}	��u!��%��n4� #1�_��@�|��h���&���ų����E=BB���򀦈:��u [%"V$�����݇� 
Pd��2�9�y���i��#�LR�[Q��@7�g\��N�D���j��?=_��ݞ�/o�s��9����m��8N|\�8B�������Id�*ͯ��h���t�w���m�O��;�c2L�1RLOb��3��:�A�k$��c�z���%��_lы�^�B��;�f�B�K���L;*�_�9���ުwv��s�
���d��ki{cstR�m�%��E�^�Iv����g"=Ծ��#T�%%��{4��\��̪� �$Wn9\:�)TB�&�>L�p-�&]lm�Pվ,�R˦L�F��CH����B�<����Z��+���w70��[]�kψK����r�ܥ��XPbYME�J���X��/왽N�К�� ���n/aCy�E���9"���&�^�i/->N��Q0�a�U�y����4���my�	~oGi�x����nÑ��]�@37��!uF|�ˏ�` ؒ�42������W����!d�����}�`%S�f����XJ�������:�J���Z��?�d��$s	�;;q��Mpl_�-��D��Xy+��ү�غ��G��������a�7�G~eNa�#�Y��6���
�7H�Q)��a�E�;$����jF��Vhr��%Zz��Ճ@P���j��1�"�U�w�؁T�D�8�,�w�XK<��� 4�Iz[{'L�
ZY!:��V=�.��=�
#B�78�'��Qx 	����g�EŃb����ǉn����� Qiz%�\�y,ǅ8(�4�@��vD���ڃo�гRx�8f"�\r�;�����v)��>p�|}��	���\�,k��yke�7TZجJ�@7�?�<q:��=��0��ܜ��^�P�\L�w��12����w�=����z�<p��ԥ��M���ϸ�8ȶR|�����dP��-_@2`]}��;�<l`�`��
�GO/h,����
����P�_��VX�'��J��Y}�s��� �?�Q�W)\�	(��hY�mU �+�[���H����Y��F��Ԋw.��a1t�y�s��ى���0-T�~�N�P�c8�����Qڻ��SnZ�jyoq粿�e��O*��L�+��k��2`��	�%x6 �5��1t��X�B,T�n�<aLjɵ�����078���;��Py��}M�Īλ x�5H�'/�G�<����P"�w�;�w��P+�s�ǽ4;\�[1�>	�'���_�)\SH���]P5�Ǩ�}����I"J���}5�X\�i�]k9�s��+/�P� �<]���2&��^�	�@�L�=�z�Ĺ-�rn*���l��hc�L'��cV�A�S#4��4Wcr���v}Z�����TeGN���s6W�-�B�!�)|�}aK?�����!�W�+�RaJZ����mdcTwc������&�G�c4辒�����>�4:�:y\����&\U��i��j�� K��? X}�&��uBIh���6r�`�Y�u�Β!
v:��f�P�*>�)�՟���	Q�n���"�ry|;��w�Z	�1���By�֝�<��y^�
���(yN���}�a�_���ݧ�L=Q�EW�X�R�l~�+�%1���ۧ۵�B��ݲ"�	��%|�̷0�k�k��M�*tc��u"%B�H�6,�7{��#Dw��;��zx���u�.��ެ�D3Y��S	�n'8|K1�@	3m�ze�r��C�M�rk�R��X��X�h�/$��Ł��\��7,���}\���<��t"��Mc�W�}��	����o�9L+m��K	�u�\Z�Ͷ$IP1�3���Db<�� �Ë��陬�;��j"����}})%�߻�Ȳp���߼z�ܞ}a�1����(6� ��Ž0{׊�(L���������gAX���iJ�R['X�U L���[k����H�eV�T�U�/�Q�Km�x#,ya���������):��-s蛾T���A5����
�B�(]t%��=#Db{F����vu0����Q:Z�����@��1�X�5�{!��À<6�9�M�>�2U���D�[��H7�w�<�
��2�I�2���+b\�!RO��鉂]O��TH�եnD*2ټ���I��r�/��VW�8�@�Wgk?+�́i���CX���{���}�Q�Q���g�Z��[�TϏ�͡{�˜�AZ�j��D�>�o�m�XY�g��6S}߼kY�eH)���[LG1PN->�*N%#���6�{�.a)РT('�×Zr#+_,obI��4S�/jMC�<N�X�B hg��׀��$"(�mZ��Q=�q�H"U�Y)�e�ێ(��2"
���#Q�&p.�;��ݥ�uNc�%Z�/�$j��,�N\�DlGh!a~=_�"����/�e`�p�����	�7�hV��Z�{�X�5�C��%&ι�Sս�[�X�6����
$�� R9���i�;KV�P�C���LW���*6+�n��;$h�D�`E6W0�b2hxK�7�xds���&j@b@�ڢ�G�/?���Z�fhm���1�'�Y:���5���}\�ɺ�/�$��As��Uցh��1�����Ox���ך��
p'��y�e��~���$_�Rs�GzUﻐRD����)�5�3�<%�� !a����������đ+
�Nn�K��ՐQ�Ryx�����786P�\b��ܽBʈ�50����V|7mZr�Y`:m�h.�4[���J�r
��i�*�p\�nv'(���h���:ю����l�8��)��|��Tf�B݀��'a�]!�v7$�ݭ�E�1���́��x�{���7�BB�}Agþ��yA�$�G9;x:��=f���I�!�=6���]��tC���5ĝ2k(�s�qE�>�C�[����6��B9�7ݱx��G����܁�Pqql�e�N��> &���(8	͂�4����
}P�_B��6%O��[�/~����f�M�䚏��N�D�U�dbu��P���]I�$X�[�'�L��By)��|�`�=e��&������x�DU�F2LԶ���?f��6 �a`��+6�T�I%���_������Wi �֮��q(ؔ;�7� '�a51��w!L��W�s����!9N�Z���rVE�=\�-����W�c5��rJ��>h!�!�\O����`�Z30uܡ�dܺ�սW�K�ae4&�(SS�3�����4�H�T�V
bJHe7���X�=y+���~+�JP?��B�JA[�y�]-C��9$ok�纼e���,qD�Ŏ�mh=;��!�տۇ!q���]$B�>\j�p��R�C&�>V����f�3l�c%�GvMn����}'����-�NZ�<k��6L�Z�Wl:Ug�Vx�{�r�����`�)�>lK�A/�;���4X�;~��e�D4��!27f��-kM6K�f�91��e�|a���$14��//i�!M�%�P�m�8�|�����_C/��8!��$Od������?E3��lR>�'��f,�y�\o0 �V�;JTK��G!a��(�`��Z�������@�K[�$ �ݡ��#fa��U���S� �mo�dr��{of�82�L�Adjv���gL�� �M���*�dˑ����n5�1\о���J���~{s�D)�:^�`�P=1(�@$۩u�I�6(ҤV�+7f���k����5Y��UO����.*�3�,�|3>tl��W�-/O��7��NS�!���c4�_xNg�>����N���H��Q�w�l�Dm���cLc�h����q�w��]�~
V4�H�zp�i%�S����Pv��7S��F-�	���jKj ��U攞�B�u�Ln ��| �	?^����+r����s�U�}-�tL2��a	����Y���
�Iږ�)iU�;��5{�*���aɶϑ��>�N�_-4�Ԍ9PFq�ϗ�#��<ۈwƓ@A�ߨiRIK`隫�90=g�/��(���~"v���g��q�9�Z2}�t��(����Fx	�Z��;Y�1iIo���m�C�JWht7���4����^������`�Ә8���>>_L_��I�1����zW"�`qH�;強�P��1��ᾶ�8z`$�y�꼛Q����I^S��7E�>�(^#I���Y����f�m�"��h�Q�\UC�!���۠����� 
��%qMUƩ"g-�t��\��GsF�˿���[8:>��N5���82`[=j�7��j�2E@zz���aj����T,-���ε>%�N����F���3�	�ʟ�'�K81\�?nA�z�aW��|Ip�;y��T�٤�;�c��J�~	2�����g�k��w��OO�fr}���t���v���d�&��"��K3��TM�2$�!��.~tC���mA@���ef@�/6���c2맫B�vۜ�lx��zr���,�_���Ϳ7x���&��Y�מ�R�0�z.�:���SsoΈ�ἷL�?�N��*L�\�=�l<E�����1#mǼ3�\B+�"4/�q|�A�|�oj���Nx#�ZJx�yѧ�]�O��`���Z��b����/}����h�`5�{έW�?Z
�3��s��8nS���m�|GЀL�EX:yA�E�^�A/�0dg4�[M��:A��u��*Ub��y�ۇށp���?֛�'Ap^�
.��ޣ�zd͇s?�$����rW	ۅx�5b��s�+����l������{o�����ܥ��|?Jͣ�K0��=�"�T��L�ߙ���W�<�{oc��P�V�q�~jt�`O4Z_5�u}�
�Lo�t�&�#�*�bܒU0��-�D��[���V��]�*	35�.��f���Z�R�k�v�3.�N��Z�JՉ�>��t�r�,���Nڞ;�[���J��aO���OA<��d��!�kg�Q+���BR�M�.�$oi0[��	Y`�qD���"�^�5�Z։:i�/ɣʽEN������&�XG�j�]�*��2��-��S��uj�<��@�D�x/���7E5
G��J���4�����`�-v�������"�T_��I���p�aԁ�+ϸPƎ����'2�<[�������46�l��������̷�Jװ�4��ёr�/��D�+�yG��\��J�K�[��[�\U�����R9tdne[k����/A��1�ǉ��o����p�	B�m4d�w�T��6�YU��dZ��z��fR=9�g�����������Oq�Y�4{QӿiG9��������iK� f����s5���'�*f�$��ȐY�%v0`�/�9�r���P/y� kȲo����8�|�{�,�t�ӭVK*/o����#�swf�t��c��>l�No��H}�~�AWs��"G�s��tK���ݔP�y��������P��\fv��n7h<�m�p���laJ�G�%P�����R��sh�s���Y�r�Zx���U@e�����(�fK?J{�����i�ie��*b:n�>�f>�dN�أt�d;�Xla�'�	z��˶�>��/��a��o��1KnP�ύ�@��0Q���� ��M��k7����~�16��c�Kg�D�K��]�>����Bz��럢���~�'�\u+�V�wg��N��������ͼ&,6��z_,^�V�R����S�ÏCۣ�BwM�Fp�8D�����{��,o�_d��~z�uq�&�����9�H``47�&V9�S�/q/��W���o��_��mL�*�A8��WsU#�6�A�<�h�e�_�����_�Y��@Ό#��R�%9�1jA�k�ECJ�&��8J¡���ߗnT�|��t�dX�b"A���,3);W�9�Z�h.o-�_���w��,#��ޥ���7�Ϻ���R�+!���i�B�/��+Ԑ$���?�����W���?�����ק�������h.�s�ϗ�K�甖x�M����t�p�a����t��P7���*?�X��~�킠�@&�J���1:u>w�� myy���V�>�ec�a?�<+P+���׈�uc��7�s�˺�x?���)��t�B'�s��yUE��2@��r���l?+����VG��B�6V	�~N@�P�[���E5�� ~��S)'L\�����5���3@�O�N_��w0���F䨟�w/��,�b������U+��}��_��=����;�K<Wb��O؟K�x���D����t��!9ZZ;�] �|�9�F�Q��o��Q;�f S,�k�x|Hv�i����!"U�Y7HSQM��f4D��7��v���1E*j�v5�͚�{O*>n��6߈9Y�E����Jt..q`V|�ٙ'f�I�q޾6`�8���/�l1������Z�<aY`kID�9&Ƽ�.����7�+֗-r�)��!��*)\yq�:�
Wh�z�g�m�~n�����M䇘O[��d�����m�H|��3z�ܗ~4/��Z�o�JCX�y9bߧ�|Uew-����|B������h����~>Ko�KNrU�y�B[V��t����0{��b|�?��Q��"�-����jo�v�܅ۏQw����wO�]���/���d9�ܯ�3Q/���!=U�4
�H�r�M,@D��2/R9�*�x
�$-�_����*�4��CuA >9*��,\��ᇞ�;�0Pr�wD���A�ٳ�XN*ޡ��d�����9�o��l��� �p���)U��/�z�ښĘ��+ja-y�(��'����}5  v��}ɗ��]PA@�#ѥ"]�EL�ll�����	��������P��ADi`� �wG& (���~�������0{�g^�f�U���k��M 5(���{� �Lғ��p�o/��mF��Ϫ��'@�O
���[�"�"��'*�oP����7}/h�0D�N�Ma��
�Ps�B$H��q�'�������(�S��@M0�}v%b�H:��kq�q�׫y�M$ݏ�0�q�e�3���O�V���O���XyS��o���~jf�䁪w���Y7٢�8�$(��4�	��GyiV螰n<�)���3*��	�sw�~� ��ʒL�1�]!�`��_�l��)#��"f'�Rٖ��?<�O���]vۨ�R�{1��������R�3ܓ�	C/Xl"�ܑ��XoҴ�ƅ0UMwxv�d1Tz�"�rP)9���,%���L�q�.s�19:3F�|�}�������������ߎ���������hi�Q�Ƽ���q)�~VPZ��a�i[�E��O�$�Ҁg͟Ls9�mO	�H�?���/�>NNx�<��V�?�弫U���x�����-����y�C<P��Q�U45�D�ϠH�EQ�J/�E�*^�7AÊ���7�3���Y��ᗼr�2R�!E�QOб-�BZ�U�*m/�(�oK��k$4��k
<�'1h�$�"7�ܿ�>C�"��p�@&�:��>��F����D�V`?�q�T����'�y��袗4y��� �a�n)pm�yf��.�L��b�"D�[�G8������*tY�z�EQ[�;��� S���b�yF_J������8h�wݑ�jH, ��!���^���-���(3�X�����gӡ�����\<1��N��QT�uw<<(�����)	ROWJ��ъ��i�����B.^s*|�>��]�f�P��R�!�xw -��,0��X`Z�=�t��s�����굦��M��+m
�lY���϶ˋ��u����2�e$l�[/L�rtm�9�ʆl�W�S���G������^<n�RPq������6��*�'�s ��dp"g�.��#�j��(����g����h��l�yu�I�E�����	*�Sk쀆�2B��9iR�1N�q޹ux����Y�W��Ό�vm0;��T[��f<���W�5��(g�v�(zӳ��T-�d1$*���:mK����v5g���Z���dK�h�!�8}}e�&ɋ=|ݭ�E����~��7� ����/Nք!���%jx��'��$�������q{D�A~{�3�W��$�2��v���VK'~�$�$�-]�B�|m�E�w��}��N��c���;��7��e�?�4�BTM�}�O������R�߾��0�c�Sh�%��FEq��|�d���z�w�[B'F
�3Z�1���	�ѿ+7~pb���޸��g3㾋��F���c4Q�@�̊ԙi�z?�l���Tg[���ɔ�D3'��b�VT���|jR�i[{,�a?BǢ�L�b[%쟽N�rp�n��]0��+(�*r�>����용�v��N�*��hT���@� _� �E�yp0 B*�dR�<���jS���'}�f�sM�,)[&m��R��vS攁��Gp0�Վ58wE�����WVJg]b���l�T�6��fC�a!^Iɓ�����J�co�w��T��	1>l���Cu��˘1�.���.��CgHN@���Ȫ�.�v8[>�S�I��ֽ�lq+%o�z8��Q�F���3�k����(J��"�/?�z�q�����2^ͶD�����ͬ;%<�����>̉�:`�ٕ���'��� �/F��ޘX�Qh�+ 2�̊��F�!JL��˪��6㣑�]�*0�{�R��)m��O(*2�7	@�}�>���b�b��zw�h���<e�;.Ø�-5��L�N����K���pHF�VI~����#N��Q_w/�T��s�F2Z�&���t��d�ZM,�;�bAq;���c�fr��X���8t��r��@]z=G$o��D���dj)�m���K4��!zF�`�"�B�qT��m_ y�'�,�b#;*�.'4��s��(�Ρ1�vO�-`�J�U�3�c�3�`6s��o�d�Fs�1������Aǣ~��c�gs��P��:KpZ�*-�����v��i�tLA��.�5K��W ź���l��L�)�H�y�k�_Q�r��5}CET'�0�����Mg�T�{�ֵ��w�+�8`��F�R��[f�.1?e�� ���\y�n�N�z�e�T��ߗ����[���p-�4w��m����co���.����7�������c�l��0_�l��\nq_f� ��:{�{
Q�\�ߠ�$��룁A��i"���砛�˦��Qǌ��϶��/�Ȕȱ�XI����pR����ǩ��#Hc��d)��hY��M�q\����'�͌�|�S��2%�`\1B�4n��a�Ƚ�z�=&{P���K��֯�R��f0�wH�aK�s�y��d���%�d ����Y����)�2���Z]:4�ys�D�ID��Z���/<+C=��T|�n�����(#��D�Ce~):Mq,��xk��뵂q��x[�' ����=���̉��x��*i����Z�H#W�]ڵ����7��`�"�M�o0P�=`<z%�&h_p�6�_;r��.�9+��=��g�՚���-	���"�������2ž���YS��@�9Ɨ>���>A%�N~uy+��,��)�5��%V��z� ���DR�K8�y����6���Y4I��ߡ���i�d.,M���b�$*I�G���>TrJT޳��)�΍v��q��s
�i���򅊒��8�y?(ms4����^��u���\���ލ\���:��+ǳ~��Y64���>pc[!�R��2�=^vK��"P�p�&ّ������&���Bz8H;��^] NFMlH>Q���&�dv����&'���h���B�SqY��,*+`��.�Ҟ�W�e�9r1Ʃ��f4f���T���I_;L��要F���e,5��,���{�)�u�z$_`���Ca�JVV:^T_Wl��+�|v��{6�ҵķ"����;��=�B?�FHל-�{��o��pjݶ}Ie�vyj�#G������]�c��l��ۘs7����X�s�����D)��"J�,��5|�0��t���L��СT�H#N���������?�q�?�)#��fFt�l��/�xCa{�x�e�b�O�+ϼ��_�@}�|��8"�!ng	V���ɱ��Yv��w#[C�fD�֥T�r�6ȧ�!5��=�R���
.��haJ�_̣�V��ߵ���,�^���l)�B��:�c2C�p���*T`��6�r�4�=г���(7��y��UCL�A?@+�4�����t�h�?�.W�����'��˶���6Cs"I�!k?�j� Uot�kM������K��	��eh�
]%��$�x�Nn���$�Vk/�9�g;G�k�;ݓu(ɻ6�LK&[6��
x7Z"�[���ݢ�Q�{Ad���a�d�HBH{vc�l����J+3�:�:&ȱ>ݱ���h(�rޫ��o�%,�{��Q���	P`�����Һ��nC���]j�j������G�~˸ye*�h��zZ%K�Цk�o.HN$�s��� �'��I���n77O�T����q.���^�{]�Ks:������;���P�ָnAW���\D��W�gl�p`M.]��bP�S���$�,�_s�$o�|ZnN�6m:��×mE��o7�DL�	z]�_��,�������1�G�F�z-x)�V!5��_�j	�x"�zx�J�M�X0�V6�|�F�m2ؓ%�<��խ�'[r��c�gj�F`\�i�f�g����m�l�_�uQ"x��8�*��LM,�}Cy���V�o����*S���`�9 W�:P[�I��hF�.�3�kg����A��W��`k���m,���=W���e��������P,S�	1z6Y>�J�L�|ʹ�10>iB:��Sz?��c��|��i?�T��U��m��@f썶��!ndq��P��.<BYt��30%`�su��ZX7�b}ؽ��y���^o)~V��쵋�1�0��X���z�e��^���%*�%I��&B��OQ�����;�<s�Q��mp��2-���kP*y0.~�j�!���#XNs[Wʾ��{���c,JvVTV�����ъ_rk�q��*h�"VCX����,����ʠ
�A�d�e�o�Z��������ܷH������<!��I%�>�U7������7��/pL����)
�f���H���p��d�4�t�3��)��FK����#��:����ZXBۛe�T���n /�Y-*!<����\5*���4bx���g<;"u�!�����+�bI�H�`�j��'V��g�����5W]�g��1^�@8т���D�&�Z.g7���+�O�5!�P�9Z���R�J���*�J��w�!߼��+� ��T��EM+����n@�t3dD���aF��1��pJ�,�]p� _pxT����I#~7��'5�@B�GEF����*��9�}V�گ�3�*���>g���R��I[Ҟzb�����}��%���bE`���Q��(�,ԗ�7�BxWk�Ks�[�2��)��S��-���2��E�)��v�*�A����������$�!��chr�	�mL���\��b�ec���S��bet\z�ǹ��"A�YR��*X�ڊ�H.1V��dĺ�Ε霟)����%sе����gB�S���G�%���D�ۿ�P�N��V�pN۵
Wd�$��.t'	�_����t5�y�㋕qc[���҆�.������_J�]�wS�����7���W��3Aۋ.�����>*�F�0����M����zf��i4��񙺼�~�bƆҧ��-�D�W��Rv�n����_N]*j�Z�&q�����]�c���k�r��)~	�Ѫ��)O��r�p��>��]�j�	��gx#vh/��pl�o)�ך��ٽC�0S���F�E@ߨ���dT�~jV\�5��h�-"]i��	��k�{Jg�`����V��/�8'�l���H��K
��!L����晪r�"�#"�߀{�+��Q ��?��8�DU�i�L�vޥe�+UudpW�^�!�Vl̏~Y�`��yB���=�U&�Kun�d�p�ٺ
C�=e%B��N���{�!˳P�����vQ�)8��}z�V�f��ǧ��G��#�J�R7��e�h�B1�Oز�= ���
+�N������}�$���cD�(P�iCg�)\S��I�%[�9^��A\F�ݺgk�_�UF��<g��^��4��>D۩�(2��5�|k�6�uh��FWR|��[���qsk��jJH��Yޜ��ɷ�?G@��b-ti��Z�ξ�)���a8�K���� ��' ����?K� �!�l�$�$
�yl*�8}Gҡ�o�i��m���Յx����[� >o6:!���`��4�?���N�~�I�=-��+*�T{��ӓ�6mfD5����ם�sg�"����}xGDÁ��Wq�,S��A����fE1�^�~0����n�.~y�+l��?_�;�1��Q�-d	�4���y�	��N�w�Z��Qj�+��=*�&�9�]t���@ķ�B,����	�]�9s4g��L�e@,7f?�Jo�*\Z�z�my?�������i��( �-�<P��{cv	��}���R+^G}�*��[u]�@���m�@�m��vL۬�����5��� �
j�Ӈ��3go�J"���X����M�{u>�Iƿ���I�<��#vQ�� :�(;�6{S��,�Lt���,�ٓ
��p�:i�G �!dL�.h�c��u���:��F< �[�#��@=��[}�Re����$��b5Z���9�.`Y�4{'��
����j���s��=��[x�|,�5�;��Q��
��<� )cf_7�����ֵC�[DL�SL�y�CH�}�RL�����~e-��OZ�Q���T���]0P��Ť�K�W<�dڰ=z>G;g�؝_���I���:��U�١K�t�En{m���	z#ͯ�mƁ��9�6{&�Sq�E���ip��D;��i�q"X\(�Z���}��jm�5 ���Q������,	�8.�Ն�Ѱ����>�;��,���6�v�.s�FJ���1�c��?��o)��0���*��u�N��j4�;�LV��X"U'��c*td�[���~B��#(�󙖶�L���ӹ=	�R��E�׾���D�3}z�a[];�P���T^�8t�NCh����TO���5�/otW|m]y�DX�$���HPw�h�"W�y�pV?2�L�Fi>��[���Gw��5�%?�狹Y��	޳��-hY�bS��h��H�m��;��(���8�)�>�����A�С�LW@��Z��ݞ�~�v3�ٜ-2��fّ���� Q���ͳ
Y���O��5�����g��`��ʲsă�ZiEs��
6⭲��ν�D>�3��;���y:���I��T��ر��lNMr����=���8����U������y4j������I�]'>x�Y ���[������
' s`��U�t�7����*Kʃ̩:�+h��Y��}'�Zd��F�<�p���y��A�&�E6+����ֱf�r������7��c�9n
�tV5x�(����:�<y%K��B�f�{���"�-��_�8���#0È��3=�L9l������-����K;�*�gh�sK5 ҉Rq����!���ecP�t���oGT��ݍ��ߴ�F8ky�ߙ&�x!�$��e���Jc�w�0q����}� 	�牍C<�5�u
� \���_�8�6 Kp� f@�b�LrC�9�9���T.��h�����̡ֱJ�/ ��ӌ9с����k �c�	�_rco�K��f.�J�@Ɲ�+�yE�1'� ����;���R����b~�,�C�q��H��Ǣ1׶$�<�!���8��I�ތg�f �\��{��G�쾙7DƐ��`���e��r�،j���=�Ms_o0�
��$h�{��~EIyW*���<���k�B�=�"f����,8����s��N��3L��KƂ@A	e�5_�P^��J
e����-�����2E���qv�u^~����e㑆����14��U|fV��r.�,�aw��x\яVA(%Q��{�Q�����1�{����K@��{�G\f�BY�g�ː :#���鞌��x�	��Eh�X؆g)��7�{.���
LA�==���X���,%����g�>P��K&�yI��?O0_��YKW�d��r�߳��]�x��j����a�P� >�U��H��w�q_5�A�,�mf�� �6�\�07I��p�����+�M#�b mb�7~�ZS��k}1��~{�V��x+�f3=�+ɯ	�5җv��T"nӁ��������[z5�g�e����ⱒl��(��F�О6o�Ҁ�p�����dU�Uh1�]{�W�t"p~Gq&�Y{�"e����0Y���!I�׶x)����u�b�2B����ol���	�QIw�	Kr�c1��4�F3Ü�:W�����
�/t0�F9 2��g��sg,��IBʘt�f��q��	���@�O��/�����DEf�$��gҶ �Ro�����Y-��D=�� 3�QR�P�q2t���`J�Z�����[!:��*|^ 4Z*Hzde��֯4qvc.�/
(p	m�ܮ�2B�;���)�;��߹�Q��M��ڈ����E͚�	��K�T�.��yDnQ�:3����H&��/Z�υ=�iwγ����T@�����C;��})�z͆r0�t-w��W͞�[y�?�md�-m�C��Z�/�~G���q�c@��Hp*�c�	�u,w��D7J-W J �f4���/ �?;G���bS=YQ���+���FL48jgVU+�ZR�_��q���+,W^�W� W�A�Dj@� ��.�Mf����f�M��*�+pO��ּ�N��!s,K�M�@�V��'hs΋���$c�tL�W�Q���[ن�}�������ӛ5�s�����[D�'17/�1*~�=_Tf�Y��Z�&՞��'Nv��PੁP���ĥ 4�˿��|+�+���x�V�n��J�N��pa<~��+�cK`1'�3!��^����W���Qd��2��? I��M;ɧ)<֡~^�*��4���� �{�G��A��ې|^>P�A�y�(i\Y�c��u��.C�V�K��b�
 �q���(TA+��*u�V�N����D��b� �c�]���,N[o�֨F����b�+,�f����T.��<ʍ�>�V,j��h� ��"�����3
/Zһ���|�2���i�D3��O�}�K�2?wyEJ�1Z�o���ێ��o�*@�|�k�BZ?��� �ưW�%��|����[��������=H�,�OKhL3
�[v!ݦ�Ias>A���$���ąX����KƦ���D�~h��e�A���EQ����Ʉ�	�����0�.�<��c?|����ʮk�ڙ{=�ZV���-+��]���*3ǀt l���ݱH`�ժ�G�nӖ�zM�O�Ub��D&�
�&�Z��aOu��/ۗ��I�CmɈ�KĶZ����� %�'�����
�^�ʊ�(IC����0VdͿW:����U�N�Ie+h|j�{G��}�.�&���0�a�W�G|NJn�F�W2 H�ʨN�1�"2�F���Е��b&U
ZO����̭hAj,���6̨��+�o�Y�W璱~:�=����ܝD�6^��8�٥F�a(j�%��,|�)S�	� �r��?�f�+��>
�vjr�F;���'q�z�~�k�-cœ=�:	��f���!�[$t����gtr&�|�_��EV���؃��:��|T�m��:TÐ����Mt�h �Hals��d�ZT�0L}��W�b�U7�3�I4��U�Oz����}�z7v@����N0�9�h59�m�s ��e�d���S�O�@u1-儫�O��;	6������h$O�/��d�]ضODYl�ߐ�R��K�_��a��b�[c,\�-c ��m�-Mq�ܺ1����R!�k~pp���yC�e��>_��K��QRi��LNk_��rڐ�	7��9V�jZ
�(���y[P!����
a�]��4z��d#Z6�-�:�f��>�,�ږ���޽8���$�vIL�)��Z֟G��|S0r#Qg
�`�^PY��2��u�W�F̼0e���Q�2p�H^Z�O�6������xn�g�z���=@@�_e�"�~ǳl������8��6��/���G�T�����j�*Ex�ro ���S��D!ܮp���ط����
�7H�n���qф}'�����WI�>��#.���9�hQiL���tӞ�L=��'��2*��K{��)�Q�
��?M+еU.2��Uo5#���mX�l��޻�,�%���1c����M��5�V�;4D�� 4|Ğ�,��Jv铦�O�[`��:w��V$���N�⎵�y�[�	UJ�ް\c̹�I��b o� q3�c��A��g("�<��F�B��=gr�hx����Y?��r�W�4�z5�+y�O܌ߡX3T���I��5 �#T�Y�4!m����@W����¾��J  G�D�u��B�L�g�BM��R���j�ģ�-i�Ù`\����6ӟ�B����e����1�Ndѳ�:�]f����ة����'���Kn���ͰK�q�H�	�=-5����ƮS���������JT�Lǩ����\h)���&��k�G��)�=��#I��`�%��ջ���z���Qn��H����@ǜ����PK�������ڶ�ݱ�$��̐�����������1vBx�%7&�	o71R���������4���V�o��������
�L�"���sƔV�rTI���Ek�Ͱ�:`qy���V��	�������'��럏v�Z>#�K�G~@r���V{��|Q㲭�k��>��ǘwx�ta��i�v��f��O�/�*6VɆ@�l�=3����qte���Ä�֊����-��&/0�X���2&�=��SV�%q3_��*�G�Da��D:����D1\�$	�\���#Tb#Ԝ�p1j��k���_Yi��I���i��;6�"]� �k8����Ȥ�'!L���TuXs�.9�V�x����c�8����A1��4d6"MM�O����x�+p�]���,��[��'���F����"��U�ݟ� 8�9�X<�n[�z�8��{"�����rPN�U���n|3�rp����;*��Т%U/�3����;�S:Л������;q��:%+���*����/��3Q`��8k���k�o�^�")�^~.!G���S�M�Dc�����i�\P�_Yl-v�&�Ha�nV/����9��\Gj-��H7��H=�0hZZA&���9ڂ��sA�ӻ���E�\SXA��林�%���(��)��䤖|cT�N�X�"z�v|�j�nL2�?�J���A���p,3j7�\p���'xi�d\؜��>���+��~P�Oj���:ߘ%��G�?5n :8H���by��|���GK�
���f�p��~�]�Ca��Pܕp
����׾j�����5���$`�~����٠�t[1��i��.t�ҵm�Rџ��*�U��4%k)�]��q��JY�x�����?���-@}�:��Ӽ1\��ɪ�xP�޽>P
׎c�{�}X����2�)���u"\yr3,�� � �9��/LI]��Ԃ�F(D�����[�/��,g���	�B��S�1D(��^-�Y��s��䲼�f�X=���CQWU������&�@?���$+����������9]���b���}��w	y�N�Ez��eS�T�=d��j΃�a��*�
k x"��o"d ������cp�j_ӆDꆞ� dݠ���t�?��:V�^���Mmq>	u�7�`�T�"�g��x�aL�
Z'8�[�A&��J~�S�P�� HF���OB?�J��|�|��%TC;�cp����cɖh�
��wF���i�(� A��:�Ќ;�z֋�b0�Na+ �������~�r����{o�ѐ!��M�D	QdHg|b�Y̫��:����{���h��2#�?���k-�$�ma���4�Td�\�}�K�;Zͬ�� S���'������[�x�p��nm��2��D�/Ϭ\��M[�`���n�.}����s�)��gBΞ���B�O�xN�w�!�#�0��L���a{��.�F�*%y��-���x�5�s���=�_ESJ��|�.����i6��ns!�}y4�f��b�i��RR��7bPp�F�uX3�_k�o�PN|�~4���GU�j��i���e�X���f���k�o�C2����x.�//Wa���:O��M8��?A�J�i6őq�%yMg_� ��x螡�?�/q��d�W��:�E����F�R-�^}V�@�����EH�L��y8�Mq5*y*��KnaӍ�	ȶ�g��e&/���=n���#�iE~�b"�
��y�ہv1
�@woq��;���e�`6���T[��ˍ�Y�K^�:�������4�PW�M���(��a���c�K��:����u�.��nv4�V���<�m�^8�]�u�x��H�[��rP2T-�a���}�U12˒DM�u[�'v�)�s���k�%5���c -j�u>�����UOfr2􇂥�T
�O��l�ϝ2dZ+ ^?���B�^�3��?��uWlK���7K��_G>泄�Ol�Q/��t���q�넽P¥��7��*l��4���Ȅ��k�U+;V�H��/�ӈ8R�s�/J��A'���� ��:��T��;=�C��j|�>Pgϧ�ö�`Ǜ�oe�uS�-ӊ��g�Hݘc�0�h8�F�R����o����|y��Q8< nw��۴h�GJ�������C����?���\�@$'��e�!�P���
s�j�'�2�%~ދ2��C$G_���#�Q�v��
��7��ɻeA2�zz���'�\K����5!Wl��" �N�k�y���@�"gW˯;��fn;��T�,��Ⰹ&_����a��AJ]�w�p������y�������K���8c,a�4'c�X��4�[#˔�|����I���rO�IV\v�;�s,>`����Kz$s�T�ӷ������%��	4�Ŷ/EV��Ym�`^dѦ��(�,XA`;+��1�r� d՘� V6YM"���?Gx���U=��I��!�P��JjE�9�jzߗu	�����o]J��g���@:�lö��iմxXBzpaG�K�aJ�P.� ҧ �H"��5H�k4D��|����Y�^M�r/<�~-���,�x�U��G4GneC*��bٖ����������Xq�M${�!i9U��H@�|]m�ϝ��B�m�Б(�@j,����\~�r_�X��?R?g*�$l⹼Mg�s�����@b�m�'��m��ֿ��� T|�TU���Yu=�2J%��k�_���H}�!��u=�6�pnZkQ��+II�z��p҂��_�w��y]W�ͽ�D�yG��O�k�#�]o2����{��N�`�KS�]��h�Xg|��ǃ�n�V��5��-��=Rl�T(��Z���� �Ρ��#0�ִ�;�5�xa�W����u�x�m�~���6?<N�������r���@)O[����E�9>*�\�G���e�H�U�zH�*�=���95��Wnֈ�r�iW��U:�F8{�{:?A�7�F�W,�ҳ±Nr\TQ�z���VfԠ�Q)V`��I��i7��������%�ʢ��U�f�,6��&��WWobz�t�B2tf��cj81����Ny�:�G���:o{*~U�$��}9$�,���eG�Y;�0ǽ�B��/1��)%��Oyߑ>n�Uю�1H�b'�,��Z�MTV$�YWB�pC2��D2�����ע-f����Pl�X(Ұ=�������1S�X���b���iEOq��Cp&�]P\�B�]�^%dk[�}Xy\/���J�Ɉ��R�S�Nۏ	h퀅��r�?���_����;^�۷�ފ�c�9:)�Hw���n`hTb��k�!�60�I��Y��e�YF�^�	�.﫲� is�f=q����,�M\��m�/�AGw�h�(a�7�V�����[���CpX]Y��H�y�D[�sUqeC���{$�#" ]^�n;saD�b�Օ�ez��]�pQ�Kk���(Hϼrt>��(��@���ժ���(�ڲ�yN���z�m-*��Fi�Y�� �\WxO�W�6���<�7J˨���;��'d�{���ﺇ���%�I��J����W×1�@ˍEv?�K@-�.�^�p��a`�1���I��->�@p�sl��nfˤ�E2٥�V�:g;Ӑ��������*��w�!��I�-2E�ހ�>C�D����_��I�x:���������4�X;B�frU9d�ؿ3�>f�:�n�����dl�=E�-�xr�?���Cz7���
C	I��Ť��o�ي�E��zAz�f�Q��l�"�2q3u
�y�4zú��ȉ�(r��&)HK�{�y�{�n��N+�]�ϠR��5p�\�M��Y�c�a-A�t�&���ɽe	� ��.�'�xT]X�/Y�?�.FJ������Nq�Y�l回_�7 �}h��w2�p=w�����\e��Ób�XYiBj�a�x�E����
a���g�r������m����eL-oCk�#����T��j:��xLJS��9� �Umo@�Z�jM���*p�[!��+i�/+�S����ף�;cqS�|5F�����®6	%�xa	�d���sfVۇ����d�M�����������-c����t,>�Z/���Ҍ�s�Z�f�9I���R6>ѐ+�C̷��	#���%ِtY?���=�.�,�g�����>\��ߞ���u���uh���S��&V_+�R\0� �b���iZǢ�i���b��=��(^�5_=���H��T5Q�˝�w�Ҥ8��ԋaB.�
i�I'��7���e�D��x��� ����Qt��}<�;���yY����4����9�YO�lOF�����l�����@F �*'ҹ���C~�uDFڞs�wC�dرU�����_�7J�}����sqW!lj�Ʈ�2�Qb�|C��ɦ���9�IrVV���B'�t������"�\������(̦����o�A�=z+\�	-#O��@�VҘ)Փ��P�����������k���P��G���
�QgB�)��z2�\oR�5�a���R��UX�7&
D�?R����ӝ�
�*t���*�}�����K5�&��h�ӪE�s�$.�Rt����i~	f�H;k�逸�$缷Y�q��q�޻��e���%�`ě��1[�8������0�Sφ}��P���ڟ������L��_ߧ� Ա���`�!%�y�qNV�By�`����%�chm2W��7��9Y���Ldb������ا���B�l0�W�h�`�*�ja�;�O����iz��Ef�p
��B���Ń��LC{|�G�~Q2�������wy߸��=�<��2��o�eĿ��|���lA���s9�WK[��ycA 8�	�u��W.
���F�z�֯��-��zlX�oaK&���4�k�J��i���4���ZTu?�cjveu-.?|�G/|�H�J��;^�H��[���t�������!�j�H^ �Zq&%�6E'~$��%YO�O�i�Ժ
@nW~\ީ�/�l�Y5��Zc9�\�%s����lCŕK�~���m@�)U�J��n��-L���Ժ1���3�[����Ӽ`��9\�{���Š�O�NM��h�œ���%ǣ>t���xFO㘗�f�))�.��Z}��&��� C�+	x+�ד� ��診-��zݨ��M"�� e�\W �;*�J_��Ao���3�T�JƼbt��&)�Ƨ1���?���c�����u�+C��������߷X{�EߥR�LzF<�0����X'Ѐ:S\w�ߴFmHPv�K��
=�ʉ�����V�k[t�m�9�f�����H�F�KK�ͬ�/i����Ur���zxU���M!c8xI��Z��<���B���d�-�,[�����㿓��z��8zd��oeOu7�����&\�04Y�;�XHZ�Wg�N��+&�Ҙ�1����l��s�3(Ǚ�bd��� 9+4@2���7�=O9��9ǵ}D�ke���������z��YA9,�7��Q�d��0K����&n��J�ȭ�{*�ۈ�$dނ)h�Ԕ.�M	�����聯
w��$��ఎ<Bo��gWڸ*����z�gl��
l��zH�$��9��A�aI�ֶ�b������Dǁ�D��B;�D���X.�U�驐M��
� 1������o�{:�sۂ�D�v�G�|HU���DC�`�q�f��v�^@1]��?"�b��Rh��ݴ�|v9��J�l}p�)�7ow ��+Ƀ|H|�7��f�=���8vd�z�HG�{��68���*����4�m"~c8.�;���f�+ǹ'���f=[b��<9�-�K�ײ�U��f�/t�sF*N����9�Mu��@rx'm�������bChj���W��c�j�x��Qx�bW�*��>�� ���Ŀ�h�P��dӠ�VjdI�:���e�I�鷓��*��Q3m%O�x	�=k��Q_-d	z������
�Yx���3�c��������;�i�9�2.��p����g��n�����­�G�D���w��6��ܙ�#Y������N�[�t8���߶9��i��Ճi�(���-���K�������k���p���W�P��,��6[��!u�����Hx���߰6�v$g R�2�yu�솕���v�?��t��j@,G|���8`�Rw���ƣ�y=�I[Q	d|��e�)W�ӏ\�Nm@���V�;nu�:�4��r�x��d0$�d��߆��ݾ|�X5�Ť->(�
jLE�fޘ�b�҄�'��HHix��h3�4+7uV�^:S7S�W�Hʬ�ٿ��Y^�Oo���1m���dr��4� ���X	Jm��"z:�d����\��-V�	��-Ѭ����t҅-kΙ��_$�9?y��C�	."�8�o���Έ�vvR�g@f�P)8x�/+�wT
4ɧ��*�P8B�纭R�iC�\��4LBYG�'����jw���5���oQ�}��&ݢ���&c�:�A/��C��_��I�I#��3TGO8��W6lE�v�����:�|D��,�F� "����Ҥ	U4�����m.�Ըw�6���^Ũ��uڽ�3�
:��&B.nKww���ٵ�F-p��3"����c&�
�ע	�u��z�4I`$<����p<ו?�����E���|ct���'����)�"��qv8����
��0��޶�ۊ8u Z �%6�Uo則$P��\,|���ᾴ��B
�$�T�
��ga��hzŜN=[M?�IQ����3�}�T��F��XQ�v�.Ϝ�0�)A�R�xhL�5��c˰�������N	La�|l����W-ÆC���;�?�&��+�m,ⷚ6��`�(�*2�4���!�\Kc�y!�]r	���L��puL��9\SG������kS��k�VyࣼW�^����͡����(C����2Z9�{ٽ���jr���3+�YýC�H���� )4�{ٓcz�_LoY�6u�火�v2��J��op��=տ8C��*�Ko�-`^��>�{�QJp�\"�Z���DT@`��x�F���.�
�g��_h	��� .�j����a�`����EC"�L�B-S�+x�w�a��F�Wݩ��X�ܕ�5F~:�W9��R'X�bDH�H��� @�� ��!S�yC=.!�������ls�{����Ї�<���@�M:�k��e�Ӫ=y�~��G	E�12H`%c<�
�!��, �����l%�FW-�l&"c���wpP3Q%��}x���&�/�㈱ش��>4H����I���2�I��ZrIQ��q�n�m���;�Ğ���=��9DD{E���vě.�k�ꍇ`7Q��cP�M���8/�$���,�=>��&>?#�rD��l�a�P4=��jx�W�$Hc�%ǔ�!��;��\)Xp�,.OSzvXV�_i,�D=��)6y��>";�g�Fа��Uz(��������aJTH����ð8J�7\)n�5^���0��<rf��d��6���
�B��z��U�$z���wTݏ%�����招�"�v�dW�4?��e�x�,ו���L\�,�Ei �N)�ΎW�μٛV2Al�PŰ��Γ��'l'R�	�T��aԦ�x�A��^�go�[.��y�����ۥn�������d�w�����r�.c�%4Nq�z}��R�.�B��|�Ҙ�%n���A�!�v�o!ԉg�1U�+�=�_"Jlqt�|���3{�_�⪐	�h�]\�t�k�h���m�H����g����/�U��
0kq��C^�ī�J��6����K�m:����R�D�	��"QP18�q��?"�Zϝ֙�N]����??G��+�?�l���O��s #�Y�G��J$@Yr��t�1�A���K̽v���<�}��N����]�I�ߖG�0��8+��V�N�M;��w�ݚ�ۓ����hd,�Z�F�C]���pE*�g�/^���i�9GҜ��]սP-��b��l��1��;b)4"nl��0A;8��<���170��ƪS�r�F�R�Aa�")EU}��}8_~)�D�����D�9[��3'?6�����kx���X��W��9K^��lgqX�d`'���Q�Sz�C����7V4f�������-���}3���`���K�͵9W"�F\ �I ���CP6pQx�oV��)�ƾ4u<dØ����m녗 L�,�fmk�A���,�s�;��b݌>�0ϱ�ͦ@�����OÎ�%�R]�%�!��pr���O�c(ft�@���:�cB𢡖���Ũ��Qu�ݬ���_�`�ծ'�9
tSM+�S�<7,�%w? fab&K:�>H����S�Y�Y��Q�[�F�YG%�ؚf��x\�8\3���t?��hgmi�6�!�h4�#��<�w_���T2��wK���7�g�(���[�E��>����Snے!P�W%����xD�(�`��dS.:>Ae�>���U�A�ޓKKӟ2
�	1����P�������~�O��'�x��Z0���-y�bV\/��;�$ZM���(�!�Z�v�2�f(�\0�]>`b�rtdĴ.���w���.�t�S=��@�39��Y�i�(�(�ԢnpȻ�Qf.��.����dQ�S�F�G��B���#U�f��c��%�&=�i^H^R0EjȀ���gK�A#�Oq�<�>�*2�}v�me�1�s�����ߊ*��{��í!����Bt�[��K-A��ȼ�L}9DZ]����]A��]�m��
\Mi�99�\��ְ4���g�, %i,v/���D����K�~��	uxڥvg���y(5�р~�|��ge��Q5�눗����L���4�@@�H����xc��ĦdS�
,9�MC<�S?���w5�Qk�v�VZrg[�u�Bl��&s��g�M���;رXO�E�$EJb<w��;+�$$�Ă�d�ݱ�]/6�>/��L��g0�l�ýS����,��g�2Á��y�YT�PXƵ.�.�֩��_��s!!�~��\�z�A/��R�~�����t |��.�MݨuJ�6l�pu��0E�<G�=�=�)�JWW)�s[�9n砻��mq���|�(�L`�p
?Ho����6��W�d�i�r��x,���Հ�{Q,�mU�Z*f�����ϑTX�\u�R7��@*����1��X�	5�L�<o�O��w����9t�f���M�.si��9jp�³T豪�殌
Ɖ��`,G��W/�`�s���Q�i���a�QF�J�B(�jO�ŀ++Ͱ���mi�u_V��f6ek���x���q����
�X����5}0Mŧo���!�ƾ���l��£H@�DO�p�T���#.G:!=���a�Zӊ�^������
碊����WJ����4x��*ת�C_<��{K�{{��,l~��S�OZ9��s�<�}_��)���/�[��:��m7�!O��q��.d�E��m�ҮoS��x
h�e��a<�Fb�O�U*#�d1p�Έ!u}�HU��q��Z�)��n��Lb:�㶘>��V޹Н����AUw,����x���Go6Iۺ�����r5;7��^�F�
�*����D�p�����1�hc��3��2U���5� b%�n���'��h/��fUq4�a�*���	p��N�3����.s��?������Ch�u�������m���d�OX�n�x(PmN����>e�;U��"��]� x}�cO�pd&[^ұ�t�De����2�Ϊ���}�o�E�[������)��������k����B)sci_��΃����&�n��И�
i��?:g[�?AN75��f`i��M������:!~�Lo�{2�s�0D���UX�Z��>~^]�����>��C���A˝DYo^�.k\ �����6�F̈́�b�^�-|�t�LQF��>3UEѴ�/���v�C94E���r�$Fö��L�D�#�[�7��u��X�t(�i�Y���(����� 5����N|	u+��� ��{Ğ=c^����e��;1u�j�\E��U��j(�����u?�{��[SքB�v��M���r��c3�\z[��B.��+�B)��(����C��U�|��%����T#/i�t_hF~f�H���6�/i� i_n�C�-[��|�CK!J�ރ+[�����-��?zC[��j���JO�.����([�:jC�+�D��0���oˑ=H�=8�0�d���Bg��[��YYß|V��u���L�#�U�U����GW�3a����8B0Rl��p _��T��w��c�=���N���!�0Ӟw8��y��Y�qH�>�h���4��C�B<�Aۻ���P'I{[��l��dX��*9z�2�z(�~x4�M%�����$���R�w���3A����-����lx�p4�4�<�pT|������K3��)�m���dL��҇�o���#�GQ��}F�]��!��Fv8%�5��*��"+�!ƛ���_VZEr���!�Fϟ�%��4�ŵ��g`�7�j�zxB�V]B1�v��
kI`F�Z���
�ڶk)jݶ[" ���I�!=�[{�k{f�S�-oɎ₵u�v�䔸�e����,F��ۊE���s�{�آ-���+�87�!轚�ӕuKl�
���:
��3���8ژ3��g�aKBs�bS�"3Y�A��� ��{�TQ9o�3yL��wr�0�AT!���u��R���_"�dc��	[����#<Y3"ۣǮa �ԙJ�𤺜�M�s�w9����4�7 @c(�#"��|�ۈ_�j��@-QR|�	�i��N�1C�;�%Ŧ��5�暬vR�42w�H�/�Xa2Fz�O�i�w�]ҿ���xq/7�8�0�56���X�A�>��t����d����/�Җ�������*�6�jQk<4 �֠�7����o�сp�4Į�0t4v]����p��;��R֕z6�(�n�Oa[�g-ꑉ_�����˕�^!=����B�{���OA ��yx�$l_�̥t�ճh�繉��M-�C�>}�rg��ţ�c�&	"l�B���c����D���Gs�Ek�,.�/�<Md�y�4�fL~�J79�zFp�Clp娃S�| ~V���@�h����N=0kC�{Q:�� lĂ�jY�����h��BR=�+!j�����|o�9��[�#n�w~E�?\=o�R24Dn��cZ3�a�(���_sY�\�/jԴi���Ϣ�|�ᐟ�34�^�Dv�U��#d�}k;�΂74_�A�Az�I`�����2p����G��(����3�{�A�ѠB���mH�<a%����#@����@"��׹�C .�gD�^*�cʹ���췃:�� ��H���U�;�qLuZo����贬��@���S)c���C���y �)����N��.߽Z���ѨVm%�˂����U���=��/8P��������Q��?�$2�/|�l��2Պv�uB�2|��3&�����e�/#/���tI�yw?����s�3a#��Q�zP���|fM�8���	 ��B �ld�!��-�S��w�7�DU��P�Ĳj�b�߇~�Ƈ��+"6���}.�����yR-��o�zb�y��u^��ȡ�M��a�bO������\����娍	�m=�w��2�䜏��-��=	�{��;�rU�4�+��*��p�v���m�[�Aڡ������q��M՗�!�f]�t�*T��f@�����(� _Q��z+L�y�P\�B �֎T����o�?)�@�g>r��ʍV@N]K�D�Mw�_���h��V���#K׆�9ăڏU�3�a=7��[m^��u~��3G=�y�s׼��m<��i�v��p��E�M"�|Ux�A�}g����5��������f��n@Jּ�+V�:V;׽�'\Lŕ��$� k��B8������(N�c@�W+���B���+�d6��rR�6�YVΣHhx��̅�h�$l�Q���}�躖�R�Q����R~�W�n�z*�8�n؛�4��ܿ���vZFX?Yǉ�Ʀ����d�\7F�� �Q ������GyrB���iغ[08Y ���HM��<+�N�G�9�
�[Ͱ6?8ۓ�,�O���(2�-/9~���������c��9�d� i�ab?w?!�:"D�W"�D�+\��Гrj���Zv�&Ei����C�����!��=�.�$�yӿl�OV8�lnG��GЫb4���0�4gU��k�����,��U@�}HL��X�mZ(|�B�g�������o�B�}^l��ÁrGn�5�U'涷��В!�Ht,w���At�o�k��8#m���D͙�{��A�1_�7	�\���xl�.G�Bʢ�I@P3H���p�uD^U)|Eg@�JP��F崝uW��������C֣���Է��!�]��}�ҒC�	�Y�� �9>�X]6����셐u˝g_�X�D�����|A(�9���|�@�ц��4�>x'{h}f�$����j?��D�N��m�+���K�������-�#� |�#��A�->�:.�ie=�w�De�O�P�A�2���� 7��,d�����!>[�jc0�Ci J�o\A:��~�,qH/�����T�:���
iq�tK͋ն�(p�~α��^�� 1���r߹��r�?	j�u
��V�EU�P���k2ܧ�{��fळ�7�2c:WT1gB���!�_��28 �i���1۟=yN���3s��T�� �0��r�[��3m�6����qgjUnλ�J1����v/D��"2w+�M]�ɪ���� �����;j!���vq�XUȳ�ˎ��:A���<[�i]C�~I���+�R�2���}�D׫�x�Eu��ɄD�pe�y�:[�^�3�˃�7��<N�)�Bl7}�=�	8I��'_�/���lHd	���TT�p�= ��\e�f([�tpE͓�p;�c��L���nIQFQ���U�b#G�N�}5ð�/��V^���}�T�}��F�L�9ڬI��i�`D��aB��gCʻ�(��?՚Ҁ�pP.<i�}s����Rmâ�	/���g(��N�-�Nmc�R<�C�"���Q�j=`>icڍ��p�b�QeT���<�G��l���4���J������9�x�N����c �u�������"`��C؆�֤q�rʋ��S- ��EKZW�\4�K���r�X�`+_�2 A���&+�8P���V�����aq�8�Y'�+�Ôu8�Pn\��/���ιm����I�ω��%��
�H_��X�I��4F�&+�-֕�?0�Ū
Җ��tx� ��*����N�hc��r�Mj�7�?�9����s��/�Ƹ�΀��ᑇ�ZM-i)o�;N�ہ�(Yz
��=���8d�@��yo&��L�R�ؘږo������e����Q7�h��]��W�a�UuS��lh�?Q���33]����o��|��˛��$��e&�����؋���Kk�A2f��v�oGQ(�+RI�t�@?K���w�!#V59Z�d������=����	�k�;�
AaTX�B!~��~o��,Л]�@ާ�*R��J�8�H�:������l��[�̂��iGI����6C�+���F��q�7h��j� �q���j�v���B���9BK�!�!�"�C�lV��M�w������&�Rm$z�̘� �p*�q��u��u�e,H��M��.�7�CH=���Q���9�g�[�����:�+�6�ړ&[����BR	zWDҺ�qIX�i�[f�nM�V*���'����D��M�5��Jߘ��g(��y�ۮ�{E����a�L�9�=mټ� ~!�(�~,�_ܞ&�;�o?�t��*��������(io'�R�#͂#�p�dXd��4^P"�[�D���k�Lޠ+HU#c��R*B6�I'  gLC��f����yM�T���L��Zy��A�&G��ǆL9�|'&���r�i�$5�g�z�DN����{;3FRr��Q��Χ�GH�+<�ynó��c�jx_Fl��L�xJ��C��߹��O��֏��Tw��wh`�}g��O��Rz�%1��3����ϓ/2�<��%��}�����b��N��X��\tkd�rve�l�h�λ�f$��7�(-�~�ʱ�+.W�x�����[	p���اʜ;Wk�R�yӳ�.z������¢��?�Ŋ�ǔ*�4'�w�P��$WӶ�����y�_Cz�����K�.%��ʠV��
�K�41+�2�e�-��ϣp�� �a+�0��ʠ@��`�(�ć=�h>���{�qS�V� 1S��!���l�E�f���a��@�S��#��'�9B�Z4�=,ɒɓ�w���>T�F��xV@�ГR��6��ℕ1&M�DoB�
7���oe��k�7B'�,Ř�' �6��)�x��=���@9ۂ�����>O����"��ʦ:�Yb#y��6uM�	����`�{J0\��8����c,���i��M;���=ۦ�'&��;�g���,����{ފ��y<�;Fz31���QB��ݲ�9;��"�����fh�`{:����w�{,΋�3��@\��/�
ԕ�TU��d������տ��~^�e��9n�m�&�����8|�GN�K�;r�~�m�P� )�����ˀGI/ч�y/|O��R���x@
˾����3r�^���J_Ub��T-����1���y���k�]�b�չ�Rx3~;_ֱ��-��UZ8��mO7��~-�>�7f�(�z��똍�H�S�:�;��#/�<���C��l|���}#	ͤ[�;R+�	��o�����
���a���'����;R2�s���挡T�l=�;̽�+b#7P>��G*�mʗ��_zr�v|����|'2D5J�+%Q8�Ґ=��м����Y��@A��������;�?�_yd�N;�KNe
F����F���ʵ����xN-_Z5G����F���Y��٤�Efii)�������&\�� B�Be���ē3G�X8�xfw0�ۓ�5r�p�W�콏v~!�����)�S�k�����Hj���H�}��U����g)��%�[/��,�V��H��|�d[��otP�fl�:t"iּ��*�������Ư��y2�=ӻ|z��Ț[�U�%�[)OP�(��tG����ɱ�����k/�!���7�1`�gJ'�8���F@ዊ�CN]>��*~N/��5a�����CC &��!�p��9عt�)R>�&,��ENA尞F��5�8�a�"_,;+�h#�")5?��)���BK�#�+��*�Ym����-}-���x�l#8�j8��$�ԩy��� s/\�u��mv���n�������O������Q^������9F���� \��i�b�}�����<L�{=��1w��ulsLwI�!�h
�n�kӎ`�څym����
h�a��v�ܲ=S���Ϡt�ŕ6�kb��(���4Nˤ�4�\<Fޠ���D�rk��TE������q��6�*���W��%�<�JxN��.V�"}e�����Nk�q&��Џh�U�߉��;*�5jn��\�����Y1�j(|ul�w?��Ēw�4-��w)�K�ݷ[**�Z���'���+��y'LLu+��w��G
��,Qs�k-������hݱ4�@�z�����ĵq�͉j����SEO���q��,SBl�gƫ�6)�)@�>*��� �@1���2xy���.c�`�_�+
�|�'x�r��7�|�w#�K�>���^U�]u:�^8`���������Mo�a��Rb�&��.��#�dY�1D+B�A���:�u�ˠ/J9�h4=OCR�saU�{C���}=��>�hi�5��h���Nz=<wԟ���՚k��M*�ǌ\"���	��S���� ?Z�|� ��D�R�1@��n�U��&K����ê�a$�-]t'�j3D�'	�A���W��؂��2�,c�ɻ6��g��57쓳?�!/��6�{�z3BZ�,����='@x��Ym1�����b�+C���؄(qDx��{�M�H�PzJ�`_ɐM|0)�� ��z]��h�} o�����dF�3Wh�{e��e���rh	��G�*�+�y���VJ曷�֪8���A��v� a�V t�#H�fg�1�f�_F���6�m�y�y���=�)���)�b��<B�\hj�P��sd�ݧ�D��2�����R"�!���rJA�$X���h��	����,�c(��0e�����N����vӖK5��_�T�1�	���#{v*�s���<w��^@G������1��O!��C;8N�7�BY�����f)7�^�C��v�M5��7�8�w3t������}������������yg����5p?�#�Ǽ����	!l�\~�����c�F`چ�Y���v�ʼٕ�QH�? T8%ˬ�r&�*$b�i��
��4$Q��0��OA`r���J���|D�N���>s=�t�Q���>�:A��p_��7׿;�,�	(MC���x�~�Sfr"�c�k�YH�<#�RZ\p�z�9�w\����e��vfaE�DCE88@�}�kaFN��)����W��Y.�M��y�V5�0����3���)��)�8��`d4_�j鲏t��0A����#Ғq��?9Q����!���8�p�T�Z�!��8̜I�nv��3�l�и5�[���J��,���[l΅	�gLtbٮ(51�n�F�5�1������d��1�h[h����OfW�I��18A�N��]�Q(|Pl��놎{ϻrz]L��C��s:��l�U�n`� �����ߕP�y�Zc#F�\q��~m�`8=�e"y��݃�~��?Ό���@��T�8I�D^�����ϧÉ���	�?v#�;���%�Ĕ5�1�w«�6��M�u�t���b릱hW�Fψ�e���`�8Q���_��OU��|)m���$]� �-m��F����x#���#b�r,Y�f���΢ɤej0&��L�Eɇ�/�%F$p�g6g�Lh��*EŢn7�^����N#��>�uP2���ig:Y������-���� ��M�ﴔ��C���0��o�2�r#�I�~��l>6�E�����|�2����!�9:BK��-(�;�`�[�ɵao<9��F����Pɩ͑�LJ>�95j�zL_�y|\�O�q�Ħx\I	������̓Vl�
ӊ�Tӝ��}����d�)�_;w�>x�L����v��I�Ø3v�I��w���Oa�*�U�_�2���^��M�)��$��NSt����u�b�X�w�fٛ'�Jy��2�LX�(�"&Z5�?��)�#��W��k��1��/�Y��i�dQ7��*Z��8%�2
/�Xd�F[]κ�qv���(�3,�&����������*N�9=_���JBg��൬t������ךLz�T�t�U���^}��O��eК����#����&�d�FY�%M�g������LC_���	d�r�;�qW��|]�,g�
"��BFF�γ��4i*���9����E�Y���,�e�ZI2�Y��(���عr��������7w�k�ĝ��9c�Kn_g

�����r�*Dt��F�4L�n���@+�>�]��Zg�+5������8l��q��X{���u�,,������94�N����U�_I��of�`$ǏFR}[w۲u���/�{R^�n_��2����e����<fa��>#���.Du����G"�zHi~�*��?#ӱ�K����S�;��3�
���&Ϣ(6Ź��4$���Sjk;�L܏�����}�Z˒���|H���-�p����v�J����כ%9�$���'.�\V>7�5�>��ȼ7>��o�݉�G(PM
y��Iu������R<���A��?I1O�uZa`��7@S��_׻Y��~��c��ai�)����<����&���U����ܗVBl���s�-)T�}��wR�������|���5�Lm�{�����>;�o�od��o�8m���՛[qߨ� ��ݏ����#].��OLq�p�iv�Ȅn}��&Sc�Qo4%��N�,표��
Hz" ���Zh���^юiFb�7��ˋ�^��n�wo�[��}L��~`VE�� [�OX m�W-���p�&�NU\�y���%&�o�����e�=�
���-�e_w�d��S�ղ��ӥ�?W�&v�6���+������GDBX7�Acy{��>NT��;T�MM��Ok��E�[TdØ)E��tMtThW�Q�*;R��W��՛�����6e�Q�P��^�h.��Y��r�@�0��rBa@G	*֬����O:]�����FD1��6��3t ��6�}��;��Z����W��N��p���ӷ*W%��a��Ng�ݺf��<+:g�A�r�֍�����"S?M%/(0v�$!�'~�cמ��m��'%�F,����/�TK��C:k�X����g,9�R:���N��F���RL�m�W	���:��_�#�~Xr'9�H���5#�l������=���5��	{x���ුx��Ut@z��"����m|�SNЦP�bnȭ�|��ND������u����g.@�m�*ʠ�nટ�����sjk��( ��g/����7�o��H$�<j%�؄֋��4�_����49b���l�+�h5W�=���`�M45"�ۛDNG����
� ���$⦳)o��T�ؕ�9��_�g.�K�ӆ�	��	ON���jx���dBu6�$������ӛ/��u#���(�{/�9+�zb�޶��e���re�I�2���]��&MȔ��qA���V/m�(!�@�����p�%�e:4�a�J�Y��+�s!{���c�(����ֶ֠����vg&�<J�d��j�<�e�"�ƍ`'P�6JEwv�T�[H���b!F}mQ='�3�s?�@'d���r̀�b+ E+oͪQ�����N����3Ou�����᧓��%����t�&�ti�?�%��U-�b��!L�5Sm*��ݡ8n+s�cda!��v�-�r[��yۥ�F֫zM(��(h��\ˋ��Ӥ�m;Tq���:=K'��-O_��dC:B�	s��k�������/����"Ȃ�n¸�8�����3�����]�?�e=O�"�m���9$�s��@�ֶ�-�^% ��=9���*�Y��_�B��fC0y1��xwL��l���W��'�.Ӟ����%N�gIOVݴh%�PmB�ɐG;��M��ٜ.%ӧ9�w%�3���RR��JZD&�)>�,H�n�fii!�pj*������mM *�6m�je�v���(�Zqj�|�Oy�/Q�i�.����"*�B���&WH��q1���]�/-HݬPR1��տ�i����O7�i�gy���_�X��mE��#�n�J��G��o�1oT\�+�!� �
���m��E�"���Κ�N���G�5��.��I��P`'pn�_��p2�7���	�����y�<�D�_`� 	:6�亇�čI{�o��1N�֔F��H��)�5�Ledx$�@�l�Q����r��?�VKt�	C������bxpշ� �40��GO��'v��>m�_�V��f�ֲ�k��6S���!!�#0�Af��C�w���l08f'2�c�5w5�
_�zz�5����׭�#�,�KR�����F79c6���Sqy]���!hk��8�%�Ze{�PF_9>5�i�*z=Q�=�h��b�W��=xtY��JTs������)�Bj�%�����$Z���K�	�ȍ�73�6F�mA
$��0�H2������ȎN��+fͤ]~q͉a��@F�4�e��xs�p��*��@|x�H�3��Ru_gw�{�Y3�$��d�*�� ���iRȣ&BQ?�,U]�c�9�t��g4��@�q�-,_��w-ҁe���	� B�F&���˘�9.����.� �����e�u����|�CM�����#_�-dl��>�&��d	��L�C�V���()�k����r�k'����jHU�r^ਯ����@ܲ�&M�X��Dzq���cn�=b-i$a�b����ӈB��at�}�a�7�SoZ��hZ�"�V��2*��_ %\nm%a�W56�A"�)M�"WA��R���+��~u�['��+��s��ϙ	��U��9�r����D�\�	�&�ǺO�T���9k�P#<Q�%,�!+�.�:����@&k����f��� �Q��i��-�@���5ɟJQ2�"S&(��^Si��ӼZM�ԡ=��I"n��]��_l���dH�{���m����X�MXg���y�OAd�,���и^���Ԥ�e�v\��nQ!�?��e܆zOP�.'[!�
Q�N��Wgya��H'�����4]]JA ���,
Ws`p]*o=@Ohs�|��Y��9�I�x��;*-���pC(@������h{�޸(���H��������̏�|�6�ԺA�X!$*|5ҌO��M�U��B3u�^GL`���)r$*N��o�^�����ǅ3W8�Jں����[���z"�I������;]G bDv��%ј�T���Ry�<'��e�a��R��57[lK���:�'�H�z	���0TKm�	�Z��T?�ď�0^�q�F����>�#��#�_6��|��ɠ����G��XG�;�{��P7�R��I��|�딧hnx8�)^��k��c�z��#^���,���~hbE+v�m�
2�k^DY���@�|�1��g�ȺIr=\axy�}��i����^�B<�����O
�Aǝɳ�u.55U"=y�2c��;��Ǿ�7�zY;�B"��!a_���f'T��!UE!��u��	1Hq���q��h���*��H��W�ĲP�$^�7犖1x'�f���f�F��&�>�͡R���,� x.Ҙ�-�&!�Y.Q��
:�.V�?a�x^�o��kf$�&S�d=-�{�.�gum�v%�o��b�(����'�ڠJ�B����R�8��]�-NG�v��NWSh�[J�H֘\S��.�K��?qkֽ��=���P�)�7��ndC�U���QZ��7���{/��
�}`&����� �ۑ��3R�~���������|���$Fh ��^����Kʽ�Q�Z��Z���;��!�r��3�g�a��<;=���i��ʓ�iEz&E&�)������{1����F�x�㜆}$c����[o�(O��!u��תR7\�*����8�
��9Yi{�Em|���"xzh�I�'Fl�'�wgA�O��� ��)��Kpǃ��Z��$V�ƀHo��/ɒw�2��	��wL��dxZ�%���%s?���' �bP7�?�)&�$�!e^���o��V^:$������C�@O�7���10�l�'��AfC2�}�H�c}���T�TFɖ,LͶ
 �YՌU+H�?��ҮP�����2�<k?u��\S�c�k9ʗ��������h-}��{��>�|��{�˼8��n%]�>�2����YGY�Tk{;��	`₁@�Z2T���]uD���^��LaB�^sլg���E���Y��-���J>�@����Y/C-ғ(6_��\8�a%'j�ӸwLAhY��jz�;�2�JV�p��g&�֠Y�x�̶�,I&�J�)��O���Cb���>�j���h���No���CI3����-1�hi�.B�'��	���2��|N�h���tI��ء�v�w�y�$��n����Ps}��Wʻ�����[a00~�б��;�!�~� H�y�|M�A��l�;���_2p_Rf�>0:�ؼ���.f����U���� �5�qP��C�޸��lUT��$��S��wU-y��3��f�M��V��H��r���Y���3bίN��Q��P����h��kf}�3@��%�&b��gaC|�Yޘ������wU��Fw�D��JM��t��C�D)Q�i���ه!�ɡ�#�������ցA�nI��}ZzC]��9&"\`������i��U��RJ{S[p�IK���X}�������(sL�㢓}��0#�c͊���k&����Ү�'#X�eD^�;�����wn �'�U�u���d%�ө�5���W���ZoV@@���נ͸n�B.�sn~�,>0�Ar��y!��CN�"i&����J��������>�~<:s,u���hp�	�ۑi��1��M�z�ͣ3����p�9�;����kh�b{��rن�Y��,��-���$J�.�<ƺ�N�S�G���Zخ�}�z��@b�TIhB�M.NT����e3�C��/>�`戴7��:�� ��^E�J?�%G�:GܛK0�6�Fe#�W(�gS9`�kM�H�F�6u:9mV�sH���&���#g��r�F7�!uw�2G��=�{M�wC���Siq��c�NCDJ�����H�@Ґ�:�f���������K��a3U?(�i���8{��7�M\��� i���!M�K\����)f� �^λ�x�-�*<��?�?�r�a��
���%��Z�츇 �<�ʶ�]�:�����#xj�d�p���l�nV�<z��Ai)Dyd�S�]��A�U�TV�/B���,-��~��%G�T�bl���-���kO'o���1�2�T��/���s~�*�y��{!.z�7б)��Q+b���s�E��^vj�)���A��OɎ�t�d�ӺH
f�v�;m��L�Q͍VJ&������f��n�;��?��?���0 ;�j����=oTb	2�{���_���n��Q���UH��-z�N��v�֌f�=��O����e惑@C��$���`K��І�=�BxI�?��4�TE�
E�S�q�B�`������)�?0��l�����|�O�ҏ����w)���4��O0�ꗵ6���2�Q%�~Dh�8`�`%��?��CY�Z}��s^��v���l�՟��kbu��3�_��h-;�):��+�K"�ܽz�NEu�&K����xFn�2^��%���׭�|d��ǮN� ��N��k��js�a�L�T@�רW�V���QwIF�a��Zr⽷���P��� ��f�V��  !HO���(cb�Z���y��դkG�\�-��/�5�⸞c",�k��^Y�5�D�7Q�cW��'P@�v\鳾��]0��4����
����}(��� ��N��Clr'��ć%j[�f��1��3;)wO��P�Rh�O�L�:�0l�
<�I��Cs�r
٠aR�*�TV�?�r˛�N��UaҰ��"I�����{N�dq��[D�-�!p3������9YT��<{[ڊ��X�[<>@]�dy��Y�E��Ób�j��<iO�a���PR�^�G�����l#��J"��c����>��y�?{��3�X	����t�츀(�j��#F8�1��qV�5�U�f�Uq�P��m���2��v�y4�^�ɾܽ*+0a�k�ϳ��/�7Hy�w~MSVz7ce��D+�8w�l���c����"���F^��b��_�άx�VI�_)�����G{ܠ�Mm��c�i��m#	T�	ke�O�I�����c~�T��/���0���r��!x�~�VӒ�4� -@l��$��V�3K� _\���:��2lFV�J<FI.a�Iw�W��x�w�)�]hU\d��S��Եf8TjRV���'!�V���M+g��P���.�F��_ė��^��`���5 S���+��Ib���*�Q�Lq���VfAˀ�Az��PVߎ]�R�M�����ƅ[	���o�x<?rW��ID����/���^>�"��&��*V�|����X L�ǌ&O�Mwb�j ����v�Xf27�����Ҹ>Z�&�y�
����c�z�:{�łO?��
C-��W�v�K�I�:�e�n�e`A��ĥUX�<ҡ��.˖jB��E����!��܍��� �{6����-"���λ �=����d{�})e���O �+Q�z>�ҳ�Q\��VU)��VD��(������Ȳ�$�i`��˙M�����:�JPS+V�	�q%~�x��]Ke��L�~�lN,~�C�'�TJzYz1G�F�_m6�����߲h�YY=�B�!4�K���a�C-����B�G����A�]�jv>� ܐe��:���$�̝㘨�y�9ޗ.��C
{r��L<���\^���N���a?��r�7s���\%�s�u ��j��9�O~��!Pe��b�C�n=q`Yy�[Kh}eI���@��,�35�J!����8J^�k��ܫ���`�|fu5�r�/Fҟ��.��zg��P�%NT�����cJ��ulr��!�W�Yhm��W�:�e�J-�g���%�����%~�����⟧=%W�`�Q;��r��z�x���ڛ��x62��e��U6��etH�����`��x��>Y��h�ƻY���DK�%"](~,%(�Q���~]{�b�q���%w�`g��/��]-R ��#�P���M�腴.o{�R��]�nj\���.+^��U��w�YBC��)+i�X׳�q)�	�5%� "�f��w��:�=M}L��l$���k�rJsjD7C�5KH���i���_�F�ҭ���9eFO�h���_hK�2��*��2��G� 
�>sE�ߴ��.��~5�.F�/m�����F\P�A��|��V�H{10��p6�\2e��%m��R�y�Ѓ
�#�����Jb�7}��P�Eo��A��:����`��u&K�&A/����q�nQ+���I:kFb	`B����ӑ���%�g��-
��;����Z:�HW�g^F��Mo��/�bg����P�������qsq��:�a��'B��O�W�!MZ&��gK�Z�F���,+��1���$k�Q���B��9�:��"��M:>�h(:���E	����o'L��{_.�\�G�������vؼ�Qu�y��� @�^�ʧ(Y�J���̪�0ͮ~�{�!���N>,綄��r��D�餖[��Tq�4%��pD�v/� U�m���fh-�D� �m�.�L�O*kg�q�M���F���?Qӛ�j��}^>��:�n�Ұ:�;�2@�p��	I�a���ZנH����'㲎w~t�c�c|Ti��phR�=>
Ji�0{����D��6��?�7Oڴ�U��� �s������N�]�����(a��I��#L��=�q��`�΀��%�[�⪾{��W(�ϺS�M?v�R��}��"�K�l�w���Iae�Z1�0�8�Vrt��N�9����A֔-���\�+���z�誝�H]�K���X�?L��kx+ޑ������Z��D�.����G)]�n���� 4��2���z���x��X�dvB���^ �a���A5 � }w�>��`���=:i(��|ۆ^5����e�"�.M��.!WfeZD+q:�JI��C 2CE�Ә�uQ��α����S�9�A�N�p�%��B��H5>c��֮R�G6dQ)�7}L���*��oP�9c�[��Q�S.ŀN#�ӓsKߕT�,����.K�૯w*f����s�V�_�P�7����+zX�[J��slkYEࢶͶa���Du� ��4ቤ�H���8yî=��-���u���F̙IK����jn>��S9 d�|�-������	�N�0��6����o��XR�45F�T�E�8ŝ�O��_��K�nld�?�T-ww^��Tw*ڐM,dFqz��������Q�TC����@2�����TMVO�쇅*�G^����cm�g�m��ˮO�����n�k�q�*��bIr��pѠ���f�P+G��6�8�>��������y�i�JEx-�#m�W�+�!��HMo�O�[�o�����8B�]�M��"kp[��/�̧��np=4�A��{ARq$p�t ExI� tW���2��$S�8�T�J79r�Y����w��u����4�q��Q11*>	v�ʦ�]`�iו�m�S��f�ZV��QŽ'(-�:��^FaH`�f�ܾvAɑ�[|����{14):��n�m��y�[Ƌ�ә��ͬ�b&潃na�	P��=ZPfk��բ�ObC��bq$���Y���*��`�J@��onk��`VH���~�g��K\W�tb)Wܸ�!g�̤�|p�������ϣ�!���'[-@�+��|�V� ^���]B[��ݘp�n-������aU�
<95U�z�
�)\�������6��e���%^?� =����7�Qq�Y_Gdh�PD�?<���<F~_@u:o8}.Y![CQu�0�����z} ���`�Ne�ύ!� ����B`9a�w���'��᭻'v���W�XYܨo��i��q��Р�z�=�SF�4d�9�@Ϋ�鬏�v��W��S*�Pܢq6.�c2B�z� ft��Tl�*x��H��aё*�ڰ`�\�٣�H���N�ߦN��� �fm0��tVu��ʦ�
LIe�22�����I!2o�M~�aC��jbЬ�]}}<�ǅR�(�Rǯ��_Br�",��.y��4E�18���G�B�z�PaA9��Ux|�Wv�k�p�t|?��y��Ϳӛ��>C���HP�D���%��6�G"��,^��1��E����RDX%�F=��]�^��-�S��@�0ǲ�.cy����s��ob/��M�>y��ЕCݸKG�D��:�M[���wv/A,��]W[��!�b�E�G���#d��Iօ%��U�8���~*�V�R�r�K�����ܫ4Gz�}�k٦H��º�]s]�P��󆭸)(��C8�2^�d�|W��F*Œ�&�5��Z׍0�I�5�<�i�P�g�H'�[U�S^�[jbؼ���MhB���L8k6�`\ 7k�>�w1qA���y��P��$�Q���0�}�P�����k�YV�d�B�K|F��,�1:����S��_���f`�v��BH[ɵ�&S�����5��(�+�=-��2v��P����hc^�^X�8���5X>�5_�U�����~�+d��<i7F�hˢh�RB�����׎Y�\�yһ�cV����ӥ���5ו����h���1�
�;rP<N�����Ra�M�f��_ ���c�gdٟ���f�C��:�V�}�2_��c�(s��W�Q7��/[
��޾s&��G暞�K�u�<4�=�i�g|��?Q�����$�����[���+Z�������E����S�q�.�jS��%k�����_����+��!�^��ŀ�����Od�o
e*�����Ѵfq��ֿI�C	�  �@�"��@,�ly�դ�q�	(��$K���s���
m~��z5���yH|��6:A�!a"�O>��C�����_?��tQ��Qv��cӇ�gƝTP�yT}��G��	'�e<�����h�eHR�Î��<=�=�@����H��ز�<��[��
>�P��ɫnp�(y�t��;ԻQq��4.k��X��!(���D��(���oǳ>�n��ˀ�����Sk(�[U������4=����63ޡ��q���76a��Z=�	��"y6��̱\aW�Tr�,>L�g�6u����>*ŏ�*&q�M��og���>.E�Ȉ��Α!,�¼���۴��W*#LK!oL�%iDր�l�7ڞ� ��O!Vx���+,���e,��<A��-�ȁN�M��<�a*s�&����-s���S�+d^������I���o|R�Y+`�o�����-���`r��r������ f���xA%&��C���}F5�eΈ��^ޯ�X��Ԓ2�!ԖU� ȗp�yoV�Q��M	M];qu�����Ye��q��<�o@
ӉQţ0�����b�넊�V���KC� ����n9��8k�F� ���F��¬C�Y�(^L�����s;�����*��cةs�%v]\ /Jz(�L{���lv��(t��4���P<����mkbr[�#�,�B��m������h���l�ͽn�եSAt���n�W�ݬ�6W0x��It籨(�J���N�|3�j���U]����+�Y���cS��4�#<���Kz��b���1e�9��E8Y�D�~�����-�b8(�u	�@�܎u��m�A�1zVrϓk��@�3����5{�3=�[��H=�����A}��r�sE̤H�T�@s�*I�̄�����g;3C��${�[ű�1�Dk��+�JT�+�'n�@��P�a��J�y1�z���@�q�����j<�/H��l���B��SɔbyEߤ֢���n`��$jdqh���G"zy�Go�2a�33�;�s�v)ڟ�]^Lќ�$y>��&� ʀt�LmT���u#��V������57-���y��?9|JA���"ϟ��t�m�Ȓ7V7HX</�hC�+B�ټ/���C�8+7v��^�J�ZN� �����U˟���x�����z�؍d�
L{�>zo��e�7�.�8_m=R���,��(��S�xt0�N"����%.գ��r��������E��$9��UE�m1n*�q�잶��7u���Erؠ�BC�ߥ�}:(p2��e�G����	��͵���"��0Eo�k���=Գ[�>.[S8�yDd>Y����N�l�O��՟���0��L�x�ΰI�$O�x�O�*OT�wA������O�|'�����ĳ��6.;z4�ɹN�Kuý��}�P�ǲ����x��9h<G�y�u��:qj
���8Kb/�'�����tP�V�l��Ҵn]����;'k}h1)���(����\<�~�~�,.N2�����{7�^}r��< Ix����7��1�ba�5x5�g^�D���U�쨶�]�I,�~�[�ni�ou��d��C����U�^͖�^jEkcz-�!�U��oܸ9�f��"�ϒ������WbRQ�op�^�W��y�>��� /47+�0��Ƨ_�F,�I|���0%ԓ�������>+.��F%1����ۥd}���E/С���ϗS`�ˡ��b�	�f���L�U<Y����/��SzP���r��ᡖodD2��.cJ���/�T�;�ƒi�~� �?�#X��8����މ���
��CgZA'�������J�F��aQ�@�;�2����8<b��U�$,�9؈,���e��z��x|��}����P�:#1�a�ˁ�:��l�TH�
?�
���	��Ґ/Z����'����V�N�d��g�m�2h�@y@�J� �\�$���x�&�_��,r$����RH7�.\�p�EӔ�O��O�,tT���y@f�n�w7M&^��>�x�_�)�X�H�� tJr�?!<j����P��b�V�n����ad?\�|L�eD�+�W����B���oV�D[:�`��	)i���~õn�!2zF��K���]M�RʈQ�i�K&T7[��
aG3�{Ba�	;�Ǽ:X!���}|�(�����,_��}8�'�f@&A�u���q��xvHilr���Z<���G�'q���㷤�(~��29�46�p�I1[۸��g�� ���!�⠪��E���b^�e�S����|_��{j��|KB�t�T���� ��H7�C�r� ��N��-��j[���T��S6g9�0�芄�T[��#�M��S�: w�0f�r��r����M�>��ǂ ͖�V�dVnW,l�.)>��	��9:#����X0��d��i� ��li����*l�H��Ю�,"�)w�!/ʯ%�owx��9����n3�C�Zn
���˾�L�t��稇�98>��ˠXL�-�4Ͻp�?\��<�&�2kS��� � ��@d���=��4S��2�:��L,Iؿ���DeTB7r�ܳ��1Q�,A�O����gs��P�����?��TJ�1̽>Y ��L�	D=X?	�~R�?���P�8��Y�M޸	���]�"qd��U���� ��n�3�m������g��X�^�8�LO�%m���D��"��l{�IЅ�QԸ���t��h��H	� A!a�����Ɇ��B���:�c8��ك�i�����=+���G@�K�tW��&k}�Ik#����n��?grZ�W_��׍a으�J�צ���5���0U�|�_K��3g,�~@�T�d�O1���N�m���J�a�t�Ն���Z�,���w��lӛ-B���X*rxy�"�O�=2*��k��x��T�,�
?��e=��D��?Ts�k16��ek��io���IpC�:�J���� Ł����!��o�d+nt���[>|K���۰�b5K���dQ��
  ���L�@ \�j�~)M���\� ��(��P$�1:�������:�~=� I=f���c�C��̺�/
7>6�����P��YTGg-��u]jp�H����hq%#����}�(������Pn�RǨ~��e@�'�w1�*#ӭ�"������5!������X�W)���
����S���f����a���@oy*�Ȭ}�Pg���%���-!�S��`w-?�s��q�R�D� �?D���=Z��'�鎽�UC,���*�5ʠQ<��^�&;ѕ7 J&�yQ�8����06�`���W)_)0��{f�O[���x���"*�Ck���_:�?X�R��~]��Z��/�n�}����߆��{�!�r�{N�bő�^�R3�Ayy�/6�MN;�����_b� 
e$Յ�@߰Ƞb$k�����y ���n��0�qGY̬҄Μ"��6(g�ETk�O�骀��?f��f���J��f�p�~�z�,���x7~f���Έ�!����I�	��mH�o�=����PH�*����}��E?��t���?	f�>?����{Γ�lV5Sx�����G�;�[�"�!2P˜|B.���*?��E�E�sM$	e��Ľ�L ����ypNv/���贅R�PH�~PrJ[7ˁ2d��Om�f2�*C5s��h�B[��I�
��j�R�o?|ۈ�[�@�T�u�۝>m�� Mݞv��p��W�������X�w�(pה���q���|khF�j.�\F�S� ���\|��}\M�;a��	D�HQآ�=�c\�3K�p�K�im�A�b�x#LO|�v*�r�w��e���L�a,:b(�M�Lv5���?� �<�d��YүG�=ۖ5��Է��M�?���2��XɢE�,}
��m&�
�4�����j������f���-IWn�\E���g�N�}y�%)}�5�O5H?�}��d?�?孧�������O�CK�x4����^�=�UVt&��^(}s?�ԕ�D�Q��l��Dp�.�^6"�^��W�t�(a~�= �7�$�O��1��ɕ���]��b���-��2c!��l}:n����We����V;6��S���.��K�����F�Ȅ��~`�c���>ε Fީ���=����n�������ׯ�+��[�2fMr�z��v`��p�f�rޱp�n���}�L����#r�j_.C⤎e���Xt��]�<�ڂ~��"��<>c�J�"��ia���P��6�4Ϣ��-R|�)Z$O̥�l��u&�O>���̐>FS�ѳ�?�a#̎�h�R"�Mճ�B�b/���$�:��!� 2�(6�u�y��j��T���b��:$w/��#���v.V��e���vc�]��.$Bi��a��܍�2	/�a;����\�ӘW�Pb����%�Q8W+~�)��hz���Nw��wN��;���V,E� \E��E�FW�T��|Cw4up m0��*���g ף��r�	�`���#��)�����R'��"br��0~q�Q5���Ǖ
h���l�&`E��V���E�L��;�Rrk.&�X�g�E��K�Ǥ1o@��2Gr�+�<GA[��:Y�k̗�Mg6S�m/�o�i	D��팀''��iG�obbn�C���>��=����DFG3�vۢ.�ɉEz<k�{��+���������F�4�
|n4�siTf��5��G9�Ş�yu��cC�tW��:<)c�R��d��R'<	=�⓯]�y׹�~�q�A�O�X��O}23F��J��`i�}�*r	Q��XԎ]*2Γ.%Ә��Ro�5s{�pdl	��;sMؚ�7��g����i��I�Y:ņc�X\�;c�m���G��$�;�\4����<��5<k]�~���߻��?;9�L񏷠o�LXXΉ������ v0Cc����}�%$q��y׍%�C�xyZ��p�V���@EL=��쉺{���Rq
DsN<r��=`�^*��G	D�mF7v�R �U�aG�f��*�h��¿8\]xV�|�����ޡM�ܯo���s��x��dkʢ�����W��YB�s�@�H@n�k������>Xm,���[=l�p`�!+���0P�o� ��n+)�<�tH����$e�bQ~1�/w�{��"���+�Z3[����/	4�ǽ���Ơ�׉\�ZN��J)
�Z:�N]�w]��;o����A�G�|��>ס �\+�~��/��ѓ�ұ5G'�ÏǄ��s{eI|�oP�h������]��3��B��^(��x�sk�B�cA��}JW��H��S���ೱS�汳(�T�+����Q[����3u�Y%P���ƞvE-�p�����a�0��=j����t�%\���� `0��7u���~��N�Cٜ����ϋ�1�y����w��˗�`�*��l��x�u� ���)��e��}��y������3�	��i)��j���@��"
�6���O��z�׏�v�Ү�h���1_�g5��hT�g릥�����ߨw��8F<ր�!�D��m�F28�����Ӕ�H����-{�7�x�3�Xs3 ���s�P�\�ͦV�I��~|������!�/b
�U<H')�k��f�@�ZH�Z�c��*$��НVi�%qJt3f:��-�;)`#H
h��{NT�X��3o�������L"�L��G
^���7sD�@��qׁ���_L�;��DA7�U��L�Ȟ��`��ed#ߖ��n����}OՅ=�>v�>1&FsG:%�9h�����n���#;b�	��g�����,���A� p3C��K:n>)�(1����M�G�e�I�E���e����RM�bzk���Q#rV��m�CY�d�0�~�G��{Pt�3%��v�X�3W�rX��w$pE����ņ��T�(M�%鈳/"�x�XG�
!������-���>�+���Ԧ��V�ZQ\~ٜJ� ��U(��_�غ�9_�t�P�䓮��?丹S�c���,6��f�!����}'-Htl�<d�B��5�R�A�p�ף8�f�"��Mn�!�r� w�DW�3�S��{�B4Z��qJLgڐ]m�F��>���7�4ᔀIn��e����'�t�"���f��6MX.�+��!<�N�
*�֨�P~`ЎG��d���@��L�/�ͺ��y����| u<w��7ܙ��k��u=���#1]Yn�z�x��HGJ��0y�g�%��1��7����+~�Awj]�?Pʳ�3�o�����<��=ZKi6�d�0���������zŗD�5n��;���p\H»��H�a[�1�x�	JL����؁�P�WuD̯TV�o���[by��1�P���,+7�E."�v?��zg!#2�.~��������ǩC(����E���LƆdIV�f^�gJsyl�輸�dyK������(Z�)jBt�I�ͯX�y������t�>�|u��-X���9��B��@���N�pQ���G-���:R[���gDF*$���c�-�]�&��o��)���& �Eq77�f^W+�%�bP�4��/�j{B �$���0������}��\R�
�0߫E�p��c[P��G���C���Fܚv����њ�c�k���k�z1�����
�������G6<�g��N)�/h�w�Q�.�.R��U�l�q�P�旒����͆t��q�� ^>K�$H76�Ra���3#�i�����Lޤ�q�VF{d��d����e�ʚ���С�i���ܒ3HW�`:~�R]���i�ڿ�فP��]+�#@^i�/Ҙ�@!-;�* �A�ֱ%V��7m��$6��K�a�w�<[�HQ��:��*��X���ԗ'7���>���z�$�Q��h3����_\�����_M0�B��w�����0��/.���(�T�X)��Ke3���Y�����Wj�=ɓ[?�Hy1����P_���ӑ�)�#�\�Y�K�i��y�^�^l׊ܖeJ�E�2�"�d�]��Z��M�z�'	��K�Y�&24/���#�C<XBT�����T�|3�8b[1�'*���ͻ��/�`��a�J�9o��~H���$��'�[=���nP��y�m/}��5�31��T �⏮fiB�2��jc�E��؂c\���D_�z�B*�^���3��X1p�.wi��]@�5˃��Dd����f(&�tq��)8���-;Z3�1r�zߩ��G����^s�ٚ�#>���T�A���(����[����R�紺�����({�D��e� �W�(|�/�O�(;!*t3����kS�$d2^�y6�zbP��|Mo�.�'�����`%/��1��sF���8l��,9������n:ɡ9���|P�[�es��,2�ŞB�mmJ��M�r���S�JY�&�[���;�(Ο�2�Aڠ�u�,ui4t/}���4������$,\��//p�3G^�����+�I��v����-Zk�Z*���P�v�<� "�Ԧp��WA)���[S�.>���H�B��jp$TW�I7���P�����:g0��0ѹ�{o?n�f��]�������\�ڋ3���`��!��� ���~��C�����4T����K�i�`��('�"t��[�%�r[���^���mw� �xA��\μ��N�	�y10DNT[j�7|�Vb��
��
E�]�+.(����[!�An���M[e3��W�^IL�`T��;(�"U��0�#�\?2�׶b79��H�Ll-3<B�>'�L�����픈��)��2`��X�L��?j�Ω�*X˄?�ys�OQM����P%"����^��6j�]� '뚻e��+�����(������+�f����g0�uA�bC4 ����,�
�Y�=ζ�ꪱ���T���ؠ��ǋ|dw������V14�Z���^;B*sEy'	E�Ұ�~;��| 8b>��B��<l����C|c2�x�/R��izf_�^`���Xr���Nk�hG2�Q{�7�$tU����ةb��ݼ���7�Ǆw�z�|��K��������Ԡ�� �D�q����O�Y�����|`�v��n!�P�R�����KF^7��&��9�_#��ݤ3��zF�Ę	�e�gJ��18Cl��=��s�rѬ���t�"�^����s�>g��Q؊�h >�����c�<�Lk���+�z;�w��o��.��kS	Tն�(.��;gk�%r�4��K3� �sm�C��7γ��!�+����JMWu1�#m��{����S\���:p40�z^�������Y�
��NS��e���V�IPX��?a�V"O��N���%��b5��+H�_PI�H�8��?s)�f˰B8��E;��Tlm;���1��f8��,s�}� *�@�jb�k�9�Mq�`���4��Y�}�|��;+N��OÀ%됏=ԬJ�� f"������d��W���iu?|��.l�����p�H�y���xZ�VΏ�S8�X*z�B�y��'��h�7n���B�A�����O*���sP, E��{����h���ɟ�R��F�����/*���W';h�����IN���!��ZK��mmޛ�> �Qh�r�
����Q"����H���nD1`�0��D+�� B�_(�{Ō���Q�LT���EgB�s�\		)�6^�ǽ��i9�Q�鎞`� Xnxz�n�{z�rG��3��x�jE����]�^K�T�3�����q��h�i@1f�[ J���,����Yy69<\N`p�=�=�� �m���6��C2o��,�nU�X.5��E���D��Ж��r����poU(�G$g�J#��Q�^���օZu�`GC`l�b.o�AAr �9�nB^�X���=����,�N2㱏8_ro�2�-�0�j��i4bX������4Ⱥ�a� YL�?
�)���#��2��s�#�r3�4(�޸�6�*�＼��+jGtV��օ��}y������}Q]]_��r�q��p��Iń���{�$v}G��l
υjy���$��X���h�b?��F;�,���ΧL�y����0v�fO��;Cџe#4��_�[���O� ��=5�-�>X�v�"C��Q[�{dn�mN����?:ar���-���xUm~�aT^D��-�����F4�|��)���U�(�Y��t��ݷ��p
�
��h�M�풮�ǃqk��\���6�(�i�=E��}H�u�K��b�t7�7vwZ� 0�[P���;�H��R�����������#A4�#)�oŎ?(�
u���j(�I&Iʌ�|,�>>�ۤ�dHI��ٴ0��Vw!�SR�Z�mkZ�������k��X/qE�2�r!�y����vc�q%۴��M=���48�J -��x�B�z�^�� LdG�R0���)�Q�IMb��h�9��ES$*_]��ׄ�脚�5���^-�$* ��/�?+�4PKy��\�Yr�=t����?������(�"���fh�Q�w��)���n��1�`��5Yh��yH���o�o�Zֿ@�e�.���[e��d��}��r;��J(?�2[ȷJ�t����I6ԋ�`�����7���YT���r�s:׺+rRS"���ݨ������N5��Ӓ �_�4gX
�'Ұ�䃿��#��	;��&W���~y���w,�a��W2DQ�8�^ϣj?sy�Jm�?.}�x����H&N� ����U	��~���m<v�����Fr��$4�,�#�ћ��ު�4п^|o����Ӝ~�J�1�] j��22,,�?E��C�\�Xۡ�����
)�}	�"�}�N�0�Ƽ�Sr.����)M�dO�&?%�p隅!�M�=�]�:߆5L�hN#Z>Նg�T� ��:��$��}�5>.�?/=��%P�<6<tC��1��LAG��ә���'� w�9Wa��cg�6��&�Ap	��}��$s�~�+ag��偭v+V!��l*w�e�̲=�U�E����|������~k��}�C�!�N���<�+fW�Q���5mE^�ښ�s)���h��t�
�j̲��T�e-6�)����;������ ����VK�%Q�kFÓ�e��&R�y��n�R���`rypZ�͞#�H���