��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� ���4�p�M'k����Oeۮ����>�Z�:U+�ե �\ҽZ�f�7�� � �nG�bsD�6�4�k�N��+���¼x4>?$�T���e��m���5<P.̪��7L".�9�_��V�^<C�����+ ��UՃ�ƐF��}}���Ai�eߠ6F�հG���ҏ��4����jz�3䬽�s�ُ�ERr�0����!z�#1�;$��T��KcD>9�`
�x�ŧ��5ا���5j:�����������f��U 1���?̑ 5~����E�7�KE9-���=��.Gn���e�(Ċ^ȜT���0�� ����k���D�甖�vR�Z���̝5�,I$��&�&˾y_Qh�<J-2�DD(:�=X�=
:����	�sI
f|��.E�ef�d�{/!��Rq
q,����3�UL�jo�;�f��a��f[�\��V�z'($����Q�O�=�l�+��]���-�E6��`�j�.��#���a��z}v0��7��Q�{h7 pM�1)�qUr�D�z�����6b�aZq��N	��dy����zh
ݏi�4�
���G8x:6}jt�M-H�ڳ<c�}�xX5j�1:yM�?1����~�Y���d��BvXU�I?(V���/2���|=�?�+u�ȁ��K\{��]W93DG��
"Lv�+f�|Q	���NS�$�ml&�yq�p�YbL�m%@k����<��R�M�۽��xH��l�l-o�:�u���%������[���l�.���ԌLN ����]"����ϒ8m�N�_W��mp��svj[A�ӯ���l�%�}U��^0� ��@�U�"��2�'�80�`��־��BI�/�Ϫ��/��a`1�AE/Ͱ�����:G$�@C�=�N�{�Q��y��g�b�61F;��f_O
�GM`RX�i%��΃^'.Y��K���?x�:�8~�0�q��i皷\7z�[e8�RL>{�Ky���U~��a�EE�
�G���g&N��n��p31!P)��AK��
�ZJ_{�eg7x���i4���s�PJ��XPH�a��},���:��3d3\7�8��e­��U��Nkq��/ք��+�6x�K;�-��Ӏ�t���y�j��9�_��ejG\:�ȐJ��F;��W碸���bha:̜��(8s�M������l��l���W8�fN�'��j	RD-��>��vS�k�GGx�Z��P��?���n�39H@a�R�0��4�B�y�����p�	�A���E�mY��}��X��q�'w�VE��X��b+�r2D�򁛸I	嚨�g�G�D{:�gQ�3�K�Ȁ�GPm�D�(��qba���1���7�L��Ŕs��&
��,��9�U:][X����`-��l��3�������ma$�c��U���]�ˉqe7�u}}c: �~aSq}�%��Mز�߹��ԉj%$�o��X�Iy�`F����:a1�Zȓ6�$����~<|h��T������5��W��M���\h4fI糿Җ�N���j��,�KS���c{+�%Z0I-�%Q�vԽ'��P|��f� ��8@��b;�����#�����-t������>p���O'��zk��i�Qy�WΙׯ�G���e�S�nj�(��� ���J}v*9�+�G��Ø�˴͞�r]�=$1��l�Y7�u���>FG�A��s+���������T�2�~n��$&�Xf�� ��W�"I������ĹDuD_J���g@�������S�,F�,�N�J�f8��آ��t������S���s��:Ы���U"З�� ;~
;���dt���=Ye�-U�!����/�"��E���}sGKΗR]��F��Yj�b�S�L�e/@�\�e[Y���v�T��#��t���O&��ةYBB+���+KT�O�	J��+q����"%�zw�s�4~�����6�	��2����2��\&��ǹ\�9�>��O��(�v�����3�$����o��a�_��b�[�_S|Nq��._���e��.~v��K� F�1�Jͽ���0�Uה&y\�H{P=�=�^޾G-|NB�&�������{�C�qrv@g�����ݐa���5�IWB�i;k.�پJ��(�@C�����ٌ{
���\�UI�!2�- ��OR��BQ �C�u9ϘFR-�d�=��*�G ���/�h@��~���yj��Y��W���bq���s�EB���_���fMI��a�i����!� A[������F� UZ�&����T�������v�v��������.U��W��b�D{Ԗ"w������M`��$v�K�}��Y�4ɯX{W�7S�O=X}�P�)�#�ہ	�V6�5mȣPQ,�R,|�V�s���c��U��&�b7<N�l,#K����K�.9gǖ<N%�8K۶�N�e��Cxٍ�a��і��Vn�#!�� �E�k;/+�0ߎ��v�9b%�r�((�����h,�����&
%�}-<��+�mw�6