��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk������A�+��%������k��8V��)嚇o�����)����qSAr�0ɫ�NG2��ј���^2SӀwMW@�I���q&����R�q.-�g)Qǈ.c�7��^xC���*EY�@��e��EzAu�ttj�T&6li�Ke�_�U(#SQ=>�?�c)f�~W��R��He�^HB�xs�qd�ԛŲ��H�>� ��C�/�����-c툨����L�ƒ��ہSr�MQX�U-��x�%δhT��"�$	)�'"J�����n9�Qaa���LX_�Z�}u��ٖ�S�Dj6�$:X��7� 1 ��l��C�p�.�%z`o��ȐKX:�9��b՛�����6d��	%!�D�B�@f�49�u���?��a:�h�|�AS�'��i����Z�s���5�㆒k��!�at�k�;�V���?H�p��k��FB�ݰ�o�ڨ.e�� �h {}4�p�E���j"��T�y�r;Aa�(��)F�
4^�SE�W�7�����<RL̤ΜD��W���\���x�m�9$42/�Sh�>�$�T���C<b����2������I���l���\x��9&>���^S�TK(D~�K&�
����-;����_���6/-�`2�0Ξ~�r�e�H��v$ذ��@r�g���eg�\OU̅�N�X��a_����!M��\`?,Ml�^z̯�wG���i�:��2o�����N�1ى�<^�-w���}��A��*���zW�̎��q�N�#粪�!�>9���Yz��́���XCyY�Q9��29�B%��?D*�ǟɠ�����T8NZZz�ʇ#�j�0�ֺ����=]�����y�G�8x��`hSX�@L�,D��2m��m�ݎy��JJ�]G�Z\���֨�ͱ.�6��s�ˁ>:6-�n|i&�|�����$��{��?�BwB*��N�u)�%E���j[gDM�>S���Z�/�QhPt�Q`�DV&Gh���r��W��GU
bJor�>>Ǧ/���I��^���H�=i9��߀��8B/��􅩷H�cK�XyEC*�����em.��^��5 ��e<�~�|z��Y/ O�~H8 ?��ē�㨂�b]"��L��b��-�W���2%|
E�y<㖉7�;c��<�N��"S^����zv���`&�����Ď,�d����5{8�6�7�Sm�۬G��� J��� �B�W���@ "!�hU:m�x�#K���P��SW�| 7X�jk�N��7��Qu�W�j��nBj�c��X��0��]��L������.m)Y!8>5"z#���07��r�2�S�t�2.�}X$=��ï�[��G���kBgD/�Kq=��)ߧg�e~w��xT���k4l�d�҅�{��aRQ�*j0>Z+����������_+o.�j�҈b]�o7�B�v�?ɤ'wس���H��H�X'��7�UL�cڟ�c�7y����$�-�n}���!@j�%J�.�$���+������j$?v���ș/����-��@
:H?�g��e"\=mU^Ηn#|a��@#�`k��̃x���Ô8�~	p���}L���ʻ=�hd�+IG��\!ګU��7vÝF� ܴ�ĒX��BMN�r5��C��yVɥ�2#(�3띠z�2N�_G��P3q�4FI5�[�.p�Tr���c�VwP�{["	J�p��X���j�7n�Z3)�j���z�}��=�H�C��o6(vA��->�[�.�g�V�n�M<���>���l��n���F]D7(S1UA���s4��$ȉ��z�1�֥�.�E�x�/9����������@m4T[�+�9.��Tݓ�BB�DA�����ԏ,�`UV���ƻ��������Q�sg���Q���_�MlƓ)���/��i2��w�;a��R4IJ.مK��fqH;�'�j`��a���mwO�rAq75�wA���gSj�{�Ij��B<C�� ��!X�O��"F���9sjđ���~�_0�b���ݹ4."f���3m]$b3:3At½3q�7�w34�Mq���h��*1�E���b{�2Ux6U�geP�ǻ��w�ڥ1,Ǉ9�;d�~�?h�U@0��(!	���w$.���;�S ���,ljӦ��Y����t���?��I�q�X��� fT~�*p ��!��+B`�5n�8"�#�����;O��Y������R]Q�ێ���mr¹S�� f��g��Y ���4�۶jr�,���*�&�%��^��ez�՟%L�4� R���a`e�q.��
 ܫ#�`yU�#cx 3�}�%���%0ԲE
���0_78!�1�꒜��a8-Xe��#;'z�B�Q7�fZ'� �-E�v�8����T@��O���zn����\��K�u�������[m������q�$=-�O�f��ۆ�
B��6���4� )#ȝ����*'oYf:� "�8};eN)�3.�g��4�y��jxG�:�G�X$��u��2�  G�������}ڈ�ňB����P�Ae�r�z��@��U����Uoh<���
Px�ZkI�)����I��rw|)8�W�4����^K���YƗ��6�9Uu�N,EAAT]{�z��jw�ӓ��usӥ$�"ސH]�U�JV~�e��N`�Cԟ�;�ڈ;9r��7K�� []?)�֒.�9fgĴ[���cmy��	���؆� ���� ́�w���v�l�<A�?x�Ä�yסA:3e	a��I�Q�\G��D7���/�;���(�fpY���uq:oEH��"���Lp���������w�B�AS��R��TO�!$0jf�1]����#:��e��8�sNF� ������:^��y-�,�����%�A���0u '��2q�cP�����E�~��L��P%9?��o:�qdv��
�D��0�/W�5w�~N�VBz�:��۝YqP���Md<���{�}�v5B�+x%=YK�V?��~-ǲD9�[ ,�r����-���{-��M$�AN!k!���6;�6L-R� Y���2�ID͏�eVj�=ϻ�~�OZeF]�P$��Q�)�����9��`�?��j<���ǋ�OILN�ԁ㱓� ���"�b�2��B6�y�!�����ΐq���7nEkya*�g�~���Α'�a����Ys�dv��$�3���\TV|]2�Ѵ���	Щ��]�R���L�gl*+�j�@ƚ���qKy�/\G�&�*����H��kYT��4H��c��yr�3�K�D*93�zJ�x�����H�aT���k]�b�B��q�_�&ٕ���8�K��.�LE�ם�`Ǫztkyl�o&y��A�D������畔O��g���n�G2�ާ#�i#Ɯ�<����}��\�����?2[�Ԗ��,��i#K8�i�ۧ工���uqp����}mn�\C
x����Ɖa!�,/�G�K�T���73h����0��}�� �b��#���ň*�{�<LC��r������4�}��YÙ��I��㽒��'�u�B��������K�lhCxRӍ���S1Xh�gWT����Ġ�#�X����	�=b�kG�D:�/&v�K��Ƀh=z�ö�#� b�\���mU���G�s����?V�h~p�x�-���ot��t4F�Mԅ^CmNi�B�7�?�u�́w����I�\��!q�e+~���y�R' �`;�k��-�w3�Vr,-k��b��}?�ddܨ�2�qas���	��?�Q؇��j�"f��3"�y�=���z/[j��O���OB�c��Rd@�uEk�TId�_Ჸ�I����JD
������M�����	<.�H�,&��M9aI^)QR�;�hhN�jU�al��������F����J��O�k�wJ汣&ț��oֳ�ܶI��}�a��2m��g<f�]��b���D��tȢ���wGZ��H�	s�&���=����ֳ�9�PD��G���`�Ȫب�]����ic�$r������H`��'j ���P	C�ke��vL_�Y��O�LvII�Y��i˞ĶS�P�<�*�9~;��_����p����Μq�K���R��{�ȉro7<����ꖕ�K�h���/c����<Lz-�j=����a6'WU���3�*�W�	�%����@��1X�셀UG�=���~-'jqxU;+����s.���d#a�~��n����GS�50%���-ozh���vAD�^f!D>a�Ҿٙ_��m����	4��k���^ҋ:�ڶ2hN�[��I�����1|m۝K�P�
ou�n�����^?��y��0�Sy�L4$	���Q�$C���Ixx��C�$�٪�()eHG"���[�Y��$n[\9eM�V^�^Z�_%�W�f�x��2E�_X�S�z��ʀ�� �ݷTȹSY��������C����=���,���z��q�6��SW��cƙ0�OQ�@µ���2���KQ��s�l�L�1u�!��$e<=f��	m�����J�W٭CF�C$Uq��� #Ӵo[z�
(�L�*��N�$^�=��N���8ESX�H`/O\e�6��x�8��}S1���{v���	��^C#���MR�d � H�Q&Nݒ��eb��[��g)���*5�M\C1��R�ies<��V˿I�#��kN�{�+{._UB��?�N�,�T��D��Ġ`l��\�wSS*�=�-e(��)�-��8��R�����e^*{����f�mB�	FoNr�Y�T��_�t7�(z�K �O��2��F��;�]�1r�����> C�f�&抻1�)
\[Î$���K�,YK7�����&��,�W�h]Í�X��z�Dq����H��f��k�Li>b�:8ew"��=y�`ɡ���L��h�?d�'��a��H�u�߲!�������R��pw�*��RYqW��Qu;�	3��-�
ĺ4bmm���ra��ųi2H,�Yr�� ��!F6��[�8��'wP�
F�֊������l�Ə��Y�H/D�Kǖi4i�;�U��t�'���NP:�Z?9�d�
�!+u�����:�ݩ�����U�Iە|-�5���<K(�:I��2�`�>�L�g��ݢ��綊�%i��a���P���M��#��N{.������� sm��~l$�I�z8uK��R� k0ˌ?=2@�}�=�x�gӍ&؎�1F�]�� ڈlq�X��p��R�>Sg��\2���:O�3�[���8�sҼ�!˃�4IM%lf�����W*�
��"����ê-�.��ۯ;�sW�0{���#l3�P"`�O�]c�Fz4�ʆ/m�@"1� ��'cގ���Y���N&����/��7�N��	�i��Ӱ@��l9�>���[�J��h1�)�����S=�:~|׍�k�*(h�h.4�3�{����!���ʲ�"�_�<F���&�'"�n}ۼG)[K�Cў^i�4���P�g	���ň���W7[�y��U�֞f�l�K�����%���d�0�c�����к`�����@��.��W\ܕ�c ik�����n���7v��{������r�P�B�<(��N���	��0���)ݨ��+i�[�<�c��Lח�C�t^J�m���'i�^�4)8�����r��aLz0���E�i�S~ϫ	ܙL�Um\�m�'��kRl�bCߔ/��q�O�x/���0�]I0+�������7���)C��K��ׄ��`�5Z-�g]r#���t~�w�ʔJ��V�}ڀf!Vd�����r{K�Cxǃ��r�t'ԜL$�.��C��Ry�_����.Z�q	p��G���+��S��M7�0�$_G/�m?_ۗf��6.5��0g�"�rj�kCh�#��E#p�� yC�Qج�&8��[v*�MVI�Ɣ�H4m���TQ���6����|= �ݾf��Ģ��T���蝋Kkމ*�0f��̊������9'?�
js�V?��=�*�?d]P�H�?���xeV�][�޴����1�z���A�mv�D'ȉCV���6/g�F���*:�A�t�N(�x��K�Q��ؑ��y�)-�����[�B.oz\��/SVk���6z���_�!��������'�ۜN�'T�����,'����E�u��ʋO8�Fp��?����F�B�n���uS>X�2Mͩ�Z̛��}� Q�W�3��%pԬ;|�$Z���^���g��a����|�������ݦ ���gI:�g����Tǭ��w�ᆽ�X"Y����\r�6�4�Ī�� @�.[1,���q�����
��
K0��2�A<#ؿ@.�H{���5ߠ�I$nf�����Aq�.��_܉��(��h�A�K�b��Aס�8�罩��.M�6N�SD����7�\�+�sS�[T�� ���\J�����@kC+��W����Q�t�Y�lY��E[��h��xeu^��1"��a���ob��:�����a��K.��x��4�	o�~���/�G�3��g)���TD�Z�xˍ|9�r�`��%�q?vP�U0Q��m��, �x�S(A�<l�#�n��M�]]�A|��C�霘�y�}x*wϷ�g1~1N���m�Xk
~�P*eB��l�筰����J�.���6o���.,�0�]�� �/\4R	T%�1o<(%��Zh!9����kN��4���@����o�,e�NZ��x�|i��xŎ��v3RuW�<�-.���~Ll����C&�v)m�Xt#iSP��F�F��!v�H�!�`(Ӝ,��]b��_ؠ�&�!h)<��"��kwN�v�?*�|�r�w1�½�� X�܇�>�UV�f�W�cd;E�\(�VvXej�bz�R#���v�4I�O�����:h��N��u��ۆڃ�ޔWuFn�PF)>J�e�R赘!�I8����8;�?��_��.;��"^��2[}-��qo�keg16faTQ��C-�X$F�fIY\�qq�uN7�6s�:ꤷR�Z�sd���p�Q�H&'�c6B}��om���(�։J^D�Ԍ�<���:>�\�Z��4�r �Oϫ��N���X?}#�U|$3���`��AXu�|�Ě�r��B�p�7�!�2��s{���.iq��{��O�:I���Mc�ϙJ�}����ܸ�]���L����\҅f�'�KK��4���L��0���3�(��pP�p����C�����+V��,�x�^�W����|o�҄��U��T�B�K�z��jP�.�Ͳ`�����
x�HH-ZG��B�ٸxXl�no��<�T=wk8��s�u�H?�~�X\�?Sy#4TП4츕9�;{P�c$B�e��삑|lP��A��u=
�Z��kla@ҳ���^C�X��7�_$bء&&˝��hҭL�#|�c( ��x�0����|h)�t܏�9!���\�թHC
W�N�O6a�Y����� �G�Az?AP� ,�Ǿ�g)�I"���򚙬at��b��>�����.,Sw2�V�����>��&5��1 �E�~�]\c˧���~J���i�a�#�������5�}�"�0G��M]�p*:��?�`�r�6��Db/���x�q��%
��n����[H!������W�㪰�p
���+���z�}��N���N�V�G��\�Łt��U�q�z�a�ƁYK۵"^!��_(��O�H7���Jڷ`t�7S(�d��ň��`V�{%�Bx,Ǿ���Z^���K��Q�;TRZ��6nz^,oW�l7���a�A=ϸ%��í�X��9���-j� gl�b7��~\�1���rG/�\�Zٯt��C)R�Q�{� � ���l܈�EJ2H�@A�	�%6� b�f�ض�F��y�����I^~�[�Z]g��k�$k�
�ǖ��i]�>�Hz�!�'��DM�߸��l�~����'~��!]~����Г��@c�M�əOF�Ồ�8i��UYmիl�ɰnG��{�Am�����f�q���P��	��g���fR9E�,��^�ӄ��R)��`��v"� *�q����=Z���;]��j�2�'��c��E�I�|�����t��p�U�Q��1R�s=53���3'�qOJ�ՎE��"��M$`7n���g���$"*s�ׂ�X��������-�U���e�52У�rRfE��}���$���8��b)��rOgc_=�o-'�H!�t���U�Ubܔ3	B2�LJM���F4�t;��l|fF��s��{j%٥}��M޷��i�@�+�l��E�Jh�`G �`��zǢɠ	�7V�~���_�>�s^V����.�2o 3�։��1H��zx�/*K������OA��%U`����L�_�Q���NTH^S�f���h�K뙛ۭ���҈�&�z)S&��52��K�܏�	4���#���=�ÿ�EC �h�aҶ�~�����_��7��a?�K�%+�y���B<����[`P�[,/,_�pLKlq�!�T|�X+�X����Z7�!Ў"rlܱ���M�H4sD���cIP	?T�;���$7�X�cwG�A>Z Q�Tg��fv?77H<��D�(>��`f^�id�#X`��h�+�*�������0�(��s:�]��nNP���*,HSB�E��wiW�W�ŪI�N�L|�f��u���#.�fO����X5�=�1p�  v�Td�H�fmb�HjL�m}ۦ4.�ŇuG��?"�1�pz�:��;�X����O N�x���81�z%�n�7��ߍ��AD�#�o�xM>��Y�����>�wcj��X%u��{*v�(�����eٶ�"dm_L�R@b�b ܱ��y+��Et����o�ƄQ��U)��]�����	/_�j�#����g_U���p��}cHn���o��]�l.a��������R��B���\���"tYl<�תVՕ�3WBw��e��x֮y��]��o����]� �o�f�}�'T.u8�����TT��ϰ��HU���� ����OV<�i�-=��`�<�b<t�S6W7$�,#׼}���M��zp.vęKX$��"g��>����t�b̟['2�!{��ԩ,*���I̚����$��V@�:�o���{ITNfXL��[f��Вr~�5|�'o�am0�.��X�ysj�yo�m��暽bka���/�?	��� ����_�>��'o���/��<2*H����-{��]j���jA�kR��K&���Z��f��<}���%#p�԰W|ߓ���e�BNph`f�Ef��x&@��t�M�+;��q�X^-Ҳ�&�n�x����?rG���qz8�&�x�hS%3.��|�Lw]d��v�r��)�
b��$�m0�	��xT�ͤ����~B$��Ä"���\1�9J"�el�r�Y�ށdxg�P��x�l�p�~�U �Dm��`�Q�3�11,R�Jr�&����اE�+ù�]�OVE�Ky-�f*�jd����5�+F=A2з��c;�k_Nϼ)�ea�j���"C%�em���~�*?z+�7�(Pz�Kw.��tX6����R�^ 2qb�TH�N꣚��*��d����vL}��Y��(��x����
[�%����2�0_���*���X����r�/���+Ip�v}}�'�U�X��Q`���+#Ҡ��$��:��Wg�8�������5_��7.� x��|�~�G�h6e=�&y�=͟���zy�U���;F�cr�Q�T���� �rs��-ɝ�1lF����0	����D^�tHƅ!9!�����~T�88�h�/�>s�H����P��a�y�j�H��A�aȡ�~H�_k�r|��_����Y��%U��,������TN23R��[���0Z������k�>a���HqI#O��[�l��CJ�͇�?� [2����~(��Yt
l��F� ��~��`NjT\�u?��:���������c�?,����n�% 4�x��mY�[�v�T�q@�þ0�{���Ts��*����>]f�ǋ��R|���!����\���0dNΑ|{;�|�>~��R?��)���i��K��\�s�Q����W�����|�0\�W�.�M�a#�@>iϷ��ī�ik��/�6�2F�5�>�i!���,!�Q���D�=���<���גej�>�3_��=-�������W?�f�2��V����.i�66c�4� d�Tj���=Dˌ�}�Vꃳ>�кm&?t��0��.�� ��2�V�m G�����8�B��r�w]��<P_݃xY�����$
?@���� ���m�� �A��ļ��JK���� ��5׶|$Ǻ�4�Z
�&`����{��I��Y&�����rV�(ZP�T��-_��s�6Ӱ��Ϛ�F1g�grem1�ʚ��\����#,Vc;�J�V5V�T6N�G�tā�HF���S{7w��wǑ�Y����G(��:��A�Ŭ���Ak]��Ꙥˑ��A����(5�~F�·Q5%cZ��I��!����p�f!�r��������U�}p�X�������f�uI���):%�-i*zb�_�����G/|(��-)y���(���v�W��,��? �	�3��n�jT��9y9���8���	vS���YG�l��mz�R`��k�~�jث�G������o١����I	�7�J�\�`����E�ϵ���#%Q���Y�aE�i�pvt�H�v���ܺMP�̅��O�n�W��D�`V-��R�3����>��!�JgG���Is��"A�Dr��Yҵ��`�h[�|�#��ɔH��N�"���/!���^�Y��a�ZJt��
[.�"��Zccg���ߣ(�	�K���ڏ���J]�f�����ȵ­;Ĵ�g^^������(ҝmWu���}<�נe��"=�e�96J���}_���^�5AU)Aì�{Y�0�{����G
�o���U�=�&
���^�I!jF�9<�r)��ĝ7Կ��6,�)�{K�@A�W�!�;��5r)N��v�[�T�,w.8WW���D�e�/�{�"Q��_u3R�����H�죝`Ct��slD��u/J&�X�g4�cY�G�]/��K3���n��=�.��m3���#��*�zj��ؿ���L�.
��������eX�@b�TO�Xy�?�93ێCn��TO-ūy;S�^R�!����D (]�\x���(-s���r_f��JC	�ɖ�R���&[N��V!d���+wj/���24��rY�&�~$��1�~3,䋵P�ь�%'�s��*'��og�ŢFh��mE�Д�W>�r=�������xj�����a&bL�0�F���W��3�#��R'NǠ�k� \^h9pv�o��������z_��Ⴘ�Ԑؖ}� x[�<ۄV&iHad�5|i?����l�:��+�Ȋ̻����q�o$����]9�e��R�U��|:�<�@d7 (�w	寤��-甋WD�6T��t;T*��N��Bu�)��o�@���B�������c�����k���%~�*�J�u fԀYt����__�7I�X*!$�aϹ�W�nr�[�(:��H*>E�in���F>�Їv�����ғ[s^M�ђ^c����⸹�)b</2Q��X:�~���?���&tA���϶�ac`�8K>C�s� 0���
ÿZ'y�&��jp��M�6�����)o���
w,w�����u�w�����
oX�.�d{��������Fh���n��\����/��p/���6��c%��'Z�
�54y�|��j���{d5��$u�kfWT��5�9r�o;�T�#%��(���EƐ� \Y��t}�CRw4��:&�$��o���ɔ������\����d���-f pNǜ��d�Yn�ǑJ~����(:�b*Rx��%�B��P��XO��:��5��z����݇סsU�ړۺ����PM����e(�y�1�C�t;1;�s��{)Ճ�rS���������������\��(	&�u3��|��� ��]�UU�c����1��nEǝ��}"V�e�s��\Ơ(�aӤ�@I�2,�~���N3i[9+h�����G^)��?����آ1K5&�qi�U�04[�d
M�ԃU��#�=b�e0��C��O�1��a�#�'<�p�P����� ��;`p���#P����J8�H<��1$�a�w������n������5ʩIn �h7���C��΢�\8�I���*&���/%��*���μ��pĂD���Y��g���oV\�+�=:�{q�gM��%#�]��b�p+6�����3ؠ����s��2(�K1*�d��gm�6^4I���J���nQ�P2���V5�� ����J !��m0(i���K�X�Ɉ2��(�ln�eJ���x�����hҴs�!Ğ�� I]n�{��-
�^^,��' X�m�ҫ�$�J5��\� �=wb�@�h��m�qc�Jm%ڕ�k��8u`a_~{��	 �Vt؏>B�ކa��������yD�����6"�iX��<	V8r�!�/��L&��6�.�9��7��$��N%N�o�f���ϫT�Hu�W�ZY����� ��6I�PŤKSrpɤ`+r�!M� ��I`�'�oں����A��i���4[HF����sZbo����> �
.n��1��R�:��נ��6���#l��4����ua��X��\?�=z�bb�$��5��?ғk��� +��`)s9�|����Uzj�z�m�̷~w���#��-u�Po��/zIrp�(ۻ�2X&8��]�(�E�H�k�ױONG؁�����25�_H镥
a�W��=��T�|��L��Ո";����n ��&֤�'-�~5K?��^�D1�F��̏W,Դ�h�6.d�2������R��&���3A��{T�oOɘ�X�K�`)��i_*�>�q{?�I�m�dcӶ���0��u��]R���0�L�s��DTv?s��X��6K"���!&9��K�6*N�\�4Z%+,���(����N���g�����u	�l٩zR���X�����H�m	�m|�״�3�Y�V祒���ϥY��-�1>}f� [HA�Vط�#ǡ%d�Ҕ䫦����7/>��(�,��?��դ0�Dq�7Q%��,1`R�L�dN>vmG:�4����7�F9,]����H���+�(�Y�H�!�e��@����`�֤v�dSB��S���'7���ox�w���$�dǢƛg�����]uڀ�ɥ�9���&_/��e���]�n1s\�1�㦰��Y[��f���+G��łQcb�j��gYWS�c��lIu����BOX�'�1��x2���J}�/��\|�)u�SC]�A)9���}��b�Yc� �b�4��$��:����h����Ǫ�fn�m=�%CAq�NC�I�8f�oUf;ϊ���o�pvp�)�dy��Qa�ܑ{�0Ej@(t�����ɣ��j+���V��H��y	[H�R"�x�hl�g��1d�K+�a:��HN*K0��Ra?y�R@�u]4K�ބ��Q���Q06�/�9jQ65��9���Xb��.��n�UH��K�>�'���dڿHc�+@Μ�v��$��:+v�*�|��[~
�����q�v�U�(�.ZYlm)U}�d���g��� ��&�7?�W�ʄ�h��礽%)�b��|U~�Q�g��1������N�tg��� ���K飔,�cE��o*�e��3z�5�9����ݔ�}te�V�Joc�k,O��}4����Xu)�/�3��a� 4�.��pM��u�7]�^��zB#�T��1a9��_/V�V듬#��*#>��=�X���3� ���/ee�����?.m9%����������8e��`8���h��Ѥ�)+��C��P���^S�d�,�l�E+867w��o^�qm;Td��\[&��H��ԑ�����|�>���!�\^��LA�LK��0&��nI�P�T�0�I�B��^��r�6� 2���19���Fn�#4�*��ECl܂9�)���(suEJqɲ!EݚT��8w�؂<�[x�_����x�q�Z��>���������2I������	�����Yª�f}R)�	��������0�^�ɢ���<���Ё�2�uuD7-�j��Ǆ�`�g��}���x�RowjfZnRѤ3N�Ql˓�#�ҝ���e��C��\.�j}���5���S[+�$�b����`�,���0�V��{8!7yӚ�S�󨙊�g���n��c:U��u���b��! ��̞<Hc��^/H��*���ߪv|r�p������{do�-����g��M�I@�ie Ս��Σ�ȋx�Zct��!@�@T�Qr��Ī�j��s�M��%e��fԞ�[�]%B~�����]
5�H%���(���57��#u̢�8C����,���� �}'i`6�=�A�0�|3��$6���p��a�<���J�=����Er�/��Þ�<������������Wsˠ���:�~�Xz���o@eL���A������Jo����c�؉� ��[��ݚ���*$d��¨�[�y�l"��
�"��U#�L���K�W��8�Īa�b6Bt��?ϛHU����Ԓ��P/���ҲE�-���jD�ҕ Ebŀ<�D�� 	p�1j���Ε�z������}�U7�x;Z���1��pR�*ہ�Y&οS`��С�!M4�>%OrlV��jH���}� m��λ��\��a��Ѕ.�҅/�c^��!)K��$���4��r�[%	1�	�N|w��끙��!��׭�+=��,|�&T�>Z��I�3K�<�c`g�?r&�*a∖LcE��ש�~[��Y�o�2�m�5�G�d�2��Ε��q�n�8���;��K��M�N�0�Ȭ�*J�u~�Um��@9A%�^Q�cwCV�?�"����s���1�v�ֈ!:��y;�@���}l����ȹp,�2���k���,��"4INnig-����2q�N��N��6��e9Gk�C3�g���-�(չ~��W	Vb<����|�C��@�>��;g��x���+HV^��μZ3`	m�z��O�H�>>��@��x1᏶bT�0����<NM%��I��@/"��6TNIrz�W�|)#����gf+��J(�-[�_*U���X�ӿ�^�U��5��H(4���i:oжm���)��1����0�����Nʿ��Y�ra�߄���F~5��
�1b}�$��C�`x_yQ������lA��_.���_�
�w�&�Vat`�Tb�okH)=|�c�(�P��C�p�W,V�~4�کi7J~A\��$cz�Vj��X�� �GH�	�����f��4���o�"tws���S�vs+�8G<9[4v�s�U��X�n��*��n*�<Nu �V��A��:9�d��Z�n�H�i���@��	Ә\Ν���ԁC{��=��\���T ]t�#������x_0�U����u��ڊ}�a��1HEnR��p��'y�����S��|�Jkm��O��k^���t��q\CzDTp���Jy�bp��U&!�4ey4��%����"���,��@!3�s���P-�5�\l�� /�n�"�4��^��7�r����bkq��I����U��y)�4��#�q��_���F�Sx$v���P�-/��
0l�����t�d�*Y�ɧ`'yFڏ0�I���Y���Τ�����:�g'����.�eݎ^s�^��nQ��T7sʘ/[O-��('�W��jgw��[�Ȑ�d�g�L�J��Jr�o�R	v��%L�w:^U=���{0�?�H.7��!+ѷ��Y��Ll�[>c�4�Q!��������zQ�'��ݳ�ǅ��&cV�[��vo�lGp{n�ː�ܦ�V�;w�uHi�#�IQ������۴��D��El�p���se��Wa-u���]���|�@�L��A㍐9�;�(�����4օW�j�2jbH�z@�ҽ�I��g����GB-�|��F$?�D�+�Qv���O�V~P��W�V3����~���w���y� ��w߽��0���.����u� 7�+e�ق�.0����t�4���e+L�UQ����tz8���^�!���x���U�mGf�X���=�u��ᘝ�=u��0��t���m&��<�[�;�N;5}�&���1��\���i���
�N�i"�}@+�GsBbJ':5@�;��0������͆鏎�(2�m��7������No�_F���E���@	�I�h�P#���q%����ޏ��2�/x��Ws�3:q�oF����L�{=Lr�1j���f�'h]�%����\�JZ<y���f��iQ�F�NHo���)-K<�ޞ�$?��ħ�~v�S��H/^�a�籶��V��R�
6y,��������n��d��匱9C_��j5��u��.����_<��L��U� �F4˱�8t�o�L��y��SI���U�τ��K�5k��$Z~p��4������^S�᭗�>.�2	�0n��H^�ܣ�!��i0�����se���>�8�Ǵk����_�k��~�8x���u�F�~h�R��$6Joŧ�n�M�Yr��)��-���Z~�&E��Ҟ��7��P�H�����������/��zx��9�v��>�^���'�����BNR"�21Ն�{v��\���10���2��������S��-R���ѿ�|�ԇH�5��a�(s���K8fg�!��	p[*�Ʊ[�͊.:|X(�,��Da�R�?_���L���s�o
�w��#�h�^\*����P�@C*��yQ�7���$���^%�no)��ePJ��!�;?�ۙc�龐�I�ou�`�Y�~a`1G=)+�w���|=ۮ��9�ɤ�U�lB�sbr	`DS��S8ĉ�UV0AxN�V���AY�ԂtUN�ls04��n���;���Fhm�U���0�j��:��F�?�	���b����}k�gI����q.-���p��������U���@�n��x�C<�:IO�;�?2B�X��D�@bMM����P	b��ۚ���������H�Ҋ�+6�6��n�[��&�nM)�Z!��ҟB�=�4|�'vb�����I~�;�v��k�je!��"'{�9�&�幅8��[������L�?��~7�%��X��T>�;�k�sl��X*�����c��Y9��wO�9�pX2�b��R���8z�A�8�Ă���S`!�<��Yܬ����Z��ݧ]P�`�9���{��)�8�sDǷXW������q��8�����|���ی���u3������ȣ����5����gJ������
AƆ�U7�b�܏cr���`��S�qp��Ͽ��d�m�0��R�^>�&O�Kd�.~�~�z[FS���]���\�8�ۢ����4�6���{�Q>E2��
�����e�)����w�Y��f��\�1�L�2ˇA�$[�f��u!_�:d]FG�Ө�$��a���W�GJ񶪅�ؑZ��'Q��N*(6]�=�vs��1!N��-U��.�N���W"@���CG��X�p P瑚��d��;�.f�c�Z�"cY��w�C�J���J3���O��U7�$�e�=~\J�x�"���"9� ?�,��v(� ��eݰ`�RB�]A�Il����6|�r߱��6�q���ȾWb�^�.98;ʉ�H��Xư>R �".iR�w���2�3M�p��jlʆ��)B�� �z��,�������kQR�E���O��<�4���DJ��AN�"c
��mY�c�g����v y�*���*�ݝ���R�N<�oG�[Q��/ڨ���@ۢ�Bv�N�)�����t5�n�H#��`�
��M/�}E��(�q@�[!����r�Ta	Va��0��P`���҉� �ї[�k�gc�|�&�:�Ư4�}fX7�E�����a�]��=CK-�0�]�p�(ū��Ù@S�f$�Tr*dB����1q�͵���)O	��4k`��
 e�f`�C��֪D%q\ѫ!�9u
��r�D<1'ɓt�U�I�7��`�V��$zA�ު���B۳���t)<������c3��g'��A���B6��U��dO'�S�HWJ�+&�����ˢ�ن�޸��q co�lJOF��k��mRz`h\]8,���z�8f�=8J@�Ԧe%6�C"�Gs%�M�$7�8^P��G;���i3���p�w�L�x�&S�����"�'��;,oU�΍�xU�`�`�A4�ƌo2>���_^�3��a���q:����ua��+�=�W�EQJ��"��[���m�a��:{%f������o��j�����)	�m\z{�{T