��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ����u�SM{�[g�hⰱz���dLm +%&S!�ߟW&Cao�&�����U4���������ƭ��M��ֻ:V(���.��(�~�`�v���d0Xr��c����r̰!��Q�LK#�qZ�:yT��"J�1������j��&�d�0c��9#��0��_�Ɔ#����C����ގF�uKz��U��R8̒��F��-�:+.�N���y}`a������n�W���ؘ��ݔ�.9Ƀ��ڪzo;��+X7'�ob���;�kbYH���*���Re�^����G����9_^�����o'�e�*�W���>Ќ�w;��������@����0��'jr���WpvÂ�x/.$I����X!��5MӒ��U���I��e���V75���7���L��eH�+�X7�`*�.���K58�����T �(Jo�
��d���\�4�~�ۮۤ��� @����JQgD�V,=MzJQ¥����)�����e8��% v�]T�������lF��L9���M�'���T�����W+ޥ���M��	i��zI�wϮi�z[$W�Y��=���zJ��6V8w�dm�&��E����E�jȻV�2	w��Jq�.�сԶ�hl|D0���^
�[uR�܆����s;#\2�| �Ǉ�ro��Y�����4�x���S0�GF��	&���\C�J�G���"�C~�#L���\�Z�j�,���X �%9=>źT�0@���Q�"�*���/�H˩�m=HR '���&���ʉ+�51lp���wf}T�v�v���W�����w���hrq�+pm\�k��摎F�K��O���&T� 6��V!��l(P��ݛ�.Z����u���v�&����$�s���q�
��=d|��I���d'-�)�z��f��'k�S̤�h�A�I&�n��l�(�8��|X�L�����# s�uV���qM.� ��.cy]���<"�����2e�)�����ckF�1���0�����&����2LH�����Z#��r��g�x@3�����]��%�+�)�k����N%����8$�`���,��"���dM���8y8����f���|�>�C��o� 5w�w�d^'�G��4�=r?���?+w��S�V,��bg�-xf�>�>�O�%�Xh���a���b���ukZ����̒�U����zLF������Y�Ǿ�h uNڙ��2с��M\YY�)x�(���<����<s�R�OV�C{�}ϝ�K"�H���%p��9��K<gEWy�Gy�E��t�J���Xv��9�*<u��β�W!�¨P����d������L��:������Y��p���7�k�:i
}I�ċE�[\���M�Y��܃�"�
0rЅ�ԋJCe�|�o���8���?a픭"xV �,-R�$t]" ��JS}��$h<cY8�g��W�p��>5��6UB�d����p��%�ȩ&}q�m0�
��D"�Q����M�/)S�&�w�
Y_Ւ��>�Y�6��,g�"�Hw#qё�_h�2萌��ݞN80�2�����X{�s��M�E�+�neqc_L���smZ^C&>|5�lm@2��|�6�4k����@�*�~�ǘ�HD�.��"Gt_�ko��j6�x��Q�$:.~a�z����1>K"�6���)�~G]J ��)Qٓ8F�5��k�x@g7+ʉ��D�b���*qs�|��?��k�5���	���aM!W�Z~W�X�3��}�V=�j��3�mK�݌Z�V��*��ༀH�)����@#��%sIj���y�C4����e�l�OHmo�և��y��&��� �A���: �Jͅz��*�0!��R��9n��L����\U)>�\3�CI0`�(��Һ3���_�ٛ�����4������j㴨�U[
X����`2k-_<�����"��N���]��h0�#5�n�����%4��׈R<I��/g9�f��J��S,A��|��9��)�#�p8�ɾf���蔕0_�iqu���i�:G���ڮ��dq��������v�OW��:���;+<洺݅��yJ��m��ƍ��+��q9���ax�4���{��.^^�K���
c7�݆:Yܮ�AF���suZ�4q
Ssbng>qT҄�p�Z�/͸������:��&�,�����ѴX�����x2����!��E?0�<.��=U3����]tf^\�����l�s߹�+�1�u^����.=A>�wv����y�˔r|� �=��;Nw1���9JH@2�p5j[�pTt�}6�W0C�l���iџ Y]�1v��;��?�`��k�ۊz��
J����8���r�p�ө�Us��vI�z8�	�a��%�I+��3D���#����;~Ϯ�B[�t��Q�@3ۅ�~���#1�%�Z.����Riz�cX���Ȥ�e�rL`ص�<�.� ��	H[��x)�&����r�9~�L�9���+�(	Bg�/�F	`��S:��q�ݦ*�{�e_�ȌJ��uM< YW�,��=:�Z�A��N����D��)2�����ܠi!m���y��|C�A���!��<���Hl2��:��v��0)�&�!𣚱;�72���L�3�YeC�����u��FI���xbr!��ѭZz��-�����=u?�pS�B�|�2e٬�,�&�N�ľCDT�Ê0����9�z�ǅ��co�/��ӈ�;+��"Y��+rˣ*d@�jF�>������O���0.�C͝w!in���rC�y讨o ��(�c�a1��`��5AX4�*�<b�Z��!���
p�V�}���.��p8���W?�K��o	
Ԇd��jcm�pwO���"��������O����T�n��\���]#0�+�2
�K�\���2K��%���j�Yk�1���m���m��3'���A��kd��$�XB�8��U��	U?��|8��w�4@M^ݰ�8Xy�,���$͡�`�%�l��O/� �C�,�QCz L��$��ܵe�ƷCX.�LNu��8���N=H��X�ut� �9P�M���ۑBc�,��������D{���t�q�8 �M��f�8�z��m��AD��紜����н&��sg���:Z���|<~O:o�
H0")�4�M��:�b�N҂s\�R[��Qj��Ϣ�x�`.
���z��)C �O�	pK��_M0%���-x�F��i�T��y�\vL)Z����o�},/p������*t6]�R��;���j1\�ܲ�\�D��T^~����`�y��2�&���Oq).g�,B��j|ʉFO ����,���s]�Lژ#
e��o�uA/c/����$dYn��bO>[�|�2{��TE�E���S�ru�uQ�ۺ��GF.���|���j����-��0(�G�8r$�^l�
e"g�
7�a��j9�淵N�a�>U�~�FjId�In'�3<ߡ-q�j�$�s�r�\��wC�X��] ��\	�|��i�ф��6gc��YE\r�RuoV�ݞ雧w}3M��y����o�I��������Z<��3P.�P2PR�Y��pףgz����dA�[�i�1{��&���<��B�P`����U��\��A�%�80��>ȩXֆ�#�����8�6��)^ˑs�K%z����_��&|*ip���-��b۠'J1�7����k 2?���mt������M�{S�\_�`��0�2>���~h�yE��@���f�/�۴�ϼ�\F�e�d�!�η*s�b�����b+K���.��kQV��+D7,�	/��t�U;g�ƍH���ÈK�It��1��F�]-�;@F.E�� �||^�&�]�*Y_*�l��׽}��+x���2��ob�X��h.M����������[��2�I���;95c�K�K��Z����c�QO�?/Q�����Y��BBj�	G���  y�b_�-��f�i�q���;`����\����������*Lp>�X=j��`��*c���g�g�dA1������ˈ��\_���D���*�ɒ��\�B��:5�cht��o�a�x�zZ���	�����)�Xj��C����~�-9AD�u�������Щfw��/��j��P���혋�Sl[�b[��u�\D�i8̹��|��O/U���.�ߋ|r!c�'���i(thx��U����C��۞���@Dl+�,���KX�C{�Pj�B!�ֱ�x���*���`K�:����D2Q�'s��y�e/O�����٬�Ym�s���/K��v�o6��,cy��%r�B�h=.�k,Wf��ґ?�ӆ��}:i���(g_��x��E��Dd�$�zIh�"��)��o��|L����]�-y�!4f���v�7P�6���ȿ��wT���v�d�Y9���]���J¿F4��Gui�.�_b�{^�|���F��KVZ��E����2���E�ɓ	���9�&��G��K�YLwl��ܳl�u@�4WX��M�������N���mGOQ^�菧Q��|�a�_�D��Mªp��<�ů�� C�xB�Ń?�r �lH3�o|%J��<H�����1��[/��~KRmh�{	�5Y�>D'��TpS�>�v|ƚ�I8B���溘2�1*#EJ#���+)��z@:��`�ha.$���Ӯ#ӥ�<Hma'�h�/8TМ_�?����Z^��H��q+U�,��%+9يҜv�u89B��+�ķ}�Ye* �~�
�B��?��^0uk��NC�dG&*�.���Z�ڲ{����<,�5uƻ���a!d��-VE�k���O�l{�*�	�9�7�y������{�UP>MM�kT
��2���hIp������s0�?^��Ty�������
��_�_��u�e���Sh�R����h�����{����ukf�)5D���7z�x�{&��N�e/�ʍ�oqd�$�{`	�h���En��A���b�a���zcAu��[���u5}?��is�JA%�����`Z�J��A��P|ϱj�d��M^�!�CH�*�N��3K���1��Ydc?8�,i)~b��([s�Z��\X�A����Pl�*����OY�#I� �r�������4�tC	��B���O����8� ��j���B�,��m���*� ,)�?��S�< h(�:�VB"��ıtDϓD���C	>I�`�W����ad�X��6K�1�uP]�I�I�6�q�)
>ևU�1b\��>7_GQ�����f��ό���r6_�)������M��\g�-�(�&��Q�#)(%?��;��:�+����4����� �B��M9Q�ɧ������OU�x�2Ǜ���ʊ݈��m������Q+$�z�-[�ȃo�'�l�7ĜS)7�`ƚǖx�.?E�ʾ��=5�7YݚŴ^q2�,�m���e)�BrP��P:0�q4��ħ��5�μ����zXܠ��1#d�����&l'��͸�iM�k�f#RD��]�a�r�s�R�	�4{ᤄ^"�
�h1���E#8�\	�X�eݨ�������#�jpż[��+Kڍ=
oC/h�t�M���*^9C��+)��+���I "Xd�p.��$�� �r�ޠ:���>1���[Q��@2��B�<b{S��� !<S�h��@l���S\Q���S�E�e���o_�SX'O�V�}��_�jZn��; ��Ε�X	��@A�
��m��e����ڌd�sY�X�\{�ܷ�ݏ����Tȿ8�M^l%�?`��ل��V��x���LՓ/�:Ty�8���V@����6.&�iQ�jF�2�(�k-��M+�1�G�~v�����^Z7܋���D���!�
��y7'9jx��PN��Et����6I��4�Sn�d7��Ț;#!ڙem������N�6��!8�2b&�w7,a{�ȸ(i�-�o*b:�b�DK�E'�S�#t�f>����D/åa�((��+!���r^�*�ǣV����>�(������*	�=�Q�0�q��Tb�7�'��ٜ?�Qh�+�T�Oq�Or��ӈoj��+��ϭe%v����h�?�ù��(u�X�R��m���h!^&�3��ǯ��(i݀�"�AɎ�ǲ��+���&:�y� �(��B�vDѷ�l���g���*-��E�l�-�qQf�h�����ˢP/Dy��tӸ�Y������t�_��C�_\�H� �<_����Ɵ����]-B�N�D�)'��V��J�n7S���d!Q8R���� 5��L�-'��9�hЧ���&�N�h��R!~w�Q�X��feگ��_�4��irE���is ���V��b��5�U�#�+�G�D�}�`h#^��|��PggA��X8�6�G��;��ĉ6|�-L3���7rS�p8|��"�~�rq-sI�~R�J-v��H����!%����V�]:ރ�ӕ1|�M��w������&����&�;1�u+���^DP(IU�����=)xY�'4�_iݔn uh,f�#�y�)V&TU5.��4����W�fN'#����F�_�߭Q�@����I�q1{L��p��Τ4����Ӑ��97$��C@eU�v%�&O3���1������p�(!�؟3����N�ns����W|]�/�ܖ	V�P�<����2~�}��Q�z�hv�
���s�A�UJ�~#sKk��;����/�\��m�����[��B'G�gB<�Xi98jv(���ݥU���O��O�6&O���7)��3�'�N�O��'?4���|�`&�'y�4�����ɍ0�#V��(.����q	�_��