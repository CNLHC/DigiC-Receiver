��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk��S??Gl���'cT��N�H�V����f��=7=����@!�Q�G�b����vh�ASJ��F6$�B�!��MR|���q�E�^�Z{P�U�l��P*��S�	}��S�� � ��K}bI�yPG<�&H(��䤖�@��S�K�DQ�����E.�%֒�G�c����Ö����a琀�,,���t�T5�t��Ӄ�o�$ ��E�j�r�?�	�z�ѣ�ȓ����!Zr�
\��
���-�'�2��Ү[j �N���o�`�~$
��r6�dW���lz$�ʸ)�qc5{��22�
�����A�5D%s�.��h�#J�PVUFF��-�^��0���7���a���%��:.1�>���)o`����z�/��\/}1�	��#��83�hXZ@i��S=g�`������(�m�OjR�
�*g��A��x��z�-������O�adЦC"S��6~�;�aj/�a�*��%ad4��)rU�Ql���<9j����ډ϶ѻe�8�T��$�[�~�:�'A��\l�ů8E�E�������H]/P�os���d�*G���jέ��ߔ0e�S��6:�{
eE�"�:�3=I��48?�5��[].+�Ai3fa�o�Q����I�.��/j�VcP<�����Ē�]��v�}~ʦ��JO���Ey��&�uB���
�(���R�r���Za��$�hج�p�{��,g��
ڲ2Ǎ^Q��p'ȟfh��CQ;\~��b�݆\t).�SԹ
�, ����U��Q���U��6�\�+�i�2��.��91�N��DZ=� � �Nx�u_�@��޹ȡ43<x�Dv��<�I�{g�8�7m�Rj��8>�c�H�����?��V�n)d>���qR�\�+|M�����-�ιa*�x����#��Z^����Ě���j��) �z�٢k��3��X�-MH�B��g�ހ�6M�\G58�ص�X�Bwp�8=�>A�k����o���[��?���N-��ў���QNؙf��jV�5V2���˚���x�x�+�H(��¢�M�8l��)o�5�k�7Y�73���\hq��︐2�H�&�/;�9��B��K˻Dڻ;B���p|�!�Ǧ�7�pd�h�����lZÄ��p��TZ�5�p#����Ev>�G��F���v�Zl$n�d$�7=�Y0J��b��&���@���6��ҕd;._�&�7���<�փB��NCl���cC��*M�o#��Qp��u߄���c1	R��tU�yL��#�>�>��`��#�<΁4R
�<�a���w�"\d��Y�.I�(A�q��v�<�]��'_��H����2���	�Tp�%���4C93��bY�D0ZS#n�vG����;^{I$���df$�@�,K�R�k�(=��������fZ�װЮєW��M�8������@N#�4���q�{-A���N�Z(����c�[o2+�d��,u�3�c�G�)����}���Ju^��v�HG�����"B��QR��,�xh�FZ9���S|!�!j��ø�����T����V�����1)�0#�	�
�G��B�H[.ׯ���~�Zt_�gk���h�=D��zrW�g�(3�jR#�LqN[F~е�f٪c�rAf�6���8���f�&�5�^E��������ay��$;��Dy�\3�6 ��<s*H�3��7��L$A�!��9W>��|��R\Ȕɦ�w1�r�������8�CG��� R��?�Dw�L��j������t��:;!RǙ�D�k��
m��
�4�G���/6o����c�;@����^X��Z�0�D4��l��tXb���m�m^޶�+�ԑ���v�A�����\9����vo	 ;�)�A1�)���՘�V����\L�ML���(�N�����+��x�p�_���G�y�� �/wJ4=��>��o¦���h�R�ͭY��B�!���`P��}~����%�u�'����ū��J��~ �)��r�f�5.h��MLVt�1m���h��3����L�����R=(~�W�Z���i>y{h=~�5F��D��Jy%6{�W������>>a�}0�ጟ��-c8�v�(��Mﲨ������*�-f5H��L�}Qggs֩ �~�}�|t���� $�|�X6���&���I_<Q���,�'k/�7�D�]^wM��� �f��=�C|�X�>�ɖ⸿FH��i�����N���\�����g$�J�m�;�N��{�W:�a;+q�E���߿��E��]6���_B���_4J,�\��]�Q�[�?���a���%��+J��;�6�4�|�_9G'7�:���0�N|l�����f	�-�v��d�)N�P�]sH�/8�~��D�b��_3!�T[d? �����^n��0�icD��M�q1����SD����n�Q���Z�/�wj�}�Y(T�i�ay���tI���	���H���Sh����
B������Ƥ��S�P�ƻK�]XY���y�q1v�	h����>~ҟ�W�9	��!�,w��f���fF%��S�[���H���`�����0&�0I,X�=-tЧe�49<bڋ}T�Ɣ��w�%A�}@�:���ޜ�2��[���L�
���0�Ȯp�s��xY��l�D��r�Ä�p���^����cA���^���&Nq��ZH���d�\�W��l�۠��v���\��
q���0v8p��������'f>a�7֪d�%ͧ���'�i���1�A܁��%�T�V��Z/Y�6��8$\(�����HTNMe��O<�����\=#���N;k�|)1�I�?̓�!�����P�N��gpS|���¼<9̵�� ��	�,FX{%��WQCCJ6�х�(�����G
�	E5U�9�Y���C�)�
Y	����F�^"�d��*Ev_ѐ�2��ta+_�,�VOiz��c��=�>GX<�#O�Hǌ8�LE̼�ވ�� ����K��)M�t1�ܳ+��'�'fVr�l�Sￗ��@�z�@_��ǧWj�4
��كI���`8-pO�?�\SIؓ�ϭ$�7pބ�z5��0�!NN����N<�:U3 �L�����}��<V���W�~�-��H}�įӀ�*S�2��߫ݜ[?��Ϝ��(�,Yܵ09����òp������nku䩺����&mx�Ӯ�Z���9��� :7@\���`J����y(�t��3�pj�X��F�	���5�!(�^,v��/��ѩ1���V,��;���`6z�SNa2r�!�n��!�>�ZL5�K��#��Ǩd�?���߉�K_��)�1G'��$�3�U���2ǂ����D�g��Kg����:g~bt����!�������-�FA��`K���-�:[(12�M�,Ā��/#9����l��
׻�j���)Ղ����HFM,p�H�T�ݣ�_�pIB#���sx�oZ3�2I��0�?��y�5�;�+`6	�*��`%�������-���t<�t,G��Z@I�o�v
����Ν����G�M\��� ��=�R'��i����'m*����'NpU���U:~bC�B�K����E��dc�%�+�^R�&�B�M�i���a�.�i����[|N�~Me�-�0ٛ����DTz��v��|��:�)&F�C�1r�����3kUo�<i���
nኁQ8@@�9����t�Mײ����~��=mR��V��2g�m��sW*lpA�r�L����=H���7����4������l/�mKS+��:Ǐ�5�O�kW~�Ov���U�J�U'^�n�dN�H�7���VĬ�Rҽa�_P�yf1Ҋ� c��,a�&���s�c�\�*I)�u����L"=�e/��kK�9��k�����?�]?��5�<g�K���Y:��c�2�%�����㌙�{��pp��W�,�`������\>|r�$�~{��a���= ��{�Ʃ�X�K<(����3l	%��ψb|�L�A�S̓&jb�ٛ�����y=���a��wC(v��lv%�JQ@Gc�hhw�Jry[��xTa�Bb�'Kדm��&e`��Ҹd���*�H�c�厞�����,A\B�4� ��iN�6T���@�ӵmu��m/զ��{������`=}�i/l(�V�J1�c���!�Y!���3���.��4��gR}�=���t�_�Sox�xѰ1�Z��ͱ�,�����K)�!���LU�!�+�K�
4Rf��K�8�~�?��ኯ/�^VB�oZr��p��a#��="�x\N�~�$8�Z�V��P��ZBt�I�v�u��:�2h��q��fP�w�Fz�(Pj^6�����g�#������<����L�g\`u��8��\���(`�i4�𣋅x�+}tf�Kh��7�er��j���G�Bf���eh?Y��\�́�h_���I4a���$�[и)N�n��D������
����D�%�u�QbX�9V�����	�?��"�y����߄�,L]-0E�.����M5��7���$`y��-кNL��T&&�T��4M>!�5� �
�;������$��-���r��N�䭆d���J�019Z݀/3�/r�����*.�+X���-�=^�K�[�dP �k
F6�_���c�	י Y�������Us�ρC�DD�E_�e�8�Պ�y��c��h,*ޒd�Z� �x-����C7L3 ��u0���Dv�����e���F�Fl��b�p 9ׯR%���y� kJ�$x~�1���S�Ed�-�gu�m�O�xL�ά��(�I�v�l�Gy�%6�|d�c���jN+V��)���	9U`���⃷9���r�?�7��=�B<0U�r�����V���j9D�O)6=�=��czC ��-�Q��pPmy,"y&�n���ע��cs�O9M��[Y\ܳl��"�LM���ۘ5N���P}("�4d�J��`��|S?�hY�2R~oWv��L��5��w��hQ��M�����"N��O��M�����~���>/�}�!�@�i�o��S��� ��L�ۦ(��Сmo(Lގ��ڸ}/�-<��4��o0��? 1���͡4Z>D4�؅Ҏ��n�<�����ɼ���� �6�̫�c�Pԗ.�b	��c�1X!�Z*r��XĄ��>�'���:$�.j>���$����p��S���L��A5���Mn�<\�b�7V�e4Ic��)�*f��40���l!�q�@��τ��ћ3!*ڹ�����I�����e�)|��k�x��+����ڠ�gt�M7�6l�FVю�мR0�p�u�R��R}���
�8���E�
��9slwe,J��1��Q�ʞ5��c���7�5sG�ɞ������su��=�>7��ρL����[�`�����X4��(�~^�K�Ξ��V��39:ƚ�tߺ'�	^�L(�W�t�����>�u��Ok4Q�i@�ޱ��rKԽP2��HX�x��*ͻZ�B��<�\��?L�#R��EŨP2ۀ�s�#�k �i��J�G�؜/r��&wv!�zG�W���o}�bhu͙���O��Z�I�0�@�B�y��˵�ע��s�δ;��P ��MS'��@���3©��t�k����;i꽣�j�TzI�MEo����iQ�8kC�V<K1�i�����|&�c/C,Cs�J��"䍷��������RV�c�,��L�K]�
G�f���@U߈$� HO��Qi|�iv��ޞ��ɠ:6@`^��#"��ַ�n�������������b��ַ��2�b�oW��� Μ-�3����ז��I�FNw��s�������{9V�a�����^lt|L�P�U����� q�6a`[G-m&dvY�e9YX�T�lc� rA�
uk	���33�z�B��``�pRir��gt�1N۔���ƣ�x�ji�\>�;��b��|��1k�U���פ���=��X�V� ��q�ڻ�>Knt�`8{fbC&9ҐäZ��I!(TQI�����)�҂�>�s<���<u2�d��k�ku�j��h>�?Y u4B�q��[�K����B��)���Ϩ�,�.��=Z��=K�)=}?�\I�f�J����<��w駖x��T}�0ܼ�����~�j�I��n)i%A�9-����Fw�OE����R�ί��*�M'�����o[�[b�y���M�{�b�a=OSs!��]E\/��J��x~ �Mk�[�:H~$u��fc�B6]�êlT7E������9��9�Cg���u9�Iܯ��c���@�'.$�*DnJٌ,֑��>�,ɖew��);H�L����B�	c�ի��D?�շ�V/�Su��gv���C������d��Ǯ��M2*���N?)���\r���,�݁�ĨH_f־��L�qJA(��V�Fӌ��_$W��Ã{̢Y��V���F�������,H���^Ӄ����p�CKa��gˠ=�>� P0H����Fc'�?=绵�eD��pl,��d���yB�^^_ �����1`��4��q�wi�[��e�3�]B�Z�v���_u�URna���c-���h6+Ttl4A�#��x)5�=�զ(PD�lWr+q79�v���g�5��=�G��圉Ӣ��rX�p~N�~p��E�J��9�~?�7��P�ޔ8|<�2�6�T�3c��T�=�!=<��z�1-����-�!Xi�?�n��5hjt�T������|Z��e����ӵ��$NQ��F�}-� ��G�⥿�9����K�iWo��ܻ;v�Ò@����q�(������0&�ʞ��cE�#y#�С0��	V�i�K� �ʘ�3E��ž��	��:�*X��~d��p�B�q H��گI�
��:�����w>���7]T�?���ᗉ:�փ�V��jjJ��Qe�	��u�ي#��Y�T�e�@]9QY�OB�0�_�M`���';ߵ�57z�=��L�/���$�2$��E6�V�J/�V�T0|G�T9_�g�yz�DM���\�ȝ���F���vr�>b�,�wQ.�%�(˕�����ˎƬ��K������,���PBrx	��������fߟ@�	々�.�{�w��