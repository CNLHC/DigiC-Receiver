��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���N��`�G��y�]"UѪ�e�����rb��E�B����V��3�_`��%C�a�B�U2�;��S�;s֑�qm�r��n�B�/�z�h Y�f8� �P��@�Fx�����=ֱ�8���`�D�$*�B����wɥ�4�A���V_6}��\f�Deh;rfT�Jv8�X(����:�����_A���H$�+��(���S����-g=�;Y8:,.��s+s*�2����Ċ2��6���s�x5rݨ-����\��(;&�5^��p�Q�q��j'¿�������Wc}	������b�
�8�{���������K��JJ��;>({`_��ˆ��;�1$�4�1,6e�}�Q����]�i��L�[7�ѝ��%��|%����q+���E������-��T���m�I�/0���jCJ�_��q]�V� 1��)�=��/?=�=�^�JO����)`��F��rR�%3��7|d�P�y�!}�g���(����F��H]z"�f���S�����0)��oٓ�=��Ę�*#�ȍ�*}/ ۖs��������/�69Y�?j��86��駴r#�.S��zߛ{1�RE��ªm����i�,����X��#�n�j��2Hx����g¦�x1����T=(�}�]KT}�z���籲'��w����n�+�a��f�4?��9�>\�2��z��O�S�]�ᚵM�!��7*kR-��E��z�jm��V4Q�0R���fc�ΙĢ��`?�s@yO(;P��>X�cZ�s����|��;��
��h;l�qq����#
p�4�1��<D��2��"��T�x�[�<�%��j��W�@�z��r���zu�h��x�O�-FěoK'�%���$Ř�(S����\��p�Υ����5�_6[��A�g$��C	�`s�Ef*���y�	���/=*�<��O� �}�Z^�!9�%��B�m���zw�2{�P߬wu��\�lG�I�{Rm��h����dp��d/7U����X������K���o��m����6��w���}p��q� Ǜ�K�R�cp�h��325[�f��w��?f�fw��� �k�V��Ջ'������Ef�z�U����h~��a]��Ww9���.*��2�:Ѧ�L|��@%İ������N�j
�^؎|�<2�Ї]!���:�`&Yx������uR@eh+�uc6ֆ��
���}�ks^�"�82m��v���W% z�J+�����i��vE��haw '�\�P6�|���;�,!v_'j��~���ڦ�S8?O�������W�"f�؆�}�r�����Y��t�R�#7L���QD߱Xua���	c��"M%�@Tm���>_7��PKOV���A���C�7��[l��9�r"d�B6�����oB9�F�5�g�J��e=�}w#�������;�,��6��#��n��挐��o��tӳn��U�׺��^��]���ܼ��2��/�p?3���I�*���(J��_5�Ǔ)��YiB�����9��]i���N�Gi��d�*$9e&���&}`#
��Tq̺�	�	$췵#W�;o�c��1
"�����H��m+R�ju�Rb���GI��8�yX㋑��brQOσh�ɂ\��G�c��ߚ
Cv�S���a��WHb�OF�}~;�&M��I��(�QǱ�)0��)�/e��|PI��D�y��|��i���ݐ��U�k1�/�Kv"�)���^��.��y�d�[�쬌?�Z|�EF�7"^H|���LЋ�Ҵ}*���1T�u�	v��b�s��/ݳ�����m��H��,�Թ�h���͟5|2�36n�g��y�����̓'�^�6�m�"5��o�Zp~IT)�1P����l+Stj�+y��ar�2G���S��{�Y��S�W&q�f�A6t}X�d\����}���I��z�T{�e)�F)p�Y���#`h3���d�p
����u�����r��9� �Y��B���n*���B6�R���˖��7�o_��?�<����U��9?.��u?OA�S�C�`�nf4��2�G7�N=r�!���0��e�N�{�>��F��^�(� ~�%�ޕ�r�����Ӥ�l���� �|�͎n"�6�:�����;�1����%�!��N�������5���
-H�G����m����z�ܻ����|�.� ��o�O����v2\��6#����&*��</��#��<�K+��c����U��Ô*:�[���6ދVd���՛��o�I�,bF�(��n,�c|�C��oUI��k�	$4���%=�{��x���b�ץ���ZH��\7��,>�� �DÜ��c��-Ϗ�;���h��?W����@�1ŏr����ڡ;/�֑>�pè�B��t0,|�f�ާ%�ɗ"W:D���ȳ1�˔���
��S�#�F�tQ�V<��<R����o�Θ���0�_N��0rt�:�r9�!��9Lt��|?�w��^�%H�^��B��e����e+_Wo��F'�Q�`��=B;>��KX�=��('3���#p�CA�tפ{�N�8�$�*S��tD�
lpqV��4���(��.a��񆁎[��]�����}�s�nʁǪ�5�A���%��8���iD�H��@Ii@��	�{#�s�N`�Z��0�T���[[f�Оi?3CO��zfAސ����'�|�%x\ćfQ}�ם�x�'$>�Z�P7��˚�Oؑ�aݓ��x	"6������íV�F5�e�u%�A
IͲN���Sy�i��m��� �~���	Q����&m����i��0p�F6��ಽ��$`��C�/�(c|�
���姑t��=j�p�7����H�]k_�^-�(��_�A�����Akp�#�o�\x��o���9>3��~��n�eJS����/�2]�Pmz�az����#uegxZ�𛂖,��L0�4O7|=z�z�$�T��������Om:�0R�Z�<Jak�(Nl5�����
�|����5�gȖ|�	���t��];�|��6����h%L�,tkM�]��4MpE����od�γ|7h�
�Q���sHy��1j�ൎ��������Afa�ZV�}i��Mj�<r�(�\ɬ��B�j�y�ɂ��)��E��7>��)���֗��	~@��n��=%�cy�p�Q�h���	5,.�_��BqӍ<�v.�u��(�ŋ��d]�rt�F�5�̄0ּ�6�w�7|�}[��c�dMRm{�,e�9�C>k�}���)���Ui�2{�,^��T6Z7sj�M�)m�gz�ҳb�d�CS>�.�|�h@Û��]�7�K��V<�̀��N�a|PP�<�k�)��F@�j4���#��%[�&�a��m�j���f�QO�T�Zk�w
�0
K>@�)�Cx~����k�K��*J�ĂR��6�*t7�W����l^�؇S�eK������.����˴��|��3=껭�i4S0@�3����*OF����_D�+�|�b��j��x�t�>t!�n�����c�<�?x�����0��u���S�5�\~�#�W*���m�=��A�oD�j˚@4���0��8D�D8��45M]c���)w� �Eޏ�y'�DB
J������ҫ�U���v�qH��/�5������	&I��v<E����w�Зޏ�MB/�Sݱ=��Ų-�~�pb�Ū-E�W�d;���&BB�����(GC!fX�`�x�"4�-<T���2���nE�y�J7����Wo�F�db��U���2e�"&�w�r��W)��ͣRc�fL�IH�j5�o��u׺��/nɱ���C�7�9Μ�Ԯ⿿ʲ�3�G}�h�M"1�E�:޼f~�N��7Z�S�� B��^�&��M�5�橛5�=Z�U�W���U�YJ��ߗ��	 �cTg�K�W7I���:Uh����Dm ����"CJ�L��PPfL�!v9�؆-�5����8��٘U6�K#i,�
5�
�a&xdX���D�$�<�����E�?��Ҟ�����l�=���*�ܒK٘hـ���q�Zcw��m�r쬣6�Ե�o�~+�ȱ���I/нɒ$̴�|p�É��p)��kܒ�>g����:�O9@}��� ��k]J��������W��!�W�ˑc
ҏ�R�#'�e ȁ���,��P���N�YZ��P>3�U��z�2�U	+�ga�A�l�r���g!
��s,}Q1	II�%VH�6��v:�K�4�|O2�5O�5Q��Oȼ0���� i��+�s5��h:ZE�@�C�R���~��I�m�M�dF�5޹�Z�t7�8"�W߸`��F�W��趺R��Rh�����%~%��[��������Nd���$��X)����@f@� �y��|��ta����
5*9����S%������W+��B��B"�̛���%���q�<���H�${��z��{8{�z�v��1�3!���x�ĳ��~t�JN����@��X��Z,b��۳�LI�! 1%[�5�O�NGI;��n��p�w ��kY��wZ!,�'�Fe1S1J�^�i���F�R���鑬߮�am�����1d��* �X�F�_G ��j��A�#�~���{s��*�RݘNV��z�?���3��ph��M�$NJ�؇�
�{�qSe2�kW�-�{*-*|�5"�����a�i�(�r}�J3�5#d]�� ô.�3{8�*@�IC���R��$��"U~8:20Ea�ʤm���y"i�P/�н��"^�Ĥi�����~�JlÜ���f��A��4;)䔤�ׇ@eG�.�u4ah��F����k]0�9{�z^��p��}M^fwͨ�� �)B�P	��W�,`c�����<`�o��DH���"�}ɩ�|W��4��>뫬Aٮ8DH|��Osӕ��`�l
h��pLK/z<�#T���Y��NV�$ �e�波�vDh��@|
���=����V?J��j2$i���"p�)ӝ�T���ϩ��{:>�;����K�}?ˢ�a�E� זl����%u���~������mD��D�(ҥ;DgE7�x�&�"a [@��*;/X���?�g�:B�= �]��ͣ蛩��85���s��V>@�c���S74G_����]����g�#�,m<��@�� ��)j�����ف�O��k��ܲJ�OY��/c����#!kz���r:��q��V��+GR���0�J��p�B�-KA�\�<s���|=��=?䳂��o"79�g{1}M���Ĭv������������QM�^U�	����M���Tb���k�zi��{���&=��3K�;�LSâr��~�(Ֆ�nc������Ӳ��u�F��2h�g�o}Xc���X��<�w�L�rſ�CWr��U�"�$*!�!� >����2�����0T�����)m�;h�˂��u�(\��MCB��[3��	i�3l2Վ�6zݣ����|�y�u:h�_��⏃�Vs��E)o=��[�en���<�]q�Q�Ǎ���fr\�7��7����5D.�(�s$��.�݀�G}
4�Vd�o�q�'���Xc)�!�R4��,
�6��r��L:#�	 �|�I�x��p�3�v�sZt;Bm�#����B@lH?�{Q�Q��#>��6u�z�Z��o%�����'X� `����d��(����*�K���?�.�2�^�s��������ؚ����V7�y��\�"�8�����>I�r���@{������g��˙������<P�֏F���MC��%�)�	c4�F¬�/d�3�8���y�-�%�q�@�4�.�Җ�~:��-�@$:�^��.�+����V���[�� �p!8Y�k�|�0��Z'��#e%q;s�N?o�*�|�m����������s%N�{0��/�<�vu�^���*2�'z�ف�=�R^�ǳB����Q��?�hЇ&
~����[�!�kc�[��O�=�P��
���B��^u�"���g���y �ӽ\̊�‽���0��#(��u���ٯ{Y ����~15���Mg�C<�)�Ce=����ʺ�������[/��O&���Dtee�,��#T��ݢ�(��M���:�y:��IGg0�,[_P�i�q �y���j2��O�,�(�z�G͸�7��H}I½!�zj^~ya �H�RSvs��Teb�dq�������6�g<�Ѝ!wp�>���K�P�y?�O0�GGc��NEߤ�S�Uh8���EV���*4�.M�
�}��f|�IRh����]U� �8�!Ķ�y�ط5����\�>�E/@v֓N#"�f�p�J��Sũ)�,�.���=:T=�O�ӔJģ�N��`[DT��ë+���b�`�I�	�B0����z
Y��߇�� �����).�b�u�ZKdĠ֬4���Z������� �7�ùۈs�Cn�������/5���9��q��ׁ��e�e����t�S��������� ���M�U�x��u��W7����>8�~��yĖd��bz��s�s}� U��GL��$ԁ
�M"i?H�˦����/��c*)`�Z2q�nO4~���Kl�ґY�H����E�9%�� ����Z[�)��!a�$���Mכ�\k��OW�݊��jS�BԪ<;�xPo�M��hA��V�b��zWt��t\
6Y�U�@6Y��E<��	#�21��r��A�y\�V��y�����N��T����}�Q���;va�^�-��+�Ģ[FMo^L���c�"@�*
�j!�E"��G}�z��i.Dwy��
�Q����WY����b �L�:� �wY�[��m���J��JW}��4L~��t*唘���2���� o\\<��O��O2���ި
T%�rE��N����Hm�y�����~+�`"S�Tz^��FYl��.�@S�t�G-�πz�$��U���g���������Jb;�H��?���O�A�� �|�������X����=���Vm�~� �4p�_:�u:β� ��6��.V%�)�/���R'��T�4��x�9,��������g>����F_H.�biC;�z�}�v�h�4�������@m̪�'��y!Tq4��$�W���U_��ϑp�᫵hqo�]�y1����h��ǒ�&�����*p&�l��2�ڱ��c~�$�Q����(���i��z��24�JJ`-l^P+�_i��[��[���EkS�������j|E�������f7N��Dic������v�m@���-��4v�����c��#x2?� �"��	@
K�M��=Z��^�4I��J)w�kn	�꒽њ�d��c�3`�m�ȴ��p3�:��#p���#�I���#k�Լ�+!��b6�.\HGN�E��zF�z2ь���ޝLKzl��q�����E�ʼK޷gj񝪓�~NV�������|��3^~ʮ�Ĺ��63K�P��#%�[2����Z�)�y�l;������u�؇����Ӓ���*a\�KYk�lDOzhr�CT�m��p�$B��#����z:��NT���v0�9�^/���zx��*�w����d�z�w�C�Oe��)/��he�{����DU�ZX��C2�mDBM��\y��f��g�`�xXl�f߄|>)���0:�P�a�'�ϑ)o7G�Pn'�����DRuͲ�����E�iyC�>���f̘�	�cD�'Sm��ǰ	$�ܼ$#��f���us^[\��_Eb�Y�j-t��;:�	�]P�����֞��ɱܰ�ai��ז�:6����L�驨S"@B�KN*O��jG��oA���o+��0ұ�RX�^4��R���C�. �i^8�D�s���5Z��ɀ`��.�ؿ�#�����75�+a���fr��:X���p��r�ᷱt�B6�i=m���i2��/������t-EYw֜sm8��GR}�.Va{E�=�Җ�{|��R� �[]�Z]�q�E�*��Em%�QW�vEoFٵ?G���!�h}���K��AR\v?ՐRּ|���ED�]5F�X��Vx�>t�?Wgɠ@���B`a#]l�"s�B��t�?�� \2�/�
�f�lC'�w���0�y+��:����5�B{�K�\,����$ܿ���1����������2�����l=��ҵ+��������I}�	��I������[�B�h��[+g�v�Ԑ�:�Ml��u�W��Ĺ��K߰"�U�R��h�9�S�d���@���n�)��#�ݞ!ݎ��y!ت�
�|�k��-�_'�_v��P��Z�֪������JL�MG׀|Ó��j!���0����a�,���;�X�>��\��]lG�\���L�\7P`��vJQ�Q���Ӊ;��ӟhR倰��p�`hE9S���Q��}P�����`ؔ�?&��ل0��宔Ū��j�㷼,�:6L]�㎾~(�D�����6H�3m`�S�8��)TdQ,������ܤ��|-$@F���zߵ����Z_f��aJ���A���lU���+GK�����ɣ6c�F� r�󞡿m�U�>|f�eXS�6�5В��OV��XG���Z{���O�5�Ҿ�a��`[�ν�LT?���������5y�+,�u�V�Z�
FY4Y��&�gL9�6��0#3Z	 G��D���P�*&1�,b7ߛ�7ʽ��,�tWf���DY֒6�F�%��\�xX�Ez�p��hlu��;?��hf0r�m?�Q8����I%�ލ|U�	���n��}ȅ�]�f�/���&�����_�Ҿ�������E6'�^AKQ״)���o� K����8������*��_�"@������!%��!��4�^u��g��Vdߨ��vlifJ:J­"�d�n��v���@!N�i�7�. gh\�͂I�.�=گ�nwr��w�X3o�kMx�E�p��q���	���a�>Z��`�����l�5pT��YY���]���B.U@�v@��-j�b��j�M��4�$ۈ��@�N	��Jm0_��
#QP��p+����$�շ�v�����#��ŧS*�V���'���&��|=N�����N���M�S���t#���7kk_�8�L���;��Gy���)T�k�L1�T��	C�z� %{��5��Ȗ� "�j��l�S*,`u��=�q�a{6i<�Y�v��T~ħHZ�ϛ�oI/#���ܗ�W��u��xl�R�Mtޅ�3)ꐰ)ü7��%�M�}�qd0/o؃���8��:��N���Z��2��V�}��n���_:���+P5JsʹL9��da�^#Lms���K������>��@��p�O�q>��֞Q�
��9�{9�k\{@\�(�/���nf����u�a��!%��(��Q���u���"]͚�{�fz�_���B��ӹ��\�ۆ�m��R��I��/N���jI��]s1O*`}��Asbz�Z�T��h/2���*����|u�u�+��1W����v�~����r@�pC��ʢ�?����!�cFρ\���k�]�!ډ�1�=�jx 5uGa\�`@�L��3���!!H�Lv)�&���lS��r����axQ&_qC6�gC��7�������a�҂���3W�G/����b|�:�~�B�q��<��*|��?��CϹrb�U�G��o[~�^���/�u2���I2{�~
iadX'���c'��d͍��һ��I��?`䉢�^7A�lg<�d�ߵܤ���� ���
����͋*��>g	�����'B��,o:V�d�0<l�6�"�NFv�	Ơv^9
B;#2֊���Q��� ��2�@w�Ww	G��H)���6�n�;P��,��EXԫ�T���[�X�A�{}�����)�&v����B��塝b�f_O!{/-d���i\P�����4ܢo%o�����W�B"��D�4�7�u��FJXb���M,������^�R��8���@Lb�B���jv+P�	F[�f��qJK�{�*��J��D��J��K��`��[���H���~>YV�-elh˞����?<J�f�����q���4w`|��y`W����4����I�%�*�z��uޒ�F5z7��kݐ3K0����[=� T�N�R��@&o*��g��Ug$S@��Z�>l����>ك��i"���&��F+%��%y��s?�[f{���L_a�<j�<������9T�{���ל��Վ�W?�4�>��\�#6��?�:���w@#�s�uU�F{��2�H
e��vr�?�G��Š�R=�~Wa�cB�A�B?PiR��S�X���=��S�~U�O����ΐ�tP��׃t��!��'��4~��s�+�V	��5�F/�ݹ]��#B(0�ނj��ڢ���?4暱.H~bҗ���`A����y�?j1�[m�Yȓ��e_������i����l�x�-�T����]b��I)��6�5�Pӯ�P,���L��l���po^6Ŭ�p�NKm�9Ȏ}|␱`��޳zϡzM%F �٬�$�Lxn���������U���U�)�kk���D�Di�#ߕcZe"������r&�kcS��q�|bo�D�p�ᒧ���%�덦a�E'�2>����kSJP�ۗN�f+2.NոZ�84�7�G���i��
�.�k;ܹ���Y%�y͜�Hj���!G�UaG+
��r@<���,ˊ�/\)�x�~�����C��I���9�ܥ����cKnl�^֝�ʝ	%���Le���{���Io9���(Aw�U�ϳ��A�K���+qq&�]A���i��taY�j~�@\�Kg/�_C;q�S�st��z7���Q}���+v�U�'����]�dzO�����L/Wq%m���8�� Κ�N�ۜ�j�W�@̘�#Rꖎa�H�yb����C8m3�]ֵ� 5�@~�{�ݺV"�������3�?r���b�s5O?�]v(�b���chM�y�G�)F�c7K���'�N^���qn��u�z���	�0�/M��˟/�=�3i��0�;\���*���F>������ XTw�&��9
�f�絇!ċ�eFS�<�����	���0lnb=���o,��`��K^���w$�~@~��P�@���WYR��}i���,q��h8,�F����D��Ҫu��ckgfo/&��)*.���{KtӟS���iR�b��a�[�<p�1��W^(�mLy?�@�2�\��F+��h��K�շ�D�Y�E@V��,�l�V��IΞׄ�Qaez�U����we9�l2���g�f,`���:,�!ORl�
:��m\�f57 Y�J4�G:b�N�T�/�"%M�w�Ӡ��ʍg�� 2�2��p��L�3�}�kԝ��I>�.Sd����)��A����Qˊy��ysu������$��H{s��}�V �f�ɵf����o����4��"��rͫ ©y`��F�'��¿�e5��9�G`���:�ѓ�YMe .�r��A�s�K� �*<�U	"�f�	��y�N�����թ�]�I���/}��֭)Je9A g��9�5�]ݾ��1��t��4�����C?U4;#t�7H���E�YK}�	 ��딈�2�nl����Q;<z�<�$`린�^�]���}��2qb���4�@g�l���2VN!�"�2����v��1�0k;�I/N0��_?r42���߳�)�o��O��\�6�w`k�r�/�H��}"5�2�/���:���.�Q3�ڡ�L�#�o��qc��(TH+�����lR�p:�4���C4�� Z�fe�č�1%�Ҽ�}��(���De���n��F�ܑh��4;:l6�c}I�����4�9�z�V,�\�rF6�n���[�\��#>�����r��#�<�\�Eң���M���o�}�&�YmG��9�²:!�⻝��
o�$����������v�>j���Kq�ź��;�Z2ROi	�ĸ�c˱C�g���K\��b؋�	�������t ��n��3�ʳN�n� �������Y�ax���'f}�%��^h�/x�c�\Ȉ�&j0}y�	].����,�V�_��PqY��0�����;��r�'��ϸ~o�o��[��f��~Р�{@�~\��-�Gv�٧C�v똹��s�"�$؞E�G�T"�D��-���>Ωdq4#���Y�Ю:�Aᝬ�r�8i�1�TZ�Y�I�),氊�%�F~d(���E�7�U����}h��mM�/�^����}3�o;�T��>����b���*�A�0d�p�Ŵ��M<OA#z|d�gG�e~du�r(א��>%oV~�V@�-Y�?�`�a2�����7��UL ��[&�F�-�D��c.ճ>fؔ����<[���d�e�`ߥ�l����Jׅ����J�Dƽ~�-���Sg� Mq����^Y^�**#��5����jLp\��ГvM'%�8:���L���S�"�@�?Z�&w}q����A碒ʡ+S33���[�Ԯ}��r&�~$�=!� f��ZJ����/��3v0�5��
ȁ������=��rﺠ/�J4���nO[�h wӪB:d��V�c���ز�Y���a��!>rY��q�MR��.�"��	`x>fP��k���bJ�����MR�9Tg���0�8fl���Np����QI�E����ˍ���'��I����Jq'+b�,����,�/�|�٭��j��Hlt���c�t�h�o�Ե��G^Y>1���{k���l�B+� �B�#�y:��d-�C�5P� 俗���H�$�²����>�0J�!���Z0��^H��a�;�� �X���%�v�o�*ݓS�mEM��4���}�w��e��-6��.���{c�y�ǣ󡹍Y�ǖ��^��?��UI�)y�K��P�
�'�Ab��݈	4�	-藼��,%������3��E(8!��	A���/���_���f}�bJ	��I�N]��f��o�r�"�=X_/��ma$�+^�[�� ��|�"�W�g�]�,f�*n�+4�[�R��x׺^1��+��б `�}�1����O����S�@�^�H2�Z�x�L�ꓙ!hW��i�D�5^?<�.͏���x�T�e��X+�<�[k�HAx�亚%�~&��5�#���K�V�=�i8���K {�$��-���0�CjȔ������.SJ��j���b
��@�K�`��+�ڝ,G�_��5�ϰ���>;k��V���H9P��c���i\ �Z`c߱<ޝ�w�w����἟�$��#�3��臛��k�d��>Z.��MW�~|$�0,5�O���l�&����zPIj���ţsrx�PCuZ��n �σ��͡��L�,��n��.��g1�h�#�m<���0���cN�zʴ�w��t��
�
D{���Қ�Z�h:�2���A�iB U
���I��4�<+����YJ�o�th�I�?�/YP��y�r0��˶�_R���[n��+��I��hj�+��7�HQO�0�A����Yez�B�d�w���]X����Tվ-h$œ�8T=v�m�!�Hz�F�G��3���=$�+h_x�����~�(�A�Տ�K��ޅD�B#�o�8�b�_��	!U�>^S�n��%���{D;��5�A��$�E�ܮ��k���6�� ��s�!��^�FYZy���yLyx�oF{�Ń����"i:��oq����k���>dD�u('��r��S����nQտ��H���]�z�V�-p�OZtS� D��
����&�RW����}sx�e�G������*��o�����Z�@l&�V�{��Z}��a��s4����^�zp�0����SН�=T;����\�򁠡�-�ƈz���5�[���Nb�;�1v��4'iզ�As�uͲ[.(֍��T���HG��i�.4���&��;�+�.���F����1��z<�P��dц�S|a�cG�y�o~��j�\h,h���;����l1�~��颿���%l��Eڠ���FR]�W��`�c�9��?/���X��U����"�I�
Z	�hIs�Ʋf�S/�h�.s�${�F��wM�/Eco���oֿeX����V�g�J+��gB�Tn6D*�&fr��O���9�����2
F����g����-<ޝ����~�Z���ڊ����������oi��S>����k�>(^US �k
����!b�J�yx��zn�>�-�Dl���N����t$���܋YyBm�c� V\)��G��{�(��7�qn<��V�T�UGZ�'}�|v�rvgY����[�`�A"b6��&R��w}yM8�U�嗌��uڄ��U\����_b87��D�� }��0��Ɂ���5{��W�>=B22jX6�a�*c�l�`��Hm"By��~�<|·^��,�(l�*&�������g����77Hͽ�7���=�Iȓѷ�C��N5�������Da`>�������I��|8��&1\��f���+Z�r>��F3lMu�v���X�� �x6���8��M���'�Ƀ+��&D�	��o5�.HE����ʓ��� �9Y�����\�/��m��\'O��ﳟ�pR��E��}$l��E������QF��X���
5w�ґEh��2;H�p�`y�����������?��6����-�,[u�ʷh��&A�Jʟ�����DI�]���]��Rr%�<⒯�Q�IL�ۛ������)N�����" �lEc%k��;�;�	x����9��:�[�{A�z��WЪ>W���>L��
GD��㏒#�*D'Kb�C`AI�(HjS��g�71������)���bX<:i�G�O,��ƥ3���_��؈+��(�Vvbyh+L�{�-����5��%R�b��@��e�K�ټ�����<b�N
��L��h�_�jHK�>�@�򰣆J����Bh$�k�q�D���^-L���A�4hH��o�"�a�]��v�YK�CWh��\���g�� ƽ�yk	j�y�<C7n�f���oCA:���l��/����d��'��9V"ق?�N��]m#����`h#����?*"+�O�d�d.OV��� ��iaǒ��e�څlF�+%�B�Q#��I1܋�u�<�D�e��᧩�����Q��+�Gy�+�p�i��Q���0�ȞY�D�`� ���ڼߓy�Hy@�G���k2.���N���$���CK�>>Ne���QP٘�rr���(�.����N�?BE	�f���H>�WD���TO���o5Z��deYn���M����(�R���6�	"s�>����~{tMJN�o�  ��Lv�;,k_�f9�����$K��K�������̖1Z
���;7?�)��џ�B�l�J��l��5p�48��y�3�]J��"e�~�#���5_������p�de�*�p�}�Z�஀�П�[��H�X���,��a�H^�{+)/�NJ�4��^�����s��E{F���D����`\`�	���2ur�r�}�d��lͫ@���S��v�|�}׬'�	��m�;OZ�AZ�D	x��-v��9��^��hH>��E[���4P1E%DC�P&}�1Լ!	;�=��2st�B��l��dA�J�� ��}'2B�.@-x,�灄o؍1���l�d�-�2�Y�/%�q�*�'ّ�9�� �#�ﺲ5v�`��qC�x�-V5�4�ܑb�㨵2�3�7(0z�9'G�~�=����
�*f��u��	����>��^O}�6m�A����-3o�K�Lr7�Sx7�+\X��)^�Y�$rç����=��ʽ�h���e�R����إ��"���15˚V���{욼�[��w��cLnU��f��q+gL�8C����b��#��3��`��Z>�5Ӝ�!iٰ#���Y�� I��n��A�qX�Ԏ�,�R�Ě�q�(��,�:C"T̷'�q��Q��,��L��ҁ��ǹU-��~�		����(=��γc�EN��ހ���(�ȑ��؎h�o�Vf�����3��]�e�k�-|��`�[�IsbG�V M��O��ǚ�sȀ��j���G���ۤ�o�NÎ݀�;,!� ����5>��*u�Y�;��C��A�����t��oG*Y���� J�SГ�jK��[��,�:xgs��D���vv{#�������Q��	��g��_^�A}"C+��,��\��h?%W���e�������]�5�I=(!J��;�Q�*����0�E{���?KY*x��|�eP�.K��k
����vcw%�f�W˻5��|�(�}U�U����u ا*ݬ�x'Ԉб�ׂ��p�����%�N��9�(Cx��i������P�er���M�,�f�����s�q��H�fgwFJX?9M�1��*��&��Y
���w�+�̆�XJ��V��k�(��<��Z���j\8@�hQ��.��*'��)������;���}y���T�+�q�ڼ��HǌT��˸��������@�V7o��tt\�G�JV�6�X�,X��Vs���űnswL)���B�2��B��� |j��1�IFb�}bQ�L�`׈�{���#yd[q�i��`�rN���䮓]q���&�Q2��ɵ�ud�5���80�B'�{��c�C堂�ol��{\�2;�p��m�Ӱ4U��H��pmK^v"#��������_kgط�P����>�I@a�(+�L��nT�ɅZ��>t�7��fy��+��
F͏0��:.ү_#�g����5�H��5($�f���ɋu��E�_�sE_����F�1��C����<)"��8�O���r�a��,�;��=V�$�CӖY���J,��`�Y��`sq����K�̷nkɆ��g���4���.��pkk^h�1��u�?�1F��0Y�qV���N�,MK�E�I��;d��?)a��]i~�"��
#�!Z��V�@?��V}v�rOo���k �y~$;֩�b�q��˩S���UnA ����"��;T�NL?��A��iɃLp���nE��a3�?j�h= ���Y;����g[��8��/!���~��gZ�`���M�%4J�S5F�B �� U���ufO�̮s��v�А�Έd@l8��.	>-�7A);8^b?P�S<1�z{{�6$Q��Ho�x�+E�>���yű`��u_��k�ܠó[<���yK4��T5��'n��:�*��EX݈�
����|8��\o�G^��w�0ώъ�O�:��R�����p�T<h���t��+��|�	��{�,���X-�<��f=�.pL29�\ϣK����5s���Ј,�m��eە���.���}�S������(У���@����^&�6�Pwq�Q2���FL�l���X�N"�E���J���&��C�~x��=�T�zG�WJ�ʇ�=�c�g�k���
O9nb��]r�4
ћ���`w@�C��8T�����٠�]���(H�:e��i�%`���^�u��ӂ���ERe|I��o�M��P��C��Ցq�NX7�KSؐ!���J�Ν�!i�L)}�'8�k����q�D�@v��db_&ŕ[��(���Q��aa����/C.��SaC"�/@�,J� �R�;I�:���&��gX G��Zh������J)�Hޟa�9.%�_�����t*�NB��+�����k�,L��{�sW#b��`�(��Ί�����0]üf�,���1��&qq�H*����J��$:6*��G�;D��� li뻮Nw�#�Y��"�!��v ��y|��W�����߼7�k$QJ�.��V^_�ܖ�r:�Z�)��NJ8q�'��a���]��*Xw�(	����&����b>V[�t��z�zT��%4����ң��K1�W��"�����1����%c� �
�{�#�S��RY������aSԸm�?��j�x���e�NKj�L��}��7l|�L���~rq=�jy��y��ºI cLW/�v�^����{���v�Kˢ�v1��Hf;��>�K7>����qcoވ�q�D-V����,,o�bueL!���7�v	����&,��j�)��v�����ȳ��0Jy�Ġ�ͥ�k�?̜d!�m�Vz�sJ����W^sj�H�/ӍJ WX���1���I���.Tu�s�w��ԃ/�p�-�*!�W�@���Xރ��^:w��B�շ@���AO���T8_WQ,LUhwW�f@կ��3*r��U��l�U��^}�[d	��h66��oӱ0G�Q�*�&dB4A9Lw_C%��r{��i�>�#��=}pY?�!�G�#q���
�As��[DSOw�}��!c�y���-��=���/L�j�ғrC7Ye�/�Q��`<XGe�J[`�R��Y,� �-`-_*����O@=�� ຫ\l�;1��G%~�TT���\���M�`CVk��#PސP�YOi����]*��7
�AhkG�����>�a&)i$9>x�ȩ���(�g�)�!���}�9���$�������˖�\��挾��-����Ԯ�t6�9��2�zp�D�^b�Oh�K�/՜�+��g,�sG�U+s�4��� ��{� �o���*�h���ac^{�l;��ce�a�]��;C (�P#؄���5;+���p�3���jɢp�������t�Z�o���1�������(8����q-:^G^�ϻ3}�(S��?�1�����&��Y2����#��bZX��o��Ekh>m8�:��3��^���C*����a]��_�Ɗ�*��. ���vw�]��-N�v)�b٣e�	��`�9����Pa�^\JJ��"aC��wx�M�x�u���; "~w����o�*̛�88���Ŗ#�:J��e�ٓǠU�����j����i���S�F*J��L�lUK�1b���xH��q����ݬw7)ȿ
����5�	���?�#���7�S'�Y�$��ajb���Z��b���7e��_KSk?�q��4z��
zK67��Zۍ��>�V��YyBX`��ߞՄ�yR)�QӤvl�De<j�n���!��I��n΃'�6�Jx�z]Y:&.D�Ճ�k����"3��#��Р��E}��8n������=��m�|�+��8Dw ^@��d(6p�~�Q��#����C.�ܿg��+���͍:�_��U�S����|'��Z	���0fr>\�c���g�+�IiJp�]=F��h���rL�.�V��SR2���/}s� e�26e��<4���'������ji������P����%:ݽ8ל�>J�sI��Ђ�_lu5��t
}?�VC��7*�&d��!�敡Jw�F�M�;���9����x�Y��<�\��<9F+0����-�g{��(z8���!��@���U�ݠ`~yGYo��C�K�ֹ(/�ܖ�Rޣ��/�uyj�He����"�����0f�8�1`?v*��ōb_R�OϑW���sb ߉ �Z�$���f̖���ydc�]:w4F;w�ܾ��J�R:جN1���{�rSv�_��5� �r�6�?r��P���/���*+d�K��b&��1����qAD��[ �37C��N
��Œ/@ �&X��R�xг�H��!����E��A�a��?��2Y�������T�텮�XM0�[�KC?ر��U(���`뛙az���cl�ݸ�Ǌ�[��ɡX���\�|��9�E4�̲#�8�]�_��N��6�����l�xl�N���ΖFԲRi{}���"4'~:����=1#�w���7˹�����#`�p�|/��5G����L�r��1�䎏�dn ~]�!��fw�ŵY��H�sp�m�j�D�KG�
�NT�W�Bͣ5k���ژ24����Z
�X��ī"�W�˼oX���p형�����u���7��2&l`�G�,j��_�@���E�Q�^ǧnlD�6�K"�a瘲�R����w�,a��n���{Rn���-�*�{�͑e��.�,g���Uh=�L���5�[���1�e�B��*4]�ߏ�����zj��.��Q�Ct�f�Ѐy��������X9����08�Va^Mu�&�Bz8!�Q�L�ߛ��|N^�d`��j���F�,"a��bsE5 ���"a�Q`o�����+Ҫq,Xc+�ܐ]��a��d��8�-�&}6G���6�u(�>�,���ݩ��<�4V��ӔbqL��9,�AQ/�������T��y�����I�:����{w�PN�6�S6dr����5���
4�����i�
On�	��[�kd���Iݘ뿪�.i�y�W��|ɔ��S��5�~��cR Wj^\g�pӨ��h�{ ���������(��������B�� ��t�h��d�֩"Al�>�)����H�D~�wk�:@H �e�����fq2,���Vй�\.X:��QF�ȩ�T�k7cJ׀�F$��Y)�Ï�v���$�4;��bi�>2 E��=S+պ�N\�zS�`H�b�Ix��:���`?����7r�����ۀ���pn�m��-�k�K4�(5�G�j'Ё�P7�C��64�2�Gn.�!l�jR��M@:���-O,4�3�@>!�\s��bmD�ST���2w�"��Ytd2>[f�Q-۱�bC�����YBR��"��|~f�'j�����Һ�X����jT|��ic��K7�^������T��o
D����8~V=��i�F�;�V}���E+���V$�jfy�h8�JW�9����*p�W�.�B���j�
_�Vp�X^`�XfQ�.y&:iO򖗸�;���e{��]�tU��*Qy[7:�ez�~u���#7[&��@�s۠����́UizLbX5�UE?�$('�`�Q$���So2�C��q)�yF:o��������lD�]FX���R�$�c�ft*P?��o��x�p$�C�8;���̦kGp�������	�̥�R���O��/���9�_�HC��9m�j���Y��a�X�l�Ȯ��U���G4�%�ǖ0uLbwkl�ps|�װ�;�)�����]��6n�V`ɝ�Q���6�J*d>�s��뻉k�rvu�Dot�  ���J�
�*���(��Bԟw�.���r��L�lPv��'0����T�����[k��\/[x������s2�}�X^�f�^�o)�?�.�㇁�7�t��D�p��Z��JzT΢s���gԗ҂�ĭ�>  �V�Ғ� �ԡ$��F�%J����xҾ} ��wk���U�c*��NWY�R����bL��j����CO?��0��O���H�)�� ��~�UD|aB�d�N�r˓�6��Li��u�u��X���.�8g."��H��R��X���a^��#{�Μ	�`�(��.��-u��*Қ�f�o|+�W/n��+��?��H���,^�2�x���p��PZ�ʨ[�qA{̪�$^M��fR Rbb�(��I��;ˋzP*u 4q�z8D���:��~:��I~cs��Z���u�Γ�rt�8v'a�83CWb�x9��@��<�����׋P\p}H2��)T�"�N�y*+�E�)?YP�`�euz����5@R8/[|78� 1K��+-|���RK_{
�r���7�W�����������5Y�����iL�����lv4hc�[���-�r�$�����Ns3[�^��Ahώ�0���m�o1��Inc0��[U�4��B��봹L:W�����O¼�o�=�>��n�Z�8���y��9���ؼ���01ŜY�zm�.�Q�����!�m��4~lïGs���~&����Kb� �+sĒ�����Y�KYVߴ��	���A�)�:����6����'�����tⷠ��"�G��Ռ��s`��狜k�E��T� e-IX4�@{�,��8�ᇏ �R��w�=����x@qx��(3�%'6u��z�l���
�m4�yO���kX��}<�8��I� ^��L�N���o<!� )Cm�D��ot�YO*����qh��h�;��1n�*XJtb�5즄��W�i2η�x�V"+�T7����{Sk;���S�ҦN�>�vV�{m���>��$�ݝ��:����h�̫F�u�^�ٸ.]���H������#E\�iQ�u���AFyJ�{ٰ���vx�w���uI����
�$�������)����^�<3 �"�L]@r��*��7�TJ���5l�ǜK�DɅy��o��(h��N��m3��AݮG�;*����!$J�ר{�R���!�V,yª��YBGQ��Y�Cٜ|_C��	��'2y|�b�䝼�Xi�[�O'S �QÑ5�=m���e��~TU�v�`s|�$;Z��%y������d�+ <��ȥ�Q��;��9\���e���2�pk�P�rڨT{�����Ŝ]�K�%��6�
��1��Q1�b����IK}Ȯ������Қų��C��Z���5����y��)��u��S�i���OO�`wd��i��]�8 Ƒ;�$1'��Xp�񠳏�Oyň���~o�A�!�24���L���9z�'��a�n�>�E=��Ko���ƨ��;�t����Ƿ�1ʄ�f��"��ω$/I�WM��+��N�+��.2�di�N0�7q�7������{��$������{Jo�O�T�hD��n�DQM.+�}�6�A��"1��X��ʖdY,vDq�Fyx��6��a8V?8�1k�&﹂�M���F:�g�7Q�DW�ʭ~Ӻ�:ZH_�.��3���3��!�E��
F�hD>��1B�㧕�m'�f�'s\=���|(\uA`A��� �
Y������-�0D�sy�|��RK1��>Z�Hg�w1ͦb�x7E�����'!q�Q���;/���[�E�;}-Kx,L����G�0�{��M��x�&o����9q����nל�	��@�P�L�|�m��z)��e�����}�_]������#p�S�_G�+3V\
9�Sҹ^�����>��ۙ\��]8�Q��N����X�x��k0��m�C�ׅ;�ř��Hm:�|��(�fE��G��q���X�P-� yI��G��h�������6V�)wz���@����"����Xl���;��J�y�W��笤�t�m,�ڂ���ˈq渪	����>.��0�f�Z���g�������  mx������N�zD��}-zX4LJ����"q�R��H��-��NՐ�cy�u�XW���Ûl[�u�lzM�﻿]c�Y��~��Q�V��sx�A���dk�JIYهk>���0��ė�n�U_q=�"����fV���5ݣ��#�Q�0���*z6i�q�h���[����_���0b��Vo�Pai鼳A\!M�hf{�{��Wrk��Gtb0e�EN�Γd��
�?���vy�' Ø}+c��r��4�G�i�۠�
���\�:���p��U�2�.^��#�������z��L5��B����:2��l5Ԣ�J��b uȾ�}��-�E"%��>"=��e�������N����z��O)_@Mot;��OT>�ڬ�>h�����/�}8t�v+VW�>��Z�c��ǏWto�WO	�h=옦�R��H x΁x���F9��ee����Q�����R��� 7��ZD%�ؕoF��t�	��~A7U�s���.w����b�'��b����Z�Jܒ!��}���vF��Jy�?R��$r�*�iBJ���4�6�&=���_���ND`R��!����xz���M�!�mn��[��R�..w-G?��%� ���`��r���	��6Ԇ�e3�YQ��C*�x{�2�s�0�f�����E�!zt�|O�� �%�"9�]���§n�9k�ö�ɣ[.�nvA�)��Iߎ'u���j5�͂�1Ԑ㴙ļ1uuhާ���Q���YM!�Z���Q}+�О	�\�l�KL�0���DT�<*��}jY����H�s��}S!��!���<����	����I��]D�^r� Q�DG���p k�{-�� l�e.L�x'�|���uР��E�#���QX^�L��n��|oKP@��Wx(P�-�$U���@��B2����`'��x1YmTG��@�x����7�!ϐ�)r#-{�^����i�Yf/��"���R�*�DF���1������xs��W��z���~"=�@��&e>��ŐL>h�rsߕ����E`cl8ή��ʷb��t`�U��&m �DR��	��c"�䖐٬�t���2��:9-�?g�J��M��<@��W����J��&���B��D5o��߮��x���X_CW��6>��w�6��8�v�;%��{
"q~I�*�H�O��*}4��n����ktO�ɢc�5�88I��$���t~kO4�S��Y!E1G\L��O��3׾��i�ه��geNZ�2Op~�򘚿]�B��I�`p��'�n�������Nx�R�nFϐ�qՖ,�)�������(&��䙎s�r�e.T��m\L�D��IXv���PL��gyX��K�e����њ@a<<*]�k��~<:t:׶tѫ ���q�
 ޽����x���Iɓ��$𖲪���e�vF�[V2Լ�5��ݠE�/l��#{��2�����QO�I�Qk��������<@t��9�aDN���MU����V� ��bO��@j]u<X����ińY�`�V@�2W�qJ����}�|(��<�`�r�8�p��H�b�n`��o6e��%�d�|(Q��DS ��Y���s	���0sՎ�+8�c6K�ܖ��?���b���-�J�H]���x�Nj{B"�k�ۨ����׫Gd�����2�c����lR��+G�2����,AK�U=�K��w�;xK�.$�%���ڋRU8y�3�'ʿ9���ܳ ������Bk�p��/w���]���/����}�(~hϫ�� $R�).����JpƯ���nt� �\?�.+�iC�B�X�vb]+�bc���z$G�QE��[����"HE �LY�U�%�Tp�1�"c��p���� ���$��_�oh./���o)�s�1]���1
�i�����~�`\�\�ZT5L�;o��W�]��o��TIC5p����ߝ�t�@���|$[�c�W\�_�m�V'�� sZ;��Ϻ�*3GUI0�����o��mX*��B���pЀ�S6}��Ul[	�9\C��Pk�p�;)�a���b��[�����L��p����yY���q���Z�w~Td
�ѹ*=8,m��ݒ���O'ӛ�}H5c#2�W7[�TH�Δ�s�`�-2�u ��^b�F��~��<I��%��jY���q�.~�H�1�1F+Ź�h.�J����~��D�Z/��
c�B���̫���¯�Fp��cA^�M���� ķ���͜W�}H������$8�*���z�(�l�a�E�xS%�Ӗ@f���=oY���t��5#H5����>T�g�LZ)�hG�53�L�f��)\�Ԕ�տen�q��'��V_l�%��Wh���h��ƺ��g���mOڸ`A\\��`�'��K����NH3��N.k�dH!��	��4�;����^����^�J�ۍk>Խp�0i�Y �=N�豖�lZ�$g<��0���ju�I�oA'_&�8�n�˹m
sҤg�x�}dXÛzx4�+ ��
ƱV:u�q��m���e4O{鍨8.˫��K�]1<�(�X���0�<g���ܷv�p�1�C�=���x�$�d��gSXB��e�Sn�w�'�|R��yf��e��� ��.(�$�TeĀٺ��J~��d���g1�W��29]�ˤ4�
��ө7P}]U'-U+�3�=U��P7[5�\N/��|����S�yS!���)t�9�Ɓ������
T(e|)�T�%�/��놏W�G �Ev7.[�G�PA�ml�2A�1�u����e�R!�P���.�o��TNԮH�+��#���\��7�	c�m�L�b�_�pa9�ܲ��,�ڧ���Y��"���0�i���^�-R��d�2�1���G��,��n9
͵�r����̄`E�)uʅr�OnS�Z@�U��":���?�!G�v����e*ʏ�VS�ӷ�1H5�o�LB��ZT����AA/~o��cWm5���q�w��T4}�8�����Г6M�WJK�+�Νo�Q�9�u�=d���[V��0[n��_"a�hm-Kθ���M(胭�bZσ�|X�1�/�HC�`�{���(pgG&��7�<b/���Ɍ��35#�� SL���73{�Y�2�'XJ"夷T�Tˆ/���C�:������fX��� Pہ��"������2v'��7��B�dT�+_�c���,����dش*s�(�������Fz~iug?,���z���>��������OU�MG�2��Md�� S|0����T"z;���EP��Ӡ�Rl��Up�:C�V�����gq�F9��s ��]��,Odظ��٠2J�>�:r_[�3Q����]�YgFm�W�hI˶�~w�X0�5Ro8��qP�S	��*_���@�ʅ���a���&$���¤��>A"��+�Ֆe
j�0�\�j�L��c�&�������Hֻ:��z�w�4�t���6��f�dy'~&�L)K>l.�:V�ll%��}"�u����1j��N������B�o ��Iri��t�w9�;��>s��[� |���`�Z�ǻ�(!�g(���1�&Cʪ�}���A�oZ�(�r�K�����(�~�;�VÛ9' qL�[�a���"�4 �T9bT��D'I|�x*�n�e�o:<�=Ok~��:�H)&J8�|㎺|�2p	��U�oQ�d�=��eKë{T�.�;
��P[���	FI�G_���U��� �D�%����Ɇ��P}qRe=�m���a�^>4O��D�g���5p%7�W���^z��p���@ހCj�c�&�UخL#���Ծv����Ӯ\$�G���_�����њ�)Y�"9L~S�p�V��gr���W�]3�5�8��۸X`3�ڼ!2�j����v�U�m��ɠ
ˈ��O��!�V���o��P�<Š�3@+�l	��[�k����T���@Diν5�y���@�r1,:#���A�� ���E��>��_M�?�� 3�@Jw5�;�X[��<阩�YfO��]��B
ulx���|Qm��h�L2>�T�?�F����{�WT9s�7� �X4>�N� ����Kz���[��ek���L���݅.���+i.��d����;���$�~���v��֣�'۸M*���6L���i�*j�%?���%�I�����6
ͦE�JV�^��_7>��ڢ�M�Y<��"�B��,:��"t�t����N�B���7h,y�So���2�ގؠ 0E�K/����>{�#��Z��O7ɸRs���R��N�4��.��ݢk���1�K!Y��v��i>� �c��Dy��K���T-�uz��rʺ��p�����>Y%D�el)x�;����B�tԿ�؝w}���M��jr�dڝ�WO8Y��.D��Y�1u
�����7x�;)GL���W� ,Y�-��I�h�f?O�����DͳWL�`�H�y�=��a�l/c�v�陥-L�z =nĶjk�Rs���g\J�j)�TY��|�މ�7'I��wR����k7�zE5�t� �O���#���ĺK��+Y����%�(��7F��{���Tfɑ>j��m�����q���י�zSø�NX�����dn���`��3V�F�� P� TN&5K�,��U����U�LYH�.'�U��g��j`k ?���`��@޳�����j#�v£�x���{1J�#Kg�A�Z���3��߮��(����J��
���!����0��6(�3�X�Y7�� �_��R���`�X^P:�%�~����Pe�j���\s��_L���3ɢ;���aQ�E�F�"K/;�Y�jA�I��ҵ�+�r���x�8IjsחJ�R�:6� M^���}x'vAC>�%Rώ�/>+;Kyn=ͣ�w��?���og����H$	�xs�@���K���a=�$���2�0� ��d�0=�N6��3�[_�^=��u��~a��S��W!�u0�w���*����)�piO���7�r�=d���N:��7i�P{�(l��8��8{b���\�	*�*��d�s�4�5��F��������.C�o��rLT%�K�q��?Ǜ�ɖ����0c���[�:>*�����,ʉcW0N���N�E.K�<N��j�q@\!�ً�~q"��!��:��j�ޔ����()�z�g��zK��gl�yv���ѧ�+jV�n=��;mrV��U�{��b�&/ �:�H���U��v<n<�	��1�.:���{�,+x#PO�������z���an���'����Ju �[(��d��$��ޖ�M1��\W��YטݒZ�&?�)��?��e�8����7˾N��nV�տ�V�e�(�_c�cݛ`�y�^�b�!M�1��u���@��2��E����t��nG�D��C�Yde���F}̜Ps�l��m-�l�Փ�-,z��γP�a�<�_�x�o���%aQ�q@h�C���V&	�m��mo�&���>oh�$J���_:5׉Tҭ.A	jنWgy?�-���6�@E������cu"$�D�L�Io�	8��w�:��s����ke��=����Nx�[:O��	�SK�n\&�)�賁	JS�2�+��F�m�%�*�[;�Za*��[[�gI�1��0���T�*��;�$%C��E'��qS'�`��ugF0x�rh�'N<��e��-�&�҄(�x xm� 7J�?�5�&@j�{���gI���S�L��ӾE�n�k̭�O��SDxk<6>��pT�p��G��߳�zQC0?4��3^�n�cl�~.Ƨ���I��Z�"�u���¡`j��Ѱn��vK�tF�`������UNy�Q����{�Pr?4�3h�e^�XDU@���$��77!�I�(���c���6����^g��u����$��ڪl,��M�$õ��6��u��0ѳD/B\��?��(^}W��e���$W��U�6a�T�c�q5{e �)��:�:�Dy(�u�Ҙ�|��*\�k^�~�&KT���< ��vc�_1�H��as#�/��Ros�=�~j�|���7���o�
�F!z�%�P���`� ��'�迍�QߛPe BYl\�1�J���͸�I�^� ϝ����o<��ȯ�y����z�)9YY�Z���rQn�|�_�μ��St�P����&��ZP��5�ۮԹoD���E���\� ?�TƁŗ:�j ���;:Eq���4`�s����hx������:v(=��Q"�M�wP<j'JĀ�߫e��S�Z�O�#[T�
Pj�g!W?�eKA�4���'�G��~o�O��t���V����ޅ>�NNtvl���Wٳ%x_ȵ��E'w�n�SD�lr���t�G��n+�v}�z^�~'LR|�__�R���c�{\�gd#W=˜�Y�6��Y�R�bj��T�}�S$������k��O��##�c9��_�hX��w|:&Ooҋ�3{�a�JT��c���ǽ���I�:SQ�"$�����J�*�N��V#�u��!�ނ:q�+�s��0
��m{"���b�z�c��<��)r��u��P���T�&xgk�s��BZD8�EQ�]�V$4W����V��T:%Z��a�%��*WI��O�3xA����
�b�޻N�<q�|O@ȩf����Ǹ_�t+"Ip��[���-�� �;U$�L%�
���Uq�Xϭ�g��C?f�)H32o�k���F�������t>�0X���!�J�,@l3qeB42�W���_GDK�87���5�
�����3��ϊ���ՀTc�u%XPĎ���L���df�U���5�Ss�#9"G�����i|�F�����~a ����w#D9��3����������ϊ6a����6ű?{��QG��;��#��=�!�x������a�N�ٺ��$���U��c1����2Hփ����)C�:?�KG��^��ԗ����W�Ú�v�B��S¡���k�����%4�3�����=�"�t����j���߽�J�`�m������X��Q맞�<z�?�q��Y�d�w��e�Lw�߹=��UA@@���7P����c��צ_�a0q�T=T��l�ܸ-��p;���E������w����x����l4����V,��'�{;���4V��s���SN���NkGÎY�-�k���R
~w�^�=6�,��CBvrQK��U�օSzJ
8�|�}���v8����m�T[ ̣ь��cY�+*�iU̝�[�^���i\*�����ܒ�
U�������-�Mx�^e3�)�oȋ 5UGnY!��� 燣6j��K($�̪�,,G�}����<�f�����t�@{8�3d�4>��͵�-�V��i��tiN�H�לajpj%��}�BGN%�r���y��7S1����l��/߁�?yƚj�P(t��0�h�Ӯ�K�|��vR�C�Hv��n:�H��r�� ���/�]& ӏ=�z�";�O�W����U��gN����+Gyq��j���-O1�I�X��N�kG�M��M�ꦮ<獑����1�7Cʑ5<��t���6�u5/��ǹ�1�r�&ob�gEծ�^����㾤?��O.���0L:�,�Х��ym��Ĝ����}Ti&�2����j�D���N{� ��R�b����~j5+t�y"�R5�%p���K- J������ڗ�'�b��T�(8?�L.��ѻ]�Rв�o�Q+w�:��Y����}���Q��k�SJI�{h��U�L,;���ak��$ED�;�>�I3�oЉ�l�3:N�A�7���R�L3��ڼc��n;�o�{M��-���q�L4���ȓ�*��骚�y;�o~O~o{ZC��wk�ٶ�AP�%�`	I�e��(`����y�J=K�C�.�ԗ�$MM4�=����;<rc�U��P$p��3�)(���䙼�M>��
�,}9M#=�7��Y����!���mx�Vʝ������?�C۪r5��O0���vm��2`�����S��Ţ��C\%����t��4˟6�m�a�	Q��
��w�FO��hj���Y0��uw���m��*P-�L��4�F_4nX�\�M@�o�O%\�D5xq�6�Ԣx�˴� q��N�5�iza_���������w�e�MsU������h,	�1��� ,*�r��y0��<������Z��>b?���*&R�����!����͓G�b�3�-�'f��T�#�YO����Ȃ��-|���"�8�t��b�Xm�CE�� n�vA��t'�EE�I�&��s$���ܱ��g\>?�Bgm!���k'lc���,����AKԵ_RT�G\�ʘ��NW�g;F�Fw0x�*,�Xϴ�j;�N8��6�iK1=��ba��j�X�����v'y�^�e3��=�G��&���R�ИB�H$<�)�k�3縩��[���Ó��,1�cG�:2��K#��$�dʁx��-��v��Z��&�Jk%�f��,$�PY��Õ`1Kw��	a���i
�F���S��]	�+e~�v�����7w���Z����E�n�β�+�y�@1kO��[!� ĉ�ꏉw%A���x �����٣D<́_�Ne�@';����5�5��+6=��/S�T�:��L�g{W����
t���,������ɒ3a( )��C!a�-d�|z=���aA)�=����k�\�+Iǧ���/��@O�����u�D޳kŮóZ�n�M��.�|!���
�y$a�W��f |ǟ�}+�O��a��-�e�edR���q���y���qR՞��6��
y�q��g�<u�b�(J�8B�e�Q�1�⧶���K�������%�:fm���A>�f�LF���y�s�g�a��^DA�Ж���ł0�!��qy�$�n/��]��]�ɝ*��"k����{I��#����̞���o$���t�ڛ%����F�Q�iv��V!�{�>��uR�������=��h_#
�KݱDv_t~K�w9�e��֋?5��<"�:M$����+�UXL�3�ʉ��v�8=2Usc��Ϫg�Oh��(}O�!�3Tz��A�@0����"Qt&^���0�i��s�T����C��k���f>�>2�I�)�ǃgk�{?�hkx����25�$ZuK�ׯELv'��'S���4����Or'Υ�:��*!������w�a������n�c�Q��kT�}zG�� nn*�c�k]����i�>:h����6I�L
i�`�* ���ն�#�"�>H�"��{��]2�����EP{�^�Q������D�;yg5=]��쒹\�GvI�&4����.4S���v��0J�WE���>)�
>��+���>�e��uXw���	��:�`���-�VY�jh�-�����&st4�f=R'1��4KY�F0� \�0S��>S-|g��	p�F�al��:m(�]R���j�TC�جڙL*�xdbŹ��� � �qb�PЬ�n1�gJ%�	,:���`�C}��4�aH�TQU|#k:�\1l��5��� IK��� �v�%�P�jIU���"�n]g�U����%��q
[����bx)�eP�O�ײ�i���1�yu�ŵ>��0kv�JҾ$��$�ݞ��`��g���W*���5�k1�g�Z_:��8�̢tB]C�ѕx��h�>��l]�Ҁ��������)���D��������[9�EI-x�c�?����*%�ߑ$3�=9iD�YH#(ѡ)�`qKR��i%��]��B�u��d��k��6�*�g����f��2��T�.Z ��_.��9��W��sgd�J�쥬����0�3�x�6�[
;��[����TH���.����mP�)`��������t&7���`BG�\��呛���P��^�S��
� ��ܵ��X3l�+�},�'/�w�r��?+�6���AdXm��gn��CQ���5�K5��Z�4��(8�9Y1�v��$b.���-���<cg��-[�v0q�ι��o{���|r2ܮ���R2�x�մ�Ȩi������i�P�����43j�� A���iY����c�'.�9oL0��D!"�a��m��[.c� ���{���s±��:ɗe�x���W;�sɳ�䟪mf��E/�X����pf�.l��^x�>Aut��8��:�͋I�Ã|C䠥8k���{썬]eJ���3^õ��)���{�EdDgY��2�G,�� CGL�M��`�>�i �b=�Uku���\93��2i�iUf��Ώ�P�,
�/�W����ל�Z���c��ޠ؍I/�K[�8!�� ����vAֿǧH`�W��i �V�v`d8Sq�v��=0J:\ٮS-z�6�1�z ����R�t���H�Y��4t�1vU�I:�r�j�C���z�I�<'�8AN؈��YPȥ����'�39���G�C|8J����ܞ���tD��D^�o�J����`�J �Y(�<M�	h)�=<��S��@���L�S�v�!;��!��}��[��������T��|>u�t}�zn�h�;������棽!Q�) �����0���=]*sr��C�o��}�����L��z�W�q1��n�l�*���ȕ���a2
�#�;��@U>	hGq�2�w��s�t���Tx�\Q*�4+ַ���%5���� Sa�GϿ�)L�����b9��w�{q�;˭��|���̨:�\t H*MI�A������hC�%dY��� W?��F����d!'<��#4��{A6���~3����SmB���ո)�%�ȍ�<'\�h
��f���˄ڶ7�\3z���s,�B���H���Ɵ������:�Ѥ�/	��/�D������/�8*J�@���eN�E;�47�42���k�:N���,_�L6]r������xu���.Ds6a�u�O&�`��-�!��r�D�)LmG9���$��x=m��f�B9��O����>At7���{H��+�)i�R�C��D�7��{��Ir�Ş*c_��L{c�_'��B�"�^2ls�h�`��`	�t$�����_�!2�q�k��� ������6���#��t�̡�_0�4%��dN�P` Ә����H�3�KM0b8�t2�ꄘ�[43��Ȼs�����1�_�s@*�?erxx�6�;�;�!�X� �0�R��A�����|3�)���g^�_"<&pyBp��_�|��5��U�*��=�6EI�pL6��?i=m�!�n���U�}׷��o�%e77K���ӛ��q�O񑷤�W�Ԣ`N��ϵy�,�8-UeA7�����)]q�#�6xv�a
u�=o��	�7�Ȱτ�>���2�2��a��������>^Ճ, ��w 	�'�L6kXNDO��S�#`s\�,�Y$ߓ�I�?�|
.��XX��5�z�g�#�20���b?߸��@���:�d/9�\V������������ٳ!�|�A�Gn������Q����
 ��>�5HgYZ�6�y=�،�9�u
��n�'���)7-F�}�\��}g0� )t�#���%w�?��˫0�2��n?��0Q�����bJ�E���2�~%wC��d��8�ܚ�iI���
녬z�e��ḱpi!Q���B�l~Ë�03���Fi�p!{Fȸ'�/��"��A/��V}aqg�"苙9-y�%j��
��Cj�DvPY��%�5�����f2"H�A�\ƣ�'B����8*S��,n�U�,�ȼ�=�	B��x�0U�_�F��2	�M/T7�����i6�±����D�Z�]7�p��Q�h�t���'*�cpܹN'J��J�}����٦*d<`���V��/��?����0ټp 4)�xn?��}�m-WC�쏛��O�������q�y���g��c�j��?P=�F�g4T�'��;��I�a�M���J����]D˱�]�L�"��_IlP�0/���X��!NS`0�,��v0�\ ��|�?�|u�����i��:���*&��,I���\���fRjq�T�ܜ�����uv���W������zj�ԥ��;"���{�T&�#��]��ƴ�ی���
�1�F��~�7�Sf;�+��������٥Y�"F��c�A�uo�� ��(��L0��:�R��Lz��H���ʃQbSu��eG��5�>	��쭏�n�U��SVߋ�����U�)������;���B�/�S�4"������E")w9=U��*�iu�vk�Ʋ9V�::"[�<(��+���W�IG�.�sS��.�9�.��(������a�@~����C�u����X�肥׿�a�L*m�}U��$��mX�%�id9S�!Goh�p��z�ׁ�2���@(:��7k�{��
{��I��9��'���шp�,(?j!� ��/�����u�����q�ܭA�-��<dYvO1b���һRN��']z�+��wh0^"�q5p��^�Y[�@���<^�4~���i��a}��
� ��փ�bI`����}�w�v�V����
��
�y/�riSt������;�� �(�?���U��m�(�L���4Qd2YC�a�rO"���rUyѵ���MhY��0�ʅΔ�f�@%�8&OW�}
��B���x]���=H$_�ɐ_G1Y�`�d"�9�V7m����D�î�q#���s\%)0�4dd��I2�-C�����?R�8ɦ���p�=mED��/M'�����i`�"-X�v��34G|�iJ1d�Ƿ��q�G�H[ژ��<J��8̵ j�
��`q�ӽ����i�T|��t١f^Q��!R#+)�M]��x�>��tB���6k������YG�����;c:=��χ�x~N��]�"���_e"�dB@��>��Ѥ�g�Ǥ �F�e<�/�Z�� �y0f�7�-�M�D�k;}RP2�*P�w��Z�ѥCz��b����&����!LA���b��</ߴUw��o40ܩ�fR�H�/c���+a8�j�&�=;�?b�4Ѝ��
�bt8����A��-I$N�n��Π[G(=�P%6-QsK�𿅓N�8�bL�c��?2l⻬ �g��G�Ɂ?x8��5%��d:v��gՆU��M�S�E�B�v�?϶ �N$���yi��jϚw����$�9S_?X����Q0�;�Y�c �7�͇�JJ�Mj�ԣ�<���O�o���޸�e�t:�`fzʁp��Zt|EX+��Vp ���1Q�3�
[�Pn�[���%y]"��V�ӌ�ǔ{���ٹC��,��D�F��������>-�o�a
�߂ő��Z��#��オ\��@��0���\�C��(o�<vK��c���X�T�cM�AI�
�&h�|�V��~X�6��vZd��7�9�����$�屇�{�­'A�yg���8�ʹ�b�Œ�x&�����v�ɡ�k��n�,�Ӧ���0OoQ�˛T��_�uiI��Nx��yz��̋���Ĵ��r�ы�������WyhW�5�� 2=�i����:��k۽^�L�@�(O�k�a>&��?S͌w�)�d��B��'m�gu��]��j4�vv�O�zi!���k�$:�	@��ERq>�ߓ;��� 協�^�o���A�'��W�kʮ�H1(�d���ܚ����u�7�8�x(l?u�W�#?�Ԡm��@�X�kc:�p����g����������:��
�Xuzu�T�o�W�Z>8���-��� �C�x��0Έv��ď�:���*�A)�i@�~�l���GLV�!ǥ���ڶB���͟ A2�ō�S��cl��/_"<f B��ᩐ+���_���c���pB��Z'���%��ӆ�ۭJ��Wh�vU}m�x�ZO��i��UfG�S<�kvr���8���+}� 3���%��m3\B�i��E�lTI Kk#j8�))�7�^�I\Q���:[���	����Dh<୒y�n���@9�����B����)B���{����
��T�y������s�(nl�� y����D	g��Г���=��5�X�i����Z
���1�l�&�������g1~X����f
V� �fN&$>\Q;�1�g���k�,�A��邽��9�Gؾbƨ8��q��[�u���Lh�3b� dP��9�	S���3�,/nC��h���M�U������q��s��r�f��h'��6�ZIod��ݗM�.�*u�^i��KY��2���}Q�����j��bJ�~��Ӄm��Iyo�Aq��ꪂ��y������L���𕛌R����N�%6vYш�*a�լR�O.��2�����?i��ii�0g�� L��r��ؙ��z/�j<1�	1��]�JyJJ��..�w�0���.�#nFd��>@s	~�Sʿ+�^;;��
b�w�rD���p*��ù����m"���u@����}҃o�^Co�V����.ێ��8��IP�iƪ=��2:'�f)(�Eޤg��h̿�8�@�ϓ�{�L��Jo�(p`s���h59]@o�N#�	W+1���T�\m�����Ѫ=�brd6��EÓj�-���wNP7��:m�K�{�X�,��Z*X�!�7�MWf� �AŮ[P��X�B�E�P��2`�����:)>��:�\zqf�Oߥsm����	���ʖk�l�������q�G����9Xc�*�aF�� fVxp kw2l��f�g`��ة�os4'c�ͽ+�U�9�"/��~�Y����7z��f@�r��Ӷ-�ó���O&O5��l�kR��E�>��J/�1r��)|)�ӡHj�8�2k��rR��T��O],ND�'�k�����ӫ�2�d�]G��<�����Ϸ��{��ÛQ5�ȋ�羁h�-���F���_�H�?�*���اֿ�crҦm�o��HHT�C�Ho�Ff�u�% N�6
�4�/KuZ�ފ��r+ �I6�
Y�N����ۉ�VK���1\�n����R��.|u�Gɡ�}F1	:�Սx����1��
�z�_a������-�
1���6�X9��*`Ӊ/�4�!ﰺ ��d�����	��|�hP&7�����[�l��{�3S�:%�H����M�.��}ʰFR�}>P���>��r��0���
�PX_���5�W��sSb���I�wE/J@:o��~f�����M�ú�f�嵣_-"����Du<����r$(P�>c�@�k�k�%6�J�H�� ��3�����+v�-�I�=��3�`z���ޭ�˥~�����
82�C.;��G��!��.ɦ|����q�ٸ�j�~k�L-� B�����K
bTQ�ܳ;lE@��������E�Řg��A�k��;��o�b��{-uI�+80�4�yC�oh%�?+����7Th2�ewOޛ85��4�*1ʀ;��V�y�� h�*4V2��,њY�)�TDЁ��æY3��G�'_���Q�v�f;��5/D\K4t�pK�f�4�NM$�F7���P
	��Ĝ���XE���a�Z�N����է� ����ˌ4_���*$};�p�_���?z�^�KW�LM��j�)���L��y�^ᾊ
�K<��>.Q8,p�CS��N� g9Q>ˢ>�A���v_�ת�5k�2�]��b^�~	@�[�$G⌃���?"$&\���A.�5��31 fQ�V����W�L� �Y]�"#���M*�'yx'�/{E�������J�_`�t'�M֦��<�|�H�1��o�"O�_��ԋ�%��jc�v������$rc���?�UDG�_5`A�-V}��/�팤��>ߒ����9��Hu��Eֱ7��V�-��� 5���������b� ���`���2y�:o�����G� �9�~o��tA�����0���e��Pq�a����#���o�]�U�P��^G��P�ئ���#8�ȿ�A҃��
�XqH��Og��h9�Pm��5�9�G
q���4�����4@J�Dln�B�h� K�TaB�44_I+LV�S���Zd�a�%R�f(�\���N�fN���=�ZP�NcdN�'ٛ�c��GE�nq��_P@�4]O>׸�[Hjx�>/e6�r��i$X�����֦ �a�ڹ��M?��B$�����kX�}�.8L�ѹ=��[�JI�s_m�k��y01 4���ҩ��-8�e@^SJA��M}�D�S����V`����(�툓ԝ���.i�|ȇz�.#8��eU��Bᭊ�&
.֣���z�x��hM�QP�<^����q�[�$��ءeB)�'�)a����r�ϟ>VJ����!}�X�bD�H���:�����"'֥7�b{۞��H\y�:� 3�y�͉��ӈVg��U��k���`JVIj��P���A���;�xq#B���<ɿ�X �
!��w$���Hزض��w'�Zi�&�:����:;��3�S@��h�o�~��9��ާ"U�F�8:��`���yQ^��~7C�-����ŭ��:j�q���7�I���X �}�B�5�?�gn�$l�y&�sPP��U���i��gjj�6{��s��ܜ���=ePi�$���l��Z���?�L΍�H�S�3EW*�N���h��Ϣ�{b}����s8��y��#�����<u��6ES�_�4'�uؔ60$�g���j��@+Ʈ��7u�10ɒя��L�-�S�FC�w%(��#!L;���y��зѷ�}3��� ��aE�!�k���{�R�wQ%��n�&
������E0��IRu����wx�Fu�9y���i�?�ђ�h�Y��v����ƙA��52�'�b}=K��3Z���m\^��򜊟|���	���Ӳ���>NU��ĉwd����"
�~�ъu�F�7��j��"h����uYha��q���C��w��\����w�_�
�,v��^���Y�0�u���5�`��i�L����e�C|��J��+E�����nu�E��ݪ�w���Yͱ�*������0�9c����=Ap�:i�9$�g@��W�>~��Wy�q���>��^�P^���ӼK����rQϻ#p���t��y9�&��ͩC�\2m���z<*�z�W��DI$(%BCL�ے:����%��(>�h���V�Y�Uzw��=U~٨��Fk�>\��T�{�>�'��dP�8��$��/��`g=�d}�;冑��#��O�e~U|F����O')]����V��>9e�6Nd��"|���eϷ�҆0Ki����kY8�@�p~oJ�������m��_W�����<.�wr�L� +<���'��������G,�n3O����G ��\�}�D�l6W'CWS(�C�!ㄯb ?	J$�9���K�������;����I�#����\�o����[� �Y`�� *1�0�1	P�=���XK_z��� �[ؾox�P���ErWC�!�D�/;���x{�h/�cUf|�Q.����|�~7`/��\LN���z[P*��~���:��S���˸<rYAPcv�PT�)��WTn�b�LFI�'��K
�w{���q}���*�dS')Юx�4���ҸatO,]	�|l��1XU�Y�{�&`��Pp�Ef	\RdE�G������H��]^$1!��<4�~`7@떖{9����o�̙�C|�+�/�Q��y�	�L֣ʊg�#:�F�T-�#�R�ic"�g���>+���a��b*ڽ�'��t��Z>Z��e�m2�D+R�-d#>\��������/H��RF����U��X�Dyl�IT��F�X����F�};��#�~�9s*36a3HRv��d�A3�s\-,2�[�Y�Iڷ ���! )����*zٚ��o���Sm4)Ϯ�~��8�_G=��� ����5Y��g��6�Xs�iSNUp+��w��Q~Ii4a���B�r;�<0	�TD�"\_�N~Y����n���R{Ɩ�� �@T1�ה#�6o�&�Q�s���V�3:�<��i{o� �C:� �6���i����R�e;�J�,Q$�B(�oY�0^55�h�
�#��Ϋ�RU7'�Tyz���)��)�g �芋�Ǩ���(<pV��܄\������ܐ�w�����b-�2��M�>����3�Ɯ�л��Y�{��V�ןlu���~\�N�2�+P�ː �� ��I��}.o�F^�^v>.�8���&4q�dz����L-un+2|`jY䴅>-�-�,�J#��=~sې�3����%�7Nu�M�սq��I�\�>_ր�]/�O꿕g����:���ǙQ�#F"]]��f,��~2l�F'ϘsU��R&4��A>�Tg��k8J��2��1"��������[��]�Tk�G���*����V��ǒy����Vs!�R𔈒�O��D�>srh�#��O�?Ko��*a^¿XBX���K�O��U.I�v��ujL���D3<_��җ���8�����Om^�h�i?u�H+b��:?�ڭ(ߞ�<�#�u.h�l����K{�-/h����atx�D�@���[��;���`dleɸ��!�e���!o�-�%!7���h03�1)?c!�>�И�$��~��s�c���n>QՐ���ݓ��m��6W-���}xr�ŗ{<�����ȆT,6mL�C�)��
,�Rx���f�
ğh�����*�����������.(,�\#���^�X�\촀��L��O}4@����B�D%x���а���Y��E=�V[s��)��V�M��.ٱC�we���:��߭��U���E��+*��{��8M�!�����k�`5^��H���E	�Y �jo�����N�ǐ��2q������ q��nfֿ3;4�C�]�f89�-�@�x�0M�SZi��.˅!.�}l����覲A�����Ng�a�3�N��}z�S�<N��]��s�����}�T�@�І����U�l��^���wcoV2I�������"A��	�J���V_���|�	<*��!a�����V?L�~DkU��cB�BLV� �~k8+߯|��'��qˍeC��!s�(�a�kN����U��)��ɵtq) @��	���`m|��	õ$؂����B!m7!��[V�¾����t@�##���J���ҋ̴PU����|aیM���ag7F�|�v���nA.bg�+�Ob�Ώ�r���d���G��_�J
�^���
ކ��N����;�k체�x�뙦�S�L��l�D��d�.c�J�%�v��}�U�y�6��u|�kFka�*��܉]��b�[鸢��@�k��##���m����p�-Cו39 |m�z98�ݶd�G[�@���5��#���N&f�_��-3h-�-�P�/�o�"B8vn�L�{�]�1¤�^C�.x��� VӞ�I��m�A?p�>���ϲ�|!��o�wпH��vD�7K����9:pNF,��S9�C���A����q7FQ��l�^�^���<��(�t�k�%.�!�"�H�I�N�6�?M���F�F.����N�A�0�v���T�K�&
���y����[�(Q�zxd�NM��yѮ��g6z��U)�س �YgXe�?�/�k"�1���ar9@��	�@6g+����#�l����R�{`�+^G��R��R �^0澫Z�ౙ��9]*��<_׬d�*����+�[��k�hH�9�k��\)��u��������&	����WT$X�:( �����&����C���^|.�-�6�n�C�KHW�U����Zу�̝��A{�����R�����8�#�Z!4���(��K�4�=�\	�MЕ�<b�M�9���)6r�	D��1?�|�~�H��^C
�1���H�߰;��>*W�<�hcO�ʟ��>á��b�����c���ȞQ�c�K�f����ZG���v��`\�y|,,�]r�N�|���� ���n�E
�g�X�*~-q�Cy�E�=�A�巌8X,w��a����bfN컜A�\h*V�+�+j���������^�@${yt��5���cLpCI�ě<Rܘը��'@�
��52��=uCːlg�v�	���#'���;�zA:��=b~t7"v��P������ݝ��T�cW��
����w��$v�}S|�c�>j,���u�kLO�vSن��B�^!��Db�/�[ʿ�LM�v:���p�������p8V�U�`ޒ5pVK"�!���^_Ϸ���o��z!�����[I4g�T�����aS{�?��!mDL\���5(Ԃ��AO�PX��#Ł��i[�l='��d/^Ctf��T�DO��<9K1�È4�i����L�0�rD�)"���틴
�Jv��_W���$)9J��� '�$���H��6�\`c����oP�Ѣ��88H�� t��Ucj/n����n/����&�-��C���6�`�?���{1�&%3�Xۖ(�7_V��޾;:hsz�0G~���C<M��0A$Z�l<Jv:2/㿳�Β�}�9�T�D�/Ho��j��|�;�`͍�X"�����S O�!3�M����������.n�B9���p<l�Ts3���T!ЮQ"��x����ӥ{���^+0?	wA�7_����o>N�`�R�{&?����
OR�4�'�}���'�0��PW�^�`J���̫OJ��T���Mkzkl�mω*�V8��h�ec6�7�޺�������C�,n���E�p��nqL������	~d�Q��$g���}��Hީ�56�Җվ��0Z4�5�;k�MF
�� v�������ΌlE�Ea�D��V死F������|�7��a7kQ�w>��!bc�����棳'ˬ+�A�ls��o���*.^2D�;Օ��Ð�s�4���~�F�R#���z�"=�-_F��IW��j������� ,:*�mQD\\=`I�I�'�3�ft�
�5.���m?1��Zަ�g�C���v�ɉC��
Һ�<Ǻ`����͆��W���ű>8�&�9���9��҇�����^i�n@��/ea�|}�Z\8�T�4�>�z�3����+�y2L�{��q�=[rbI������U̪�^e�5����|�?�S��#N܆$��gV����v�bC��lrF���5�뒑���γ<���5n�b�5��=���',��d����A7�"^қ��Vu�n�p����g{��YK�$'��T?�PO'��~F�Q���>6d��P��@%N0�̫z��e�I�֙�L���n��܏L�7,I����$/�c�4�`7{����4tr�]:lAޘ�032.N�mcsZ�Nv�����!Cr2�礊����^XS�W��\+Za}�d,6��3�p�5���p
�wP�0��b�A�/�"�V,�$�Rs���J:(�+��ş�-bF\�|�-&jP}CP�:�@�/d���Nr9�F,l�"�ގT� �mc�"��Y��>����-C�m��=�{�w��xK�P�c9I�gc��sq����̩�X�՞Z�[nl�	r���\���n1p�qȒ��Rx�r�?M�½~�iA��2q;d7%��ay���1CH5&����lٓ��H�bة��̪���gD@�M�aN}���iWȳ�1�X��C�!�ɷ�e�����L��E
�ҋ�Q��_����03]Y��U����'ao���g��$uEB���#��4b~}4g!�պpNҁ��W�*S��T��O�<�YQ,��F�q\����2�Uc�)��A�+ک�ޯ���ݝ!�:�6�|���I�Zw�����֋�A����Ra?v�8ɱ��0��/����xh���WÉ�]�M��%���PTVN^?�Vp1���t�;*H�>}�$G�k��9N���h~��D	��2B����g��w�K���"���i�(r�;�~�F�s��Z��g�0��<і���Ob��V�Or�[�;G�v�_�s�L!_cI�2W?�����el��ӄ"�)��{]���&����J4$�@��}*݌n%.WE�k\^�|fhm6U�V�KK��J���
hQ_����>'x�f�(�I��X�G9� ~��R�-?�#4�_�8xI��ju�5���O�$5_���0����A=v#U�̹�?9�x�2��h��iv��dXu�XE{����w6y.�?����]|jT��N��N�uު̴��h�%�cb��̖��iS�DZ�Έ �7sc<�
8E#���A�f����f��:��Qa��j�)@n=�uO�<��N�ʯ���feqG��2��s���t{B|[��D���$�0g6��}հ.�jL9c* �"���:5�z��qpI��3�K�RM
A��[q$��^��?p��ϒ(��=��i�os�H᜷&`ɅWM�]	�8��>%U#�]o�$���]"ć$�)�K���Lc�6���e�@� 7��7P���#֏U���ݜ��	�ru
k��~_Ϛq!��ae�N��ӿ��H�AW�������N^cUs���X�9C�Yϒ��W��qپ�$�A?���n����ԥzf�L���5R������$�_h����}�c�ԙN�Z�7��n��'�e�j�C�ɢM�x9���IJZ��{���3�|�|P v�C���Դ�ACl���^1�2�2 �XX�c��g���Y�첱�rq@�yx�����!���X�����V︬�H���	v@S�smtɨ��Oq=x�p�aI�9�n�:���\kJ����(�t�3���"���զh�{�]� "���@��8f�Y�c<X^�dY�A�Qx�G�0�4�q*S܍�Ĉp�t8�Ъݝ�w1e�-bZ� �*TU�&�HwT���.qߥ�ӅƬ�,�r9B�V�OPm�@(Z@C��i����R�jx��-Mj1��zf��]ǻ��{}��n��+N�i�X[_u"ހ9 ^۹���I�����2�[��n�̎��Z�Y������n�G��Tp
!�GPEU{��(�_yad�1��K�TU�������@{_H6����Uqe���}p8k;�+�@F]��!6��l�)1���]j����AH� ��*���~`����¡̴Վ6�y�����hy2+�}�\����2򐪃�b��P� YU�\|�/3��p4�����X�7�/N,z�ˮ���A|�z��eF���+U�A5�5l�v�q��I~}��H�t�*�8v�����{�����9⮣X�QrJ�nL��F��I��Bݚr�dU��]�8X�Ao���$���ƴ+j��I����07wx¿���T�Zf�E�LR3������C��t�~�^1�m�ś�_��-"@�7j����4x<p�|�9ۤ����~l����Z�2����y�޹q5F�9Z�0�\����w������d �hQhO�2�H�y�$K��}O������.DBoR���_f���pȾ��H��X���V/�"��	�C�};��_�*����,�m�1��=p��s�IG���8�~�mJ�a��ǡ�g~�:*�F;-ݴ+���A1�⫛��w;;�Յ�<�L��,=_��䅫	9hOܚ�%�7�/�E�,��������Lԩ-_��B�������T %���L�������?���&�J�{8�k�4��{dy�w0���ݰ ���Z6$��s�`[2>8�rr�1��r� a>^��,�}i>����\:����M> �FGML���4J��;��F&�u�9ad�[��������z3� �qQPuL���3��N��q�G�&;�򔩌[����	�w�k�ۭ����,���O������y�u���z��<������W���g�'��]*���!�[�ן|��=�7�d�>���8u��������kR���Lj*�#�[��+ݓ?���Ly9_�bŨh�%Z�q�]o��]��ޘZc���7.B�yu�c�8W���k�X��Cp�ް���sv�\|���Hb"�IX�A3ȎȝD�d����N�ؿ�Cu�Oc�x�IX�����{����[p6���������e*s~�� �'��:u����X�P����
��B����׻��ļ��2��؀���c���[G������m�ɴ�K+8e^�g�|V��Yl�Di5�]�d��;�5�Ez��WFzLv��"��}�X�'�<w�xnw�Z�Kx,	��(a���+4LR�ѺE�C�г4���U��� �l%8nт�6�2�J�'Q� �%Sĺc�T�`"�l�)z�������D@�~��wnǃ=������꺥��=�ġ!�됋VT)Y�Hv&Ӵ�?�젃]pD�z�P� "΀X�"ͭ^�g.�?z������l�����q$���T8��b�B����~�'�w��~-����^����t]��ׯs��(�CCT�e���%ԁ�~����a"�85Z�֎~��{���k�g�'�6PXP*�Ҭ�[�5�q�2Qrs7Q��_n��,Jt�/O�Z8����*���u[������G{�x8�q��)�y6�J��w�|���y�2�iJ]jF�_4�x�숯�����7�ϯ���ެ��4��-Bn������%��G~^��0��B?,�R���ʨqw���
�c�������6�.U��w�����{��n!*�q�v�S����3j"��DC�ͽEDe���g6�;/������;��Tr��	��o\1�Kҙ��H��W&\�`��!������;i�U������{�e�t�E�U�E�Y�����4�!j��;�@��|�/�m5��P�L:�Z*]�u���"˲#����L�B��	^�q�OR1ᣥ��ġU�|�U.C9��g�`Ɏ�f�:�_?�t:P��U�O�"�������[/���Q�yXH|�e��X4 �,D.���
���更������J�wQ,�8�3���JVsL��0�N��M������Q��S/��1�$��%��"���[ ���3ۯrv��H,/5�y��H`��U+B���Ow?�Է�3w��d�J�w�H�C- ����G���V◐qV��0x"�^p��Ym������K�~ڞe���r���p��v�gBS#�����wR0Iiū)��YvF^ί>�q`��xT/�)"?kk�Sf.�fa#W%0H,�ʋt��Y�=A��c�BY _����xՁQZɢ��i@nO�o����NT�CJ�s�[l�������~�r����U�c�yo}��#�/ �0�@�̽�������i��B�R�z+c��4ѩ�WIКE����R��mRU��3Ǡ���݀��}	/��8�2)�C�_N~x��	�������ش��ƥϞHXYh�naKx����=�_4Z�Z����nѹ|CG�2K�0���� j�e�j8����U��m�d��8sFض��QT�E	` V�ч�l��p;���g��jE*��R"80/}�P�������iK����kf�Ҟ�JPR�U �vZ�h����"�!�wf��d�Ղ�ǵ�ui���<˒V��fO��������p���ؓ��VGH!�����>�E� 8S��vn�yw���v�P<,J��5_��ס��5���o�#�����-�n�
�Z��OO�j�O���\:;���x$sp�:�<]�A1�&�#���/9��W(�zf$��V�fJg#�yUNf<`�1%I%S3�:8}��A��[!����'�Y!�B���%��$�L�e�nZ�n�-i���L�}�>��\���&�v4�k]s7שgY�9撱@ꧺ�eؐ]�?���2]��~���ɦE���r%�UG������2Z��]K�+�;ƽ*��:�~6��F�=:yq(�?P��W��；rT�s2�D)W�����s0RA�0��Q7����=�Y+�.5��X�q��[���i�G^���Lk��� �E��J�|�Z/':��rr�i�������A�(rn���`���I�u��� ���f̗C�M��kɨ���6�)�C�F�:�ush�
��G}�%��ŷ=m�s)nV��܆g-�/+Ap�.}�2�/�����=�d��)	�t��K����E�)ZzU�5�@�/��8)����\�|~�u�{� U��n�:�|Q���$>�{�ڪ��ʏ-�o6$`�Һ��HF8�ɮ����f��:��>�X�@����M�Aq�T�_�o��[XH��EX׌PIFƴ�.OvbM��Y�gE�gk�l��,i�eq�`�m<�"�Z�	��̩�M%�+�z�����y�6:�l�oΡR�H�����%��ځ+�$Zq�k�<�:ʆdB�кDm��ܴ�|ͦ=��D��z0�Hz�bZ�.����1{��[l�$�i�U�
;�ʤ�)	�ՌGB�
%^!��n����է�u�PaV��_�pj�`�Ćth��s&䄑��#�2q�b�т/X��7��h1���Xy?0�� KF�\På�|�y�zם4�x���f����9��IW��q�"7ƼBU�'�`�=�}��-�r3O�yXG��+]/C6����b�>�.��D7נ<��W9��q�@�4��+_AzT��]�A���gE�i�Q�i�OhF�I��7' ���i��)�I�n�>�c�'��:Wy{֒
�ҳ"j%�\ �����t��!y/fE��`>��]#I$���>�����Dg�:.qK�EC�x�Z�D��t����|���"�`fV���;��5��bլ|��H���
	u3^y���F ?e�!S�����vg8���H�g\�`�𨴀�O�������W����x �b��GY�&���j2�%��$���`�l�\P�Im�4ll�UXٝ�gzC��.j%n4�ߎqۂy.9�',.8r*
(��OEM��G�A>y��gP�y"R��H�`7��b�ǧ�U��Ȯ���e"�e_��.��]�a�ܔ'�Q0�P�wo��u�Ei!i�7����!LQZ2/�'{q��$$�,e��N��[��4;�~�P��hH���+�Gz[�y��Ƈj զ9�ڇ��U�V���vOLl�\�����ch'��;�#a�.K��V�5�{H��2$G~����K�!(ܡ���nO�%�c�>45E���:���*I�v�OiT�g܌�h'�e�w��+�z@h"`��B��Xz��y��V���1��b�h6�3���h�,Y���h�A��<�<�/������Sؙ$3S�I�
!�َy�'!�=���S˹R@��f����=XAʾe]�]�Y+��Ԃ�J8��?ME�&�I�5��LT7�Q�d���(Z��7!��-N�vG&��7�w8��������8�o6M�.�z~�0�� t�~E~���Q<�E�Lۏ<���+�\⍤q��Q�#;�9Vk�V4��~/r1J1�PmE$_UR~���� �]���p4��&T�+�v��h��q$��| ���xځ����=l���|���_�xT?�Wj�y]�M��42�;2����+��ޒ&v���X�Z�����:O�6fȒ|��H�<zx̶�K�9ƶ�Cx6 � "X'��9�]@�t�>ۑ{}9�=N��a>��	���Í��ĈCi�p:qh��1N �,��r�8�?h��9uc���Nm#��e9�9�b�.�5��h��:�_�gŮ뇧"�SAۊ *��5�Bl���?���M������6�݌�L�w)椬���zӿʱx.�L��S���Oh�������k��~���ڈ �CPu���^��-4� _e$Dg20ƑW������(�f�v� xb��v�̿O��O��8<������l0�M(�}v��*������%�zJjڋs)�?�j��E�g�d���6is�9i@��I�Ì]��#�_͠#��Џ�V�nݹ�kC��SR̜�,�1�\�՟��vJ�LuQ<ĉ�a�j�$"��%Rn����z��s	�e�:T%�����&�^7�l,-9���� j<��у��nA,��}¼�$���}�8}SGꄄ��/���F{��n���B2]��F�q��T�4�"�W���-�����4J�r3�|)[�������u/5��ϔG���	�Qj8�Q1^�ތ�B�t�~�-��1b ����Ɏ�k`~��gb����K�r(��< �`3�)5��c"p�0��1uS7:�/ͮ;X� {��S�=���χ�:uw�Μ������(�˻���wr���\4wT^=)I
����I.��p6I�oe�nL)� f��}���,��f�1nԾNUL�i(�b-��5kt'?�{R��[=���9%��Vl¼Q&3#o�Ve�ƾ%�[��/wcd+�-KJ�	���jo��Z�,&�⼺!3�l��2�����A�9��a�RS�z5*a�WFJ
}�Ǧ}_/��p��3Wzxh���w+6��#�-)�!���o�A�1���eW,��	�ėe��Z���q� z$�Wk|:9II����c�q��U? ɉ���i /�H��m��w�:�8��e_�ӝꝾO��ἡC�\m��>�#vp� c��U6��?�
NOY���zY�pŽ-޳��7&_�X�F�S?���i�٪�ꂾ\��j�!0[���!�U-	���S!���D�ʍ��r8蝌��Cv;z��]�DEEzK�"zc��:�O��s�!�
�ڱW��U#�|����`ڕm�C��MBE�Iѿ���ںEY�D�7C�0<�1�[QH�n~��5#�j���r��`1Q�Yzi|�x6�5�K->�E��6��T����q.�q�Rm��#���N�Wp�@��I��ʻ&3j�P��24�9�W�����7�'�LPkb�Ѽ�Ƚ��˷�-����U�I�gg�_�ꊃ/R!���O�KirG}��N��$��!6<�_i��� ���H�P��b��%�	_p���yD_f��Y���*0ߒ0A��lUε��%h� �����3d�j�y����y�g[K
����]�f���*Ԫ�*8:��4���{s�=�D\�{��B(X/���p׬^}AD�RK�<�B#���>�&��P5��e����.���Ӂ��]�?L���[�Zϑ�bj>4�^eDE�h+D���¸�"�]9Is��y���o�Y��I�W��Ձ���	+6�C&�	Ϳ$ҩ�Q)���M:��_�B䀽��9�kܹx��&�Y��Bx��hF�,5b��/	�G���ơr���FU�ן�Z0��;������zϻts}�u�+�U�ֶ����О���Q�D� ���(Z��拑�(Q�g3��M")��6w;���w��W'+z��+��.>�ҧ�2���Op��-V�cTF4�Eخ�b�(]'�,/ޑj� ��s�;��� p�:�AZ ��m2�X���JRT4Z���b�$Ѹ}���P�Sݕ� �?��U��U��3]�R�Q�K����2��R��7�N��LA@1l�SwC�X�\�?��5q��L��G2�������Pl����w#�LWC�з^��c�H�h�16��t,A���,�"6��o��X��O�dzZ���[Lߘh���*Cm�?�-���}�r�&h�\�$ZJ5����T�#�7�4���ӌ�J������Q��/�ʫ��������xf���,	�A���L��;U��C�.U_s�_X�_c����Ό����KՍkz�!�D~/����[9�<�M��*M���G���ث�9i� ƾ���%��X��F���*�O)M-��=Ghʡ�:?o��r�z�������V��ľ͖��80%��)�l�:�\`�xlmWƊ؉/�}4nYw�\ѿ,w��M�J�.�7�䑴W*J�W��*�]���j����Z7��c�>���"�B/�>���⎞�@�)o���;�8[�-M�\S��������'�=L��'��Y$G4�kc�Z�퀊�ѫ�Vu�\��ƸT���kл�ߝ�M�����PXJ�FJ�|l����dD������Y��kyT���^P��/��۹��_�Stؔ�K�%���J4mx�Q�l�cf;qd��F�lF�G�՚���A����IΒOEM��ľGі����a_��QA�4']z��26����ם� �ʡL�&� ��֪bKe�ltLs����T��@c|!������5�L��L����/�hyC�w���$�t](�\s�����)�hʩ2�٪T�O���n=Хu���w*�Qj���5���x9�AK0\�j�ߗ��-��9O�U���X�7(���]H���8H�jޠ�{R� �"��m���/\��إ�|�:U^�ۻ?�Y��b�+q>��~�K�p�/36��V�����8C�Td7�/I�y@@v��_�!�GU��[�L�>������<��$��Zx0I� ��x����
C�1����S��į̯��g1�v�f_fp���\<��9�2@�Sr��|p��j$�����}yP��k
ר�����4�����R��\��\D}SJO���KCxz��b*ڶg�Amo�U�?�}8!��#������D'����`|d)��`Ў_��И�ɧ(��ۂ��G*��'�g���T���w�qǽ��B�V��Ud���@�����֜6��:1[�#��g�/��f��ZH� ����%3I�ц�3�8��q��t�����tG���T57�K�0�]�y�āNth�9I�L�o��s�����7�_yO�7�щD~���pO�N��J���:r�~�ћNXɻg������wU�K®a��O�����0�<S��3��ECb|W��ו/ӝ�j��ྠ|Ͷk۬��F���� \�u�6G�:'�O��ĦK�u�}�U^�G,�Nٙ~���S �AUR.���i�}��4�������˞k�)3A�kr���}o`���ZK��t˖|����&�,�e3���{ۆ�Z;]j��Z��E���D��������-�^�fjK;5T�b�"��'��l G�]�}�P�z��ͫo���>��p�;�~5�1�y��G[��vc��|]_�NZ8|�=��Z�z0F�������7t< ����Z�`KґC7��=b�f �"'�����X�e�9��3�"��r���G?ЈD�c��l�M�ս�,��2�A'�G)v�y���r��{S���5�`mx�|��;/�r&Xo;ӱ:[<�dU�F��G�v벤2�wpQ|1-l����R�?�m����D[D�_y'7͹XYԏĵq�Ѣ����@m@i����E՞�Ñ�ӄ��*�H��W��S�e�������.2��0�%\\� gB��p �A/}r����ތ��)�������.Q�U���؏DM��;?M��騕�	Y��d#~��5Y�W�ۗ)��7��_�@mjv�������msz~��ގ��5| �b�9�����M���ר���xU%6�V$����&׼���/kK�M����p��_]
�U�_4򥇮�Os`�8�!�����U	�%���?1�b%�H��'$�b��V\%�a�az���ey�9Nc��Y{~�7�&^��v���rL�#Ţ1?%�����S�Af��Q$,_��
S���/ZjJ�`>.��� o@���,/������Q���8e7�!�J�A�2C�w%/ƢPbH� '���0�]�N(�i ?;t�a�m����:%��$	.�o���2G��9Q3@T�/���=���������4Fu�+��0{�Q��2��RZ�������/����ǰ�|�N̓���N�	=�t�%�&)��w�%	����&��hT���J�Tl�����J���P�A�H��:ہL��h�������+�!��r�J��>�@�a�[�o�����^��S{�.{z4-M!�x���UVL�oQ��O���-�����}_V5�~�cYy�,�K�SQ�|�ƍH�,z8�p��+%�
��S�L�2T�V��3i��c�SO2��S���$��_Dp��E�gVg�j����;�[�xB�=�c�/��J&����E��׈�DD �6|�O��9��K�3:5N�&N*��xލ��7.�����<S��w	8�$�e���#����X!S�-�@���3,=s�jp^%�݆]�u��]ؽaF;q*�YP�������F���9/A>�O���%"�I��7|��h-:����eƕ%ǩtŠ4�(��6��k�ul�Q�����ۋ��g����ɩ��M��k@�+��j�\����u���ay����l�^��	0<L��Q̦0C ��+��&~}�����z�mUu�kkL%�^��|�+'_��!�L��S0�͏�x>}�̶z��3��ㄨ� ��ƿ=�z#���](F�����Y}�bl=�#0P�Q�^�Q��+��ҕiik�Iv�j�z�r����m/$?3��Xj�(�����3���X���>n<���#q0d�D�b�j�ă�[���s�'�oS�M�ML�\��Ew���Y�����zj	 �\ѣrq�<����&�7������)��d&Yw&S��Myf��R���)�"��ZbtJ�[Iyx��	�`w8Y�VE!�!�_�.��� [�E�Ŭ(��=��*G��^�ح3�2ɂ[�w������.% �%��:���TY�t��w�ٽ�`���8���T?�6�59��i���^ �!�Y\ӗqe�n��2����{��.��>�j-;D���xL�-Vp_R|����J���]\�I��t��K8�N������U,��/���ϴ��l�b�2L�'�0���U�_��1S����Z�������^0�oz�:�A��Ws��m�̔�<,d�<����Ulb�g�ʴ�lN"���Y�ZM�Z���)ҦDh��c�t�4]��v�0�W?�5���)����ydg;�{����@*��
�M������ig#�z�_�4�@:_���Yy�]��N@6&�X�����6v����㾉c�3U�5��+�wB���,EE���Z���n�gf.�yZ��*=��U��K0����Y;/y@��,���4=�F�"xKA�N����7���D��糥+��Z�LjG����ᔥ���>��(pp����6����	y�=ž�K�W�O���a��[ϓ��ͽ��
�~�D���BG��Gr��6S�(���[ר�X�S�f)����zs~�F+ʚ �``�������i��k>n�ct��\t�^x4TOh�Uٴt:f��6f��Q�i$��w�:�c!�
U%g��w�>�N�1��M�Na�1ydꚬ�w��&��xth�ڋ��b�	�+��B{>X�&?��Κ��<�cCX�I�^Ivk8�Я��oK11�h��-�?p+蒐eɑ!]��F0�C��o$uH2:n31��h�m�ph�hE�I�x�j��l&w�g�!��Vǵ��[�m7�����u@�B�[>�g�����������#K� �@C�|���]�3wD��w��I{�bA�#�k.'���
�7g؋���TG!N%�����HMƄ��M	CA��]�t�
��hBή�f��n���S�a����҂RlG�=Dqm��V��B�dZPs�.���:��A8/B��$P����|Ƞ�M����}�KI*u��Bk�QY��������L�/r���Kaj�:� a'�P���y�j��a�*�B`���%�&��czU�Jl}�G��1*o�ox�m;!1|��>kB�r1�DN�&\`�W�C;�4�/'Ѧ_#�;Gוmp@�߃+P'��,����Iz��z�$�inhBz������ڟg�x4�6*@=���-?0w��|uo`�z�ʴ���p��ͮo^O�ԝ���Y��*[F�hP~v����gCf~ƺ��F�	Ԑzvc���4@���X�Ou���Lm��X�M��hu��,��Q���5݌��ʈ�����s�ElK(k���g�y��2�V~Dy
���< 䰨����ql�na5V�A?�:�J_�����>�7��g��ΠU��ݞ��d�^���Q|�0磜�;��&*{�&�Wo�D���:�����
m56+B���P:������O��-R7>�K�y`����F+[?�j�����y��H��|^Jb��k�8��3|��^��&`n���,��8�cP_�JF:�Z�O??�C$�Ӎ����`�3Y_§�G�(U}c*�7qr�$�F�AA`�
*~cVOyKM�Й��#� �9�N�"P��~7P�R?�2
�o���2� ,8�)��f�;s������^ �=������Ᏺ%��E(9�(�_hh�&�3�/T�~��%K�E�,o��Q���b��P�=�ʌY�M^�Ɍ0j�/�,Z�m�,JA1����e�ð��(`��� Ϛ'�aL�;^9�6�R�\�P�쫸Xnc�Z!�|�i�h���\K�ƿ!���룕f۶����l���7�8���OS����CRʮ�I�%i������='��9+���V]ᙦ�w�[���u�u�"��C>�XR9��ںDu
��$���qZ�
ʠS�Ly�U̹�iV"�z�N�䌍�Y�*jCk�v��J�W�EB�-Ҋf�<������G�^�W��wZ�ۙ�O�tZ���w��1L/��Kf�u0��u�1��Q� 	�0��3��8�۫`3�|OAAL�P	)22���@.��T������}�/@���M�F��F@K0�y�T�;��lN/�Cry�]���7�bi��Ov8��}�e:_1và0ۜP,�e��\�ቜ��C�Z��nB���K
���r�e�iE��V��d`��:=$�|�T(͕}��!uQ�h��w�`2�k�ê��Al��KO���DA2&��KG�����e�@�R+u
)����"GJl�}C	�;(Ґ�X�Ź�-]�r�n�*��Ōɺ��#� �՜���7@Rp2 ��IN����	a�a�������،�SgGDX��鿅Sf����ȇ��:�e14)�x�T�XĬ;,e>P9R��"��0��.��I[={w�
�{��eO]9ͦ�c�o���O��Ewn3rv!�j��8H�y�9���ԙ��f�8I�NJ�y�ۗ�L�pn9*�a��Zo�B͹+�ZU��}6VgL���/�}.r���>��*�޿�����ٰ@�n�|�p�L,4�=jQ@�ڲ�P��5!��X<?�I�/X�(�Y��A==��1���7�]�V1q[��	��
���yZ�
 �'��P6�!�������F�����mr��xV)@��䬲������c	ڹn]w�v�L)��keH�=\�k��(j��_@ �"�&�Ef���[D^b���&~tl����)h��Bx �j��쐢~统o�S+�,O������`J�޾ ���\��b؈_h�~ʣC��a悔��5��=�]3��fI�Ha���c�1ↄ�>�Y�_y�s�_NA��^��@�a����_�2�t��:��<��5�1k���)5�n�X~�|��7��5FQ|pՀ�;�Ś�f�)-��6�\7�^��}Ȓ��X���H\y�����؁�^s�Z���@�oǇ%��>�P����$�z�7z4{�p���5l9W~>^GՌ�M>�22ET��٠sJ/x�9�R�jL��9Q����H0��΢�h����9"n�^�x�C/��<W^A+���e�ȇ�sg9(����r�{�Z3�!�l��Bh1o[�{m����΄��y�1��J��톥?�����3q�dP�nH纟I+�-�����H�����Ś���� zT@��m�� �FF45���+������8��i��c��}#����M/��Hw�����P��v�`0�=��|My���wmu����X>�F�����S"��_���h����*�����C��*�\s97$�)E%��1����:����j	���Vޡ�&jf�G9�����lB�?G S��i��V^�����*؍��D\rb�p>7����x"/���=�T���#���H�C��3��o�� O��F��8��R�����%�K�
�@���!��L��en1,>�my͆�`�z�&���v@(���AJ%���R�+]�EE�>2�Sq��n�]�$<S�k)t3��M"�PS�m.�i������>��$��������F��ཞXg��ܸ�R�l�I #2|��hN��b�c�XodHE)s���	�z7iDj3��pd�Bq��,�����=VK�&�x3	�o��y6���?���ԇt9{�[~({�6��exy�4k���kz*��� �����ʂ�A/@�w�	x��3�ː�6`���N�fd�寧h0f,1/����3|оS��,P���˚��g�A��ߕd�#�&"�1��¶�Pq(u/����c���C�?�8��D�	����R·� (U;�и!��6 )L�Ƀ/yG�]�K�D�WLڔ.r)������`���ŦFc� �\����k�޹u�w�t���ލqx�&����3�
Q�-S�rN���[��Ҧ�	��{��`6�ǺR��M^��
��,|U}����m��s�,7�p|��QW���M{�D+x�IV(�Qu��Ę���y�$�<~P (	�hԹnOQ�f��4�4�s1Xn��wS/y��i+�C/��d� ?�~%羥KzɎ0�U����T�8�i�Jprs0M�{�+��s��`�qE��7�D��<z�,3�.���&ɍ�;F=���$q]�lEU�k-�Ep0B�y�>�%��X���|͹���ws㎾uY�#V����V�3ʒRh`�s$Ȅ�>cT�����A�r��iv�,rH��S`<]T���\PlvCkN����Y �R�t���O�5ݰ�^�Oƌ�Z�8�8 `�!����)����H�b�2��6�̯�P]mp��F��1ERD]X�	n��6�g��P������nb�睤9�r/E�2�8iSH����T�)�GHw�Μ�&��nx�e�F�j$Yo.�񝵻=O�B�-�r�F;�i�Ov�1��z��0���l�=FdRZ �	C�T��v ���]�N��rOЉ���QW����u���� e#1�U�7�R�.ݱ��ЁDDv�Ю�H��X��k��6��3�o�꤇�-�߻1!d�ܥj��/��*z�J%WgBEa�Zؔ[oY׾�PZ�U���Ezu F�8��� y	��aJOK�`�������r�!�fw__.΁$do�R9�䁀�KSӃ�Q��s}di3+rހt�i�.�酦�v���`���,�6�i�Mm37��I[�N/d{u�$v��'��a��uK�_��0�����\�ᇅ���ܘ1Q��$^j��/�KN�23:s[��	��9�Y�b-��Y�݇�$٢\g><U�&b}�����������쩳@����;_4��ҍ$���^�3�\c,����_1&�#���Jv�a����cd�3H����m�mOx�Р �%���\�6"b�y�G��a���~�{n��Y��7�	�#kt�f��
��m�ߒ�x��"�W�>�x٧g�507�,�G%��]�R�����]"0��sb
�wOϸ�, �~���r�~�N�hq��#����Q>1���G|!���f\���L{��"��v�q3c�5���3 �s�p+"-/R1�~u_��������_-?h��8`U�[+���̦5
�����+|�P	C��!@̐�=���R�����N�>m]���aS��>R|����蜛%5�lҰ%5�-�Ho==��D��I�ӏ��2��+DQ��^Y*����Ym��1�o�F��>oo���Ƌe��R�z)h� 1��))N'��������o�����.��`�h��{t�E��`��
z�1{pA.*�?�df���9�#�r$�	"I��m�E�𜞑�ru��@�+�cB�Ed��~}4��g
�غ?r:�Pe~�ᩤ6.`d�Tj��=��(�9�_=�w֤�k͊�v��JkG=⡛�s��CT><<*�^b��đ�Z)�k�b�D^w"��X�	�Ň0`��V[6��I5�w�zD�~����Il�=� ݧY�*A��Y�qKU`����'=��U�j��|��h`��4�ŜX�l������	�z7��g �c�q��SEB�Eʬ�t*hU(��r^�j����`�ZU*�'f�#���,"85ה,]eBq*D(!��`�Y�؈20� ]{�נ�4W�b	!Ti%��t�n�X}U>F$s�IK�c"�����ҍ�VUb׿;�y�;�sN�� PA6�Kr��44ǰ�U������r���J�u/{ɊM��ң4.W��7�����:��*�n�~ n�8�
0�ntM�]��T(<G�A47�/dIh|wC:ށjv�y�H�q�'�~-�:ɏsOԓ��X�q2*
�@����!��%è|�zl#.K��zh�{�W����5 V���g�A���@����ȭ+P-��~�1�Dd 0��n!��B#�-�V�ϔI(DRd�.<�1z��&�{�@c�zۇ��b%�/5F�e�2q��0�'��-`�Х�UN%+��I���}!� ���w��c��O��Х�٪��{��t�-H�z�I��c����pD�D�&�-��[�U��hmJ���w<S�+}�1��-MH���� �E9�c����E�&�Pʇm����\�_�q��ڗ��N�� |=N8ؿ�b�[2;<u�ǧ0�)l��Vٷ:����ϦN�@���G�/(�@��9�u�C��OS\*Q�!�R�l4T���<(�Z��eÿ��]�;H�{⬑�VW)���N��񣡏d_OT�Ei��Y/�[b��o��1Zր���$��̟p�(��ke)��Q�K�(:�E�[�:Y}�e�^� _A��h���w�5�bV8�M����\�ބ����!��U�7�2�� ��b!�./���'F�4m��A�B�6���ɨ���D	� _�t�(�ScX06�쏌�[���?��>�����B�$Q�1����uX[�@v�)it�9�jqϟX>%̨�[4��� �ʗ�����4�0����Q_�c�
��X�l8��ZM]�8��*v��S��yT1/m�XP������6|Еzk�Nvm�����Ŀg����@B�����}Z_)�+G�'KH+K�{a�b���U�ޢti�����9����۝fǌ��a�s(;�_ۑ��W��ҿ�}��L�vS�x�Gd��I���R(쯦Ā@3�����r��C�X�3G~JR�(4DC8~{K�%���͆�M ���	Yo�*-S�Y��)=�swLᜠ�	G4,��Jl@�)�j�B��	���,��N-c{$�G�G[�K	�.��&G����h��bp�8�烍�c�"��BDO��ZǊ�H����w8J,�ȟO�[�� @���wD�V���F�S��|�}*�@���ѧ�]���T����"���[�i<�de���s�\�����e��s��+s6�!����g���c�ġF�<�6����a����mxT~��si҅7)ش��X��)�՘)�E�4c�d��P�Q�R�D�����F饮�/J�wX��g����`���\��9a�/h���ڼ��n��ۙ����J�bp��ӣK_z.3���.��Յt����s�����ؑ>�w�!�׸i=�\3�k����Nu[���q���k���p������o�����lK�U�4%kF���U�Ku脚��]��1���:~�<����d�]?���ה�gGi_�5U�sg�u�q���"��M��GNI���Ai	Ȃ���[6�����N����5�{b��l0���,T�i� �M1�3P�R)�W��ҥ��_��~���)�����=d����5&�<x9���<��4�{ܘ=]�K�����sze.���M.s�!�Ys�d/7�f��'�"�k�Wf��Љ����w�q[@z�-��5 �-ԼN���{3#|�-ִ�k�{�7Q����К	����5Ύ�:8U_c�K�h�[a��AT����w��o�iVl/�)R���=��.k'y�����y'x���oy�fUrX����%����EE��b/&"�IY��km.��x��L��J���1*٪��-Rs�ǃ6�p��a�x��'��2���5�}�3�`3��m��p{�����`xv�3� υ�B�E�.����,KǴw@.`�����RO��J�C�FI�@HF,y�ڍ��t�^�o�ZH�iH}pݽ��{m�i�o}��MbiٰOM�?"�����qI��bX��}�$;QCQ��}�x��U�fi���nX����-�&s|���7�6�s�3�|�?YLpWСJg��uq��`]��PB65@��u<* ��})�E���[e�#䟲��SpG��7��W�z'4H���_�Դ�*�
�r��5��#2�L�hdCl��+r�l����>�,��R��jI�Sn��M��I8��_\5�
��?��C>+ߪ���Y�,};'7�� �W����T��n-N�t�bO�l��8�Q��KD�A?�bLzu|�i�A��1�d}�DVfg�Tw�t���x��Ld߲�w
��u�ߵuou��80���.�81>2���`cbx�g�2�_м��y�fg�QA��$&(�GG;78*X�P����|!�O���4��<��=��u܇L��u;�����6�	Y΅��{ş�!��F��	��E���p�0-�y߶���ԪCQ��7�\}�__4�iH��#��Z;q�#����>���xb�{�����=�W���J���"��� �,l�B�U,8;=� 5���6��d��E�����;I:}HN��źF����`��q�+��&Bo�%�h~�#�i�^����l�&�VدJz���MH���ҜH�W &����Vt~�Mw/�.G_��g�P�eT�izbd6����͊���X�8��U�V�5<�]6¦��\eO�1��ߥ�L1Q��������)A����$�j�<�S���,c�b��Aq�|�,�[�7"W$Jȧ�r>���s��M�4�ʜ?���ʟFD�����8<��.����׬Г�� ��(��ޔ���M6J&�y��	iY�%������	�W8DL^��	S.w�0@'K��ي}>��!$&rc�Q����&P���E-�[�r�H�?o�����bK�(��zc�͜տ�0]�ۤLI���y&���7L&�x��=O�a6��>�	/cO#�+��H*��>�Zi]� �F�Ψ&�V�5\���d�����枟#.v�F}�Pk�"`�Uֲhصm������O���~��X/Z+~����Z1GԸl���p��wyJv��_��-�K&�(RG�P�@
h�U~<��__�cՑPG�Pd��U���9�����-81u����$`n���Dit߶�0�?Kw�����}�x����9�7&��y�K���3�����_%� Ol�z���7��Z��.�Ⰵb��"DW��f{1t8��
�$�����*,�`�f�;�+�7���O�?��,��Õ� �������si��rlFh)�����,<I;�?�j������m�y
������>�p����h��6/E��0�=�����z�{x�0tq[��@P��j^��Ot0��M�ms%�}ݴ#m("����;��aL�'�18xp����f4��t���e��U�9���t��lyl�%D2�ПNW��?F�}?}$��ico�:����
��Wbim���!�+�M!��T��ξ��382�t��r�*�2�6���c�q�_��o��w��^Tz�ٜ����O�,�g�弔���	�:��B�8 \��<�6��=^=
v!֚�H�nPm���BR#A!���9;am}@�GR3���k|I����e���"�JJ���-��4/�V��*�ؚV�񰝤�ЃRSٛ�T%�W��*�*@\�v��ȍ�[��0�̖܇5�0�p*�I�MV��x�@k����+�R��+'�s�_� U�M�V���A�U�S���1G�c�M�%��I�<��%.ߎΞ�d�����J�]��S?�Lgs�{��i��Cd(��<��Q��}J�����#���\�ߥj��h	,\�Z;��8�Ap�0��m���zU��:�4�vy�Z߶��	��52�_1d!c�P>���L�����ec���GT(�/���wGe�?��"���JRh9�O���{=:ߐ�B�%����!5E�sː1ث�4�⹄R��I%�
d��>�YG�˻�D/�v��M����$�0jD� ��R�r�d�8r[H�/r�O�毀�%���z��k,���<�t�� �ñ���e6_�0���0	+�pL��"?��$7�eF����!e��&^賩d����>ڸ��Y�����#��z���\W1��\���]'n,�1���"���������� �ės�T~��~��/qR�TQ@���i�)��h���S����\۲�� 𚓋������/l��i�C��R�6zo�ï�1Z6L��N�_{NQC�=��4�
��B��m^]�$�~'�+3�u�]�>�\���HѠ����@�Bn,{��`�5�Fg8XGu���<�2ó��cأ����m7�3J4�zʦ5 r3<�RlV"�Gp������:�?:*h�*	�{
͋t����`��ت,;�.���"���\焚���M�l�O����;;����P>�`ƖςT�C+�כ>q�z�,C��@ϙ�Dv���>
;A��~���R��~!_�A-�EO�E���ҐY��hRHv�/�T�GX'r��^s���|�Y˶f�6�jBN�8��ޡ�#����A�l�sl�����O��͚=r�~�}��6�W��&��ئEC�"�LO�g�&��-�a�{��Au���ciZ+fq�7Ļ�a�ԦkSH==��u��,δ켗ŎP;�^R�����ٳcNo)�m�h��jY<�#��xʪ��ʅ��9|��S|@�.�4Y����WF=j���+.ť>��y�(�<'���d�8���\���oy}��X�72�,�;�̕���0l�PYe��!�!Q���@�V�7J�W�#��x>��!q�ci��?�U�A��XS�s�^>�%����&B	�s��2�����$�@����n���Z����k��Hr�ޱ"�oI�l�*8%�b�|�z��,,+7W���n^��覡�>W2�C�p�g��'N�hE�rGO%�VҹY�^/�1�肝�qj�N.�3-}�,:5\w:`T=�iv��Zz1D�?�y&�l�m�G��9�ū�q�}>��k����hG�%�0�D}�XU��~���1ٶ� x���FA�~�G���`���Ĉү�:a2�m�v�^�{�]7�zkc���JO�H�g���/H�W��:!4��$fz)�H�Y�|���璴��C�Ѭ7��AN-W��¿ji��RŖZ�(A�U�٪ܧI�PQB�=���U��>�A�+��
5��q���2�+����g6q�ky�&��px��J���B��IO)��GG�'lM���+Cs�����;,Kh1���K�߂a��2�Y��	fv�Z�/��03�����oH+�O��D�9$O4�6�L�����˷��H@�YHʰ��e`��:��?l�Aّ��]sݙ�K�x>�?`<!g�]ڀ�c�.�qq� ��L%:a�9�c+�6�-��"E%��/˭�.����iu�q��ʋí����guG2ɱ+U]K2l�1���O���8������4e�2@����԰�f��5?�<��G�i��=�&��Z��~�q�,������J՛��[���d�?�/ ��4pEXqi��8�'����� �lm<�H�^7m��'���r	f�zjѼZ@��`@w��o�{9��I6A�`=d�<��n�����cq�� �9��|����f��S�����h&�au�J�_���f��
[E��7�$��b-�i+���ϻ� ��d���#��r�N55���t��*�RȘ	a��\����kNP!�ݸs㷸�-/`�n��5@,�= ��ʶ_�m�I��=s�ZhiPwn����	�	H��2/�~����\i ?~���A��BJ�@�"�^�d���q/ ������P�F�F&KЏ�V�v�
<��x�}�9^K�*�K��f��g ok5��)ĒZ�e��<T�������qx�\��Kqv�E��m6�$j�9����O�o����WH� J"�鶍���͝^�桡�dP�+�)�Lh�3&�>�Zć}��υ@�ƿа�Ob(5�^󶵮G���A?	JxH
�!eE�i�D@�u�vA^��Z�ݮL9ڬ=���Y� ;&ڶg�����RϤ�X�!Br�����d��>
r	��0�.q��jB��?xl���(8���+\@diz?�+;e;>= Ba[AU��t+Ծolk�h����Wp3Ož�S�7Bвa�yg���}z����
d/�P��]`{��Z� K���g������I�Y}?G�5#���lA	��ͭ�ӭ�o-C�s�%xd�@��vl�N
֢�QW���l�6�bJ6�;<�=���PFk�/��qX>��uN�Ƒ�C�b�>�� �|��*F~��u#���zߵ!�kZ���^�` ����D�?�
"�r���3��?�A�hSCYrw��[)jjN���s��^������#_1�B�Cj��h[�B�H0
'�j|����+�Uwλ��@�߃�3�	��!yz �ִ�5S9"�^�[�K�N�^̱O�V���{Т�/N��-&���sf4�Π�{�9wū��A̻O������yF!]���Y85��ҿ*����ᐅ�ߦ/ �-9� ���SWpG���A��jM{E�f�
�����V[
|������_�FI/��q!d�J��c��k���	��+ÃY��Q=g=����ٙ���z�G��!^�2
��F|n��{q3^6��m����{�V�D��	3��%#bF����f�a���j�SN �)V�D�8������Z���H?��p�_�Bu(C����X8��*u��h���)���{Mچ@�J�#����1Ws�9�{5�/�dM�W����t�>�z�(���k�#�f�
�F��*��e����1���0W>}OzD�U��=D��fWo���t��TQ-q6�I��J���5�7��F_����Z�m.8x�i�M2��E/6��3���L��  =�@�mcDA��%�TA�tK��=��"H?�g�������V1@;r�@*���b]1�����j��;|�˱s��z�#-�P�r��̂�G����l�Pl�G�e�Ue�^B4IU�����K�tz��w��)�>����Z�B?�{G\�(/�Kzd�w���+�b��y��E�z�#��+�*`e����`���^k�]��p���5���{��-�Dh�e9b�(�LfP	; �8OO��A�MPM���C�Ő��C�l��"��3S�ۻ�,��& �����>v�,��.�F�F�.���b����j%�Q�眆���Kk�����i������uÇn�qx�����9t�����J��z��?폦���u�V[�i_U�űu9
P�u�G$Z��c��\�����DT�a����L(*r
of������Em���m�/I��Y�a��d��s����3�/z)�?�G�t����Ut6\`��Q�+Ϗ�>��fn���P#м�ZƋS $v��`��7�{�lǢi��~,<D#(n]1Q�Bc��v���i�V ���L�AE"ѥ&29��K�ob���%^����y�^�ܹS�p�b��b����\�N�vɗf<��s	���wT��lz*%�d���#�&�1���C����)8	�}�}$jrg�y	�?��m�O�T�[L��R��0R�j��a2�>S������qZ�qN��\����tzŬ�7��h�� ����Ը��q�(E��[��ڿ����?2j H>�BC{�v��x���^��N�n��M�Y���������V`��?�I�=Y�.��i��*������� 3E��d;*�[��ej�j��M�7��
@��AU��X��:TXs�|�6w�~?z����D-��q����Y�&{��2!��#"�eiO���4. �Ѿ
sP+���=�E�8��bj��y3�ߟb�5�1�e[.�����94�nڄY��E���ơA>_oT'n qb��SI"(B<�vF:�X	>5�V�Xʆ�A���Ɠ������sԟ���sM�M�vP�6Iߟ�ݥQ2�X����K�ڡB�e�Z�)p�SYz&�{F��v��vkM"�±�Hdt�o|]���6�Ɯ����`xw��~�sN���G����G�r���r�3� ��v�j�&	B��lF�7���Q<D�6� �r�ӣ�xpo�sjC�c�)�]D���M�����[$�b3��S��V)x��}�Hn>!)v�;[s���I����Oi�fE��dk騏�{z��%Yo�ʁ��T��^5�Ɨ���!l��*�`�hT<����ο���r�/�M�m��'�k�`�F���.$�xT�V����3�4��*=��_��7�8����d@y������\��b�Wgk����|�~���.�?w-�	�^��UkS�:�E'��VĹ�\�csŪ�6t7�4���(Gdu�����+.#p�#���7ּ�y%�A���)=pS���vi|���@ jaC�}��e�3}*��K&�&U�!'��kիf*q��Y}��gӲ�DV�C�eCNZ�(7�vnh�ê#�9��JYo09
_r���|�ߝ��uSCOJ7T��sTD^���,?Y�hÃ]բ�RhXcF��~����.��{Et�QZ�ci��N�z��U`�.�ۢWdO�ꎋ�t&k���c鸪�����/~�^�h��4á�����k��`Րm8k��^ަ_�-m���)L����H�L�ؒ}��!�ZH�8X�"I ��%��]�X�uJ`�{��P��)f����_�f9����˘^:&��Ğ�p����R�fP')�GN׏�@DO
R���^3�Ž�Ozvx�N6�ϯK^��]|D�!V2�_�bJ͙����M��b����3���$�:E%q>��e���=\jA�2�����R%�s�=�d�'��K*X�o��b{9>�3������2=C�!C �����_����
�I[�h��&��MA�L����j���X��HDׅ�ܴ�|E����V<M{��ROF�R\$r�'@����`��n�(��O�S���O@��Z��|Y�E�ء��[���^_[����	�8�+��rM*"�}�X�g������l&������K^k� ��{ې��t]����^�j�����AP*h�Ň�d�C��Y\,��6$�g2S��Z,5���̱�Z��4{%������ژ
2M4��ӌR���Gk�	rj��l���(�j�� �h��L_6�N~q��o�o#M16&hyZ�N`s�A���^bޭ�\��w.��*5F2K���֗b��[h�G! }�n��$�fԬm�5��LF�:I���j`���a/LU4��,��{���������uE�����]�O ��L���o�ގc��4P(6uQ:�k��L�'�lh�|��������JrvkC*!�z��Ǆ��7I�����rp��Jj��`��I"��6(>�����E��L�Z��!ν�B�'i6���:��V�!�""W[%c!�X���Xx~^�� +��}���	�Rx��`\g-kD�-�?�1�����&�6D�ewcw<X�	���1���ݫ�	XB�w�o�T�/KQ4Fӂ���ͺ���ߔQP�L�vlQ^sIRE����x-i�/E���ʷbd"��c�TF(e�LWGmҴ�,���N�M�fp9��H V�r��[�'�R�z�DEB�TV��us�c=��I|�n��upz�Xw/��~�Gy�SQ����I��K�Y���Y�5���	P-i���S����w,1� N7�8]Z��WÒ]Hy%Ur����^�)[������,f�7�VG��4�����9pa�fbm�Y9o�fz�dEm�]���zpJ�K0�'�������!�M����
��FbP�]�m?��u�I�{F{3����&����e�#��=�GnM�MG���Qę�O�n [L�t�q0"��p��&�{
W(��b�^���Z��j�?;f
!�c��T!SO�a<�t�����Er+������A%V� 	�]�?w&d$�s��$�?��m[I-�8��Fz}��l��&c��Iʰɲ+�2ʁ0�����z3ٚ�F�����i��?��-�|�����/�y�FT�a��}'{-��1v@S� JC��?9M���=�������5'� 6j��ai��V�9��∝�̭e���Ӕ�τxzc�>Dԛh����s�3�*?�>k�d�>u��_n�� *�*�p&�MF���[i����'��#��j4>�)��7O�p�e+�`'b:L�=K���X4�a��	��G��q�ǀ�#\�Ϋ�Zsљ?�SN�z��{����%�c�Jc�< ��s��Kv��)�z�{q�Lb��o?�v�%�߯˴fc�>�Z�6�gk��n7�2�p�B!�dR��~\� �U��G�g��f��sC2H�6r��,���.�3�c��3x
F��񛔠 V�!�G��1q�k`I��0�p�þ���\�`L����`?���j��V^��g��|���I���_� !���*����x6W���O���r(�Ə	y��J�K��'�����}��j]B �z�Q�>�2$�������r!P�}��M�/4&ۄ�>�2���B�h��xɺݴ��F�N�V$���O�$�-�A
v�w��9�W���Fp �������1�"e�b�L����B5S��R}ы5�![q��?u��×_,{c!I5��e��JDy��?gP��������^Ϛ����Z��@�q���K�X��VU��6��6��qL��'�浉�3IEq@��(>�HT@����s�����om�_Rs �a��j����kN%{��CB)0��t���P�-Zn���?_`3I��bz��g�b����k����<��l`8�Q��w������Ș���Y���Y07N�{*tҗq%�s�IT
�Y���y�dT\�LJ]��Pg�t?����
�NTf��*����떂z:��1�%�?�z����#Ϭ���R��<Û�)!���4��L��Mc�t����

�CPj���z���?CUm0��`�e
�N���:P�~T��$@�Q�=3m[�:�핸|�`�O P�x���ص���HUM;ZY0Q���z�G*b�܁俻?.4}��ￚN�o��3=��qh<��t,c8s�{.��$�hN\߫v:���>3��aǑ�f�� ����@���Ţ��0i���&��+4��+^wY�fc��عm�D�������x�Yޡ��&:b�ר�\7�e��(PV�1�r���Zٷ�aNy������\o4�p*6�9˼Q�h����f�����\<J��T5)�4�w�W7�3P�%�lA߁꒓?_;��6��˴�Ë�'h7*�m^�$�_u��Mj���6�m怀��RF>���v�ԜU�����C-�sP�M&����K~���n��9�s�w�FJgh���G7+�?~��z�����K��=dԓ�DI���#����d"�JAs'&6ݒz"�= $��]eS�9 	��-�������.���80`O��wm���5�C����]|E@�3���&a*��j�NF@�R��B��:9&�_:�1A�����HUUeѓ��"�9%Z�Ģ�)%{1��d�;�7n�`�i_S��q���Ũ���������t��xz��$��?ҹ�U�#+w{YT�����N[�G��!V��J�oI'r�G���V��h�3�u��������֠�{�l�)�/�	�d��<Cj3�U	���"�N�1���>���̓�(WM�����*��զ3l !0�N�3r&͍��E4$���=�� �\c�u0��"�}(S��3Y�ݿ����yG9�n�}�}FXj�*x�Δ(M&N'wZ3^}1J,�+���%`8a�m�O\�s�¸�[��(��Hѳ@�7i���?m�gl���n|O�v�V���S�q������Oܹ㨡�������Ze<�Cl-�
O*1��'��INSr}M	���Sz�P����?�r�ٍV�9��qNj!!d |0@q�����h2��U��7�1���k��\U���i\ףw�N��Q.<�م���/<���^[�[t���gR�J�7��#���>Y�#�G������:ϰ4��G-�a��e4�}��4���
g ���;k�t^9��-���ks2��@+l�`�y�Q���,5���]�>Â�4yJ��ݎ��(,���( v.�Rң�g�u��+X����_�+O�RK�[V�4>�K`aU�k4@���a9H#X�#{-�M�W{rN8�����a^`'CO��
@6���fO�N�q q�4���=a��V=�E���םL4���f�IJ1�zДy6P�<��c.r|6P&��]p�Z���/e=�bd��t�D�q�ʷ�:,F�	�,}�D7��!3��x�D�g{.�]��3&D�����Nˋf���^����'��H��X�Rh,)��+V *���*µ��k�<���OĔ�-����V��'��B��	�L�ۛ���Y�P�-Bɍ@�'�s���IɪDֱ�1��8���!���5�a����� m��]����U5����!�W�m����T0'E�N
�	+=87g��ۺ���V)6����1X��5�ȱ-�R�)o�w��t�Ęx����K�����|ƖQYpY��L�J)�)�����Y"�S�4��� ��-p�[�L��\�x����crt�X����y^1ױ��k���Ε�s�(��Tyq#��xؐ���5�W�̍nX��:�8�S1v�Z��C�p������
g0T����
M7.0T��& D�cez��X��r
5�!=因s��˂Í����m(غ����]���A��1���b�^��\�=��;�B/��`���g9�p �$��F�u���d�V�4����jd�EW���WǿmF
ɮ��%��#Uf�!��ǣ��"+3�V�8�	�qQ��D�FQ΃�ɻY�V6��Ǻ����/>,��}[��;
"��-�\Lҧbk�W�E�Ư��8fk+�-��U�l���������[�k#<��W=���[hۥA	����e�6<.o��I�k��~�6)�b��-����kS�B���� ;�3i�(e9��#oJ$�X�7P���'� (F���$.��S2w�[� �\25k�.ag��t����p�z�ޯ��W1�\$s�s��V�����R�7o��ˮ��2#�|f�OY�tx���N!�(�^[=K)��;d��_T��n9��A*רnM�A_eCxI{-r���,C���kp$��E��G��f�t�F�E]-$�Pk	[�i���[ w�����m�_,�Aٞw8̑T��=}��������"yV���4Q�|%�jC�j�g�v�mӞ�r�h��G�؜文HgbF�.X@t[]<��0�*H�$Y�H/�6��%��?P��YE����8Jr�,��%�>$��.��씴{OԿ�@:�6�0����ģ{3��!2�������� ��h�*�|9��
����p���I�'!i�������Rl1BrLCJ��Q��up^^�a���(0[X���������j4a~��Vgo��lt�:����K<�_�gL�X�)#V�	i�2��B�J��*����`�q[H�=�x`��S�2����=��jEլ�fL���;�H��]7���"�TyZ[̯�ҝ��'OݻOY��S��%'�oO���G(z!�u��U#j;�ta�x�)'��Q�?��~���C S~�u��q�� ��aL}�\9�+mMqE��7�R��ع�S�[�)�h��3�K��� {�hq�S��aܘ��@�������sZtC��i�WD
~������@����ZS]��������b��G?�:VS�:�*�E�Ȯ��@�'$i����[���R�-�3!����)i�	���t{�:m#��d2h�E�o�HHw�?T�M�lC�xva������g��wjMK ��}5��F7��Tq)j�xY�2�� �$�D&�bl�#�ug/Cғ��2�TU0ϔ�N�"���1�cb4T����'�p�K��S-e)�d)>����S��q:�5F���C�iUI�0�b�8�*�:\4��mqَ��r���u�\g�u3�&̆�E��\�����Fw�;D�@�|��k
}7L 
[5���R-Lp>L�}Q�ǴhIy!���5��Hm�vMٱH
���G�� ��`���`�@�#C d�t�|N�VCb�a��l��蠇@ z�}�*�}�R:@rp��/���0�mM���������0��V�yp�����5���1�9��N�cI�S�noO��kP��qE�W�X��%�kQ��a�G~%�p�`� R?�'b��z6��,�4=G�w-���V�%�s�=���iK8�U��83�����$p���&5L����JzӨ�"4v�Jo��(��M'� ��[��������	�Q��T:ls�l�uD���~pS��Fc� ���~y�T�9Ծ�}R��#�i�G��(N/�@���r�7�_�xH��{�Zb��
��6,�%I�U�w��.`�L:���R�YEՒ �C!�.��X�㇠Vo�*��.d� �Q�ㅪ�)GU���⋊��7��6�y�!��i����5�dB{�~��y ?��tBs�fQ��6LRne*�E��� �l�}t�t� v?���纴f�n���:*�r�0�57Q��n�xVfI�{T�ʪ����-+NW��[D)�a{Gn//���[O�&%YV�	Xޓ#�d�P�Boy�g��u�Lק�ﵠ�]G��%b��! ?�ڶ�m�����M���OA����[go���#����shc�=r�`C��f��/��#ņ���n��p7ڐ�
��1��]�^Yf(JD"�v{�ӟi	x(����	�W'�ijd�(����B5+�	�D:��RpCs_�+�I'��a$�5z������۠�k�kG��[�h`�p~=�z������?��l�VKFE���p9��U�af�:`+��tq6��Ö�{��|H�/dO(Y�D�M\~��B�m�(�j�G\�*�����(���ېJ}(zǇ������'i>^s�0�!��w����h��a���$�А