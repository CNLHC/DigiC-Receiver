��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ������
f0�L�J
�90Zy �?2����4{��8��;ӎ�)Z�7t�Ot��L�˽��#�{x^� �O	�,ѯ�-!r[7�F�ǝ�EL\x���!3��L��È�a�j�� fi�ƹ����{Š�'�x�E:�����z�;�d{�I�-�j7G<�P"icFl>�0�������5�ąK��䐈���/m'G|��!o��G����7��H��`�z`�N[σ����mg��F��X�t�������܃
��\NP�2}�4�r$H-�X���QA��s��ϧ3�v�}���ťa���(3A����?]P;k�_f����I��	�m v�5�uɓ��MY�z;�]�V/9��-ll'%h�_�|��kr�Qʦ���-Ft�2]kk���u���mViE�j����}eO��>�S�&Йĭc/"�aҹ|#�lD�#�)�6���{04��!.�����r�M� �d��#�K,y�jbDѭ�Ԯ^�2��z�s��` �u�P\��o|�XX����v�_��KNf.QsB$���ǭ"�}fu�ysme����/�6�n919a� ӝ{.~�fO㛇LM�����.q%w���j�fCg��.2;h�0���h�#�DNb<7)Yg\��s��`��1�z�#��(�ɝ��o�omܪh�i����`-��_~��TqC��|^�N�:[21B*�4����O1�0���q���i^��K�m�� ݝ�*R���D������u[dA=���n�����wBL���\�0�(5)�x��*��$7�V�,30�q��M��^�����<A<5�����ů/�ϸA�y�y��Jp��%k��~�8����/�z��[.G��#�}��Y�롬佷Ӊ������Th�ɢ�mqн��3����i'M��Ѣ�p�d��fc4�2E�����KĎ��7Rn�Q�/�%P���K�8�⿇�5��,��S����3 g;�FD���"�H���}	RFŻ����b�0�|�n*�& �㉙���r��z���l�<���b�B*�ҊuȐ�g���\��f��[)��YԴ�A��H�{z�)�["�R�{�)�}�$�!a�Tu-Z&E�h<�����B�l��*i�z�*%��Zmb�z�����x�vth\(��Υwq�as���#�<'�{��ǾM"�Z��i�P��R�G���G51xc�l�0�n�!�w]��:����̧p�o�wٽ��D:.c�Zi�����a��	�X�t;�+U}h�B	t��Y��q8��@­����b����� �M�'5��R��+�S/�6�JL��XA�*V@���PkmI��><�')�%��0�\��Q�c�ʇ���5/��]V`�c���	x�H�ǻڵ�_��T��)��2�l%�~�bDV~�ۖ0fH$fep���2t<������\gφ&G�Y~D�"�[ ���q�8��6�a���wI���O�z�4@�6���"�˨d�����lnA-a���
�y�ċG�&;��!m�7�����&�ypk���4�AK���w$�ݎ��(_�Crq��VW�e�G`T�3�V�⯸ж����Niܳh2~T�͵��݆=m0�e���0u�C����rX�_�.���#_�]�J��� ��5)|b�\���F;�.�b��K&��,.�EJp��bG�;�6^)6y�&��Z��޻�sz'��C,���$�� '�`������w#[7�Ӗ��,���@�TH��}}����k�х�u�ػ��r�p�M(3���4�U���2_cN���R؟Q3�J���~�;@v$~���Z����6��P��K�/,拏&kٟ����m��g`E��8�jG�e���
��?���fyɦ2�H5�O IX����N�a/n��x��
��;ƹ/��L�hZ���z�!�s;��u���uLWx� ���"[�%g��zZhx��� G(r!�`�x���6ℸ�d��'������_	�I�����"�X9�m�ӡ���.��{A^6��Y���,@p���{�� �֦�WI*)�ΦJ���^����+r��II����w�������+O���L���f�ջ֫k�݁A��tn�����X�'�d1,��{F�ts�<�B�1o�)!���|���7+QsY.r�S��ф�޽��E_��'\����^_�D\W�%��	{KI�vҲܙv����eE��\�W���I.r�_�&������� �;���%\��/ՓH$o���++��T�m�(�9.�c���UR<�4�&M����tg����x����5�g&��HeG���N�-��7����O��j[���9�nI�e���@����<iK-�1��=`�[�ш�ng�(RPmn�|�f/�����Vse,)K�Y�\�qBCU���f���Y�ð�߮XW b�C��'�� ����u�vUwI��� R��}�����Fobc��Ǩr>3� 9�y���{����d��]=�ǜe�V�®_�g�y��%.D�p7�,	��)�'%}|s��_N%U0jN�fQEC=t�'����ɤ5��*�W>��r@�Dm+s�j����OY��Z�BA����0B��	�Nx��s���ojB`�S�K��<0uj�@�R%�X�
������A�v�lO�E�!c6�t��ZއK��fozr0���x���
A�қ�j<;�,��Ǭ��^�=Cb�NE�Y��y� {���\8���z� "3G�gk��ɷ/�WS�jt���Tb��:�2�oh�Aɦ������6������4h=�gFB@k��/m�0O $bǈ@��8p��o����C�tv�2���7H�J��z=
P"%z�t�N��[��7�G�-�.�]��Sq��$����'�(�	�s$�*�o��æCH��p��9`�j8m��v[,M��2�4Zi[�΀(e-�&oa�}�蓐���?���D�8T��� ��К����#���}�B�x�YK�y>�Ǖ^N�J�?^�UP��c���L<��oK��[D�͚׬!�������7��HIF����	/!)H�A%�l���U���O'�d����)*>.-=J������f�O!�I�_Y|�Z:��k�m ���L�������:���{\mTA�R��_0��="Z�T��y�̶�$3��V�L��=�"sO1F����}�B4[�J+Y]�L�h�����7A!�%)Z�����Q�u�q�h��bbLP(e�Q��L�-lz��mNn�_�qj���N��q);5i�B>��:�p�y$o��>d��ͲGQ�z�Q퀦O�O�1��a����-^CzU\�7��U.q+�Y�����	Fr��k�d0nf�Y��]'e��ҠVO�xf��ӕ+$��,c�}�{:�odMC��:���w����85�s��dQ�~w��G��{o+r�A,n�O�^�7F��*(�&�)��FUH{&1*��eI;ĺ��l�����4&�i�����k� 0$h�F("�]}�-e�/=&,AK�T��K�?#�t�9�s�z^��w
����x�V yFg~u!�Sԯ��Ȑ����-�ݬ#/l�mH�<
�Vֺ�wQ�5����6��%rlÒ\��X�l#;_M�<~]Q�Q���<��o�]c�=��FRj��=Y$�R�����zT��&�H�zo]b�����ni��DeI:���D۬o]F��f������l絧�������m�^/V��0>�eQA�k`dz�oՑ�|�-�dH�������IlߠåC���$1���7[36Rҿ{�eVi���Kt�2�m8�����1�+�Ƀ��:a�{,���I*!z�6QqO�Y<�p^<A{�FxZY�˾Xԋŀٜ0>4�M���F��q����8��.+�����cܔ���ڑM,yO���Yҍ�Xƥꮨ2���
?�T�^����Y��n8
���iھ8?�˃��<�NB ʦ:w]?�PH��a�Y[y4�F���=����V��I;t�(GN)hC��%�F�6����7|�s<� =�� 	<d�R�ӷm����+ӫ3�"�lc��0��EK�z6��/��X)��N���h�N�^K0ޱd��ѵ8���1����7i����$Oma[���������Pq��S����+�p�`[M?}x��3:�r�E
��C�a3 9�z��t�}�9���	�
��ٴԞ�Ft�=V��EXE�{�Θ72X�d�L+�	�.�cʶ�'(vk�����������o�'�쳋�l��-�y�1B���[�+7<�z��P x�ȱˎ�8������5^"��#r֭:vT��X��^S���m1��f�X�Lc]J�ҁ�����c|p�$$-���o���ڙy�{�ĊF����6��*C<�V��l�Q�����b����Z�#��/�������V��x9'�{�?� �}�`�h��\f��%;>������R����nk�fÉ��v��~�Ѹ�����hȍ��=+ا=m��^2��C���m�1��<0�������O�9�آ�s���kr�A���MF~ц%t$N}|F�jb\�V��4^Et�4�r����A+�K'W��T��	X���$Iϛwo ���I�)��c����{���a��*r^/!��(z�Am'`1ƍ)g�hҧ}q�A�ԁ��К9@i廤�?�q�P�� ���L�̡���o�����Tv����6S�;���nB�����,ƍ��90���p�j��w|�^sͲh����e��uX?�Q��LeK�v"|��L���TZ�,���A���� �Y��\2��T�ҡss�]�y��<]&��ː�PP�;?#�����&��p�q�5��H����h��ߝ���*]���Q���VsV�d|�v��T��u�;Uu,f~�[\c&~WU�+��O9��;�vCp��m�g�f����y`�U���Bn(,�G�&hb*'