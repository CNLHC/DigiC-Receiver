��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���8}6l������3�i|�lST>�tL�%a,���때�#6����e�­�GX�P�<&�_|�|���L�W���b_z�:��j�8H#M�~�6i(ִ��zǓ�T�-��i��5�uB:B��^=9�j�3*R,�}����PCԛ���x��m?��S���bٜ��2�v��:�w&]Í�l����l_�pBƼ�|�Yv|�	����ʤY��$�3���	Z-o�M_�٭Wӥ����@ڪ�U/^���/Y>𚙃�BR��Wa��9���C	�R���~�l���s�cJ�Eؔ3���:L�;1���&�E�S䞍�Z:�I��,>a�:��B�#1���v(H<+ ί9�.��Хr�w��W���/�-9H���LDD��L�>_C�O&L��m���D��s����G�7i�=���\��M��硧M���9����u�C���r, ��C���6-����z�B�Ř0�N�a���>�=t��@ᕽk��3��M�i�L������c4g�p�o?�rJ�Cr�<$����cb �P�97O��[��pL�0i}��:�����tQ���Оb�iZ%�g�-PAd�Sy�,(���~�=��mA���g��*!�4�r���2C���s�F���]��S�W��}W���ɚcDr>�c�8��b�QE�-�'���>����UD'�h��g�%آk����-�3�&�dBM
Ǒx���f�?�xսT��T}K� .�U.��R� �s�{i��`��N�©g!1��� ��Y�y��j��m���<b��s%���'e����9�-HS�R����Zt�|bߍE��S���<D� ��<��{G���m��GR���O��L��]缟�_���p�0�ڡ���^��E�"F�n�C�p���۬F_є��S��))ɣ_˶�{j���`��@SL��b�7iy]a$���x����ذC
���]А,#�_/�[��<���*�����"����6�����x�f�h'%��A�	�N:��c��V�7_�(��
f���d��?A��&�>�p�]��E���ٯ;��+�Ջ��i�~o?*r~��<��Ĵ7uN�99����	iޏ�@�_��7��(�)x\��%�uĳ�H�Q��n�����a�b���lQ?o�+���ԃGB�?�D��Q`7�����Z�
򺙿���R��mX~�w�+
��c��Z��g�F+�����Ը¡d�'� �IX�{J�q�s>������i�D�[��?c*��%�#�i��B:&��P_�DQz�����k���ʯ.�u�Pc�.Pv�j|��N�������XS*I�qq���<�
2�����G�Ԑ
��Itn�.%\��f�c�¯�N"�6b ����^�2��p��|_�C��բ�J�J��DoGJTK�aX6�E4��$��ϢW=���\�҅
�GТ�����������.�ҹ)"�|ض��Q`W���9�f�G�sz;sN�1�@d�1C�l��`��J?��@0��Qn V`\K��#�V	tOA����(�dtt���υ�_�UE����Q1���|�D��?X�L�������䑜\l-��'��=����o*�m{�ǦMn�jML��$[���ï���᷅F��i�`��#�+\���O��$[F@?ߗ�]۔[�Þk0�
:�F]A������ԋ��Q�N�Qz�J/���T�/99\�����H������*�N���,�|/�7Е@��i[�p�_��0a�Y��h�� 1X��LCjf���o�2s�C+�+mc�Je��CQ8���o؝o/�ӯ����4M\k�J�5��s�'�cd[�B�dND�j�-�Q.��GS���T��(f}o*T��Y��v����H�	mF�Y�����E�9���O��8��|�+��)�����^C��Y�y�1#3S|�v�|/y�/����$p}��*�$8#u4 1���c�M/�J�¡���V��?dm*����`N�h��Ɲ���pI�{�-_9ڂ�;�aF���K:'?��@Z
��H����-���|�8�	I�~����<�z{
��q�Q�KcBli�d<<�w� )ۜ��&�p�!%U��+��^,>n��+��1� �U1d�����O��,�i����7˜Af;a"b-�'~��g�+e
���T4��R�0�#u�ۛ�ƭ�nq(�-���υO�ʭ.�0�qjxsCZ8���V��'�ƭ���y�U�e�iΈ�&@A'֗E��{�"��&�z�xYG�ͪ�-u�R�����W��0�|_ ���D�W��wg�_�|wR���u�fC���)���W�$�]�D��*�ƕ�4�����w'�����0yBڇ?���g([U��t�Hơ��%f��O$>��h���`�p2�3���ʯ"af_ڏ�WL�i��T��ĢbIҁ,l�r���)>�o�Yj�d1��|U*�J\2��A혹z�k$�s��B:��T -f~�[�BQ�q���?i�nT���{Lه:��Rxঝ��;N���q&�`��v�qS̪@�2^F�3y��� ��p��7[��#��f� +��"��m䜍?xk6Ψ����Ѿd���Y���ZE,��>Ē��d�$�~\��[��-ooG����z�g�h �嚧���B"S1uۥ���<��P�4�� �/�
��]�ctPҢi`�.���i�6޻�Vs����^B?����p'�ǬU�hoWoF�5ؠ��yG][�a�m�_B4ϑ��!�xMX�c�S�++�lF�z�m������I��������0�?"P�����1�J<X��4s�%O5�� A����V�a��10>�r��؏ZY���M�Ő�
g��6�V�ؖ�u��($��>0���ٰ��0���26�D�O��m��h�#����z�ք���'�|~/��Y�|U�W��5�T�AY�9)���\�E2����8V#�M�~v*goC��7���(&��k+c��)�0W���}S��ZG�ءʱ���QM�.��Aqq������Tͳ�O)��?c뗜��-S��؆�w��xrPu�[�2���d$1=�HAW	�1c�ʘ�=X�s�����KY��Uww��4��^�EI�*;jo����(�l�+����1>�
���2��cw�CY�������Vͩ�,��l\��̉�\���x�P�e��v�7��jbϞ�E���p��Z��!}��BH��%S�Xd��!�XuWw�.��諯��'��%Z��Q���sJ�О�ךԟ�.��ˑv�l��Rp�κX^Z����1_.�r;�?�]^j�9D�R��.�VN��8P�	�;߁�ȑl}3�U�0�2�,����t��OFYpz���)yC��������s �XW��rg-�|������ę��=��%a4w����e �Y�d��9����g���{��4��豘�M����x!W g���'W��S�>� <����X�����d�PQo� �M��z�8��fx��l��A���)��x��k]�AV{��W������D�"�%df��OFnڱ^h6����B"���T�oA2U:F{il�D�.��ZD�7֣£2�S��M��z��m��S�o�n ���
����A;	���ً���l�����k�Y&��]�E1c	Le!a�+��b�15�Av���U0p 5ZվH��/+��'�s�gЮ���m���Q��6���i��>�e��	�tN�q��jmb�^�K�k�Ĺ��c���}O����Z?����C9�/-�lJjX�ѣ�n�ōd�S�ھ?��B��ӤN+ Rz<"-�B�%i��l�M�����;g��&�(1[��x(�sR�sv`��C�pj�CҲzݻ�?�71"�s�힕�n��uc�6��T��\�^�Z5��#��&`�{΄&��s[`\��*cs���N�RX@�h�w�|�L��w�9$
f�}[r��eRf�0 aK[���h����������N�FX�4I�Y�� <���90�z�K,�}=I�J;M<�UOX%a�%k5��u)�
�*'*��]F0Nl)��a$��J���^%:�-�ޜ��G;�<@6/�f�F�[�j�s�e���Q�nv�ɩ���:%v/��
5̍�r�V>��S?�r:l�����A` ?�%�=:�׹� ��d����/�C��41l��޷����s��5e{����fu^zמ�S�h2r�ؽ[W�,o�����%�sng���vibF�T��O.��HY�(^¦�E�ǁ��a&�$��	w���4K�\p^d�@��:Yg���7��+�Z�^����c6�
����=R���@�O%�?��!�h�"Q2|��c�Mh��� QHCbL��+��۔�Cί;�������'�L��*�F�s�A:���5Xa���XU�媄��0ϩQ_4UH�78��l0�g��J��~s���Ї�dKh���gBl����p��-����6PǼ�"ݿ��\~(o�T,��fVY��E]1Gݰ0�!܋��W�W'��ڦ9�ޓ�ޮز�gZ�s���������;w2�������}�#e�œ���4�*6�u��r���O�`����=�I���<��֫�^���=�K�6�:s��9cd]�X����L��i�~�p \Gl�yxK��C���������׶"(%a�qWQ��&n�~E��j6j]����q��s�!%�m�T��<X���/�����ɱd�x��8�<W�}����W�?�LC�]Mw�vs��M�HJ@cuE�r�n��
�ʎ�Kc\2k�]
�f ���)��Г+\�ު4WO�R9o*緓@!�I�Y�L��5����Nv��T�iy7��,��sBl�3k��蹆�p�נ�F�s�`�6�YvT���{o��%wY�)ZwR���r����Z�1��Y���(��j&�dq��(+H�L�]�ָ$]0�"���w󉓁>ۙg;@�ar2�sH�k� X\�y�8s��.�cr�������R�v5� ��ퟆd��!��zb�܍�8_�>�t�x ph�Aqt-���
9���*�!�z���K�����j��뚖S�lT�s�z�r�"�^J�sp��k�}_�Q,ӟdD(��3I�̦�4f�w�	��� ��CJ%�Wv^�g�u�[%�+�!q�aC-���n ����"���ZʞŻ�u�<p�N��R�jӣ��	��d�K-*n?ř�jA8R�����,'��ꑨbjJ��ɤV��?�%�4avd��`�
��J��GeH����;t��R?Ah���a�/R�d3��}e.��-�����|�,�pȎp�wy��:���׈�o�IŠ���M�ɼB6�;��SE
�)%�cTY�y�\0��'������~9	��0(���,a^][�i�Bɹ$��έ������P�לk��0{�O��'g��׆ X�!хr�2��ټ�ZsY�&̻<�d����	h^/l˺�z��Ѧ%S(7ڌ.��?*'��38�KD<*� �}�ӝ��.��fP *Ӵ��㒔��XL����*~L��$�$�\���)6��Y�t�N�<��`�>�@�>=8�C�WT�Y�J`��1��v;Z��̂8vz�M��u�Hx�zc�n�g�gsg=�����v YQ��nĵ��p�����>$0��
VZ����Q���0'j��bWh�E��o��M���7k�q� �֎y�|^vq.y<����@Cz;���I�'?"$ZZS��Z��L�
��/,(�ϔ�]H�޿]���y�P�zu�>0��jF� �zwu��՛��U��Y!�a�����`�z?�ȫ� �e�䚓$�wJ���]e�𓐿/�g'�PNBD,���H)��qX�-�IIuz�ެ줽�Ss�B�u��n�b/�~��ᶚ���v|�lg��!�MR��0�e�G����d-�7�����_R�k��&��7��s��G(@$o�F�y�V�-��h��'��챑&�b&.~!�i�{^
4{�Yw\�<#+K��j���>��ϕ�i�Evtd�㢊��.����YX6s�J�����]oFK����ߑ��\4xM��817ڑ2��ʿ�<��OL�7a��} i��?]H�b�Ђ8?�{ͻ(ײ��̙����6�k�:�F���� � P������j��To���XJ3����[+��l]����=0�H8������(i��JqJ>���2�/%ٝ$to�����|�lYO	1E��Ӓ0]�q&f�����uJ+r&����r�������8���қd��	 z5��	N��>�f�㞧J�yW EU����"��V/F<?� Ma�M=����w���>�8����vaNI���p�2���oｭ����'���d���oV������@ځ#�"C�<�_�z=�N�%�3�������cu	���@�`��OZ� D��,�@ '�pu��Rs�P$O�4i^��l9�d���.E�8�{��e��hQM�P׌���m6��_|)�ZkP���mSs���7���at�)�7�K� ��8k�5����=�j�r���hQ:���E]%��sf�x�lC+��C	� ����\h�|�y��R?'#���19k�1 ��|^���p.����O��
���xq֋��L���~���=�E���Ͼ�Hvn�������y��v�[�IHx7�fW��Q�1�3*]��e������X��V��f]R&k�1]��HL�TJ�a@%��@i���=���V#sv����DPM���Ƃ�nPp�ݓ&�;o���-����`r�v�8���
L�h0���2��S�1i4���aNmw��՛/ *�ă�ʹ��~-�(���aXi?8-xѶ� &�J��MMl=Q0;�kw �9h
���5���Y�o��Nܝ���yN0��J�CZ�s�i>9������˪ˍ�W�V\� ֣�y:Hڇ�_���	���w��P��;+"��"�[�Q�+9k� o�HS��Q���z�Z�6p���i2l�>K��:����ן"��ysR /�n?�bݻ�%�)�V�'dؽ�t}�4�ږ?�fu�5��}eӊl�e3X��,��-FT[d�p:{Ϧ{���A�&E�k?xH]K�Tp"J��3��Mx�dȹj�4��DMV�rœ��W��18NK(�*�+���	�Ȝ�|����X.�y*p����
�i���Q��_
�R",ЛԬ���W��,���:z��{P�7G��D�����b���n��u��B[7���~�{u>Y���	pd��Vؙܸ��@�6��]� S����(	�bu'���RU�	Zw���γ��4����?1�o8��DW)y�n����
�o��u��c��W 3�E�S�V�*R�pq��j��2���:1±I��ov=3���	�+N��&댏����?�X�<W��dK,�ެ��&���q����]2�@3Ӓ!���a�P�?��o|���a�%Чo}��*���y~{v䧔ү<�B�IS��UE7mQ�/��p�ϙ,sNG�sa���R>�E�A���+t�2O�'�A��y�p��ĦV��2
�fq�p�}PWC��{"�C�E[z�_�vT�7��u��w{�U����6���y
8�>����ĸ�+�y�-׉��i��5Lh�������AŞ��o1>!�D9�38OfҦ�!�lE��[m�����l���^�|��[�B�l�����df��a�K0�7���		�������S9%O�#�A�	�eg�$�/�V�;4j0����й��ץ��O���k�my�y�ɐmm��~;���-���T��m-l���g4�4�D�����8~��՚+��\p�{�����
���Q��G��cN��`g���K^��67�<?�lT��:Q��i�+��a�Z�B㚚��mM�N�'�"�������@�֗1Ao�)�k��$-�=����'ւՙ��G��a?>��SJ��q��G�����%�����r���wm�����[e�#�<���}R�>��|�-���UV� ͭ'�p�{R}K���J�g!On����=JCR���]�	�<?�+��Ă�M(�+�a4�1٧���Fx,�Av��=�Qk�'y�<𧙓's
l�K�[��ad>�K?��������z[ڰ�X�c�2�����L�������e��ŌG��]VYD��]Ⱦ	Q���T����7T?�I�G�I���� ����S��`*�W{v� �m��?ǘPQK�Q�`��\�-V�#�+�DM�N3R��
� �Qo����F~`�D.5�O�ع�bq	!�zV�'�7.*m��1A�D� �v(����6�I�(�ȗf������v�@�]�el^��.d��BB�r�,G턙�:�:]���T�No\�,G|<G��x�4?�;1����| �#L�F�ÛP��GQnE���HXl�nNJ3�MSi�,�X�=�!�1v��bk:G��Yv�_	���G�Gލ��e���b
�7)?��6� jnYl�~���>�%�|v`:��]��g����>";P䉬����"8V��])�����H_��鿆���j)1bud(��UK���O����Snq�τ���\�÷�9�P�T�XFE��#��Ϭ�g�g��\e���.��_*��{!��|4f�y0B"��:�E��L��qg_镳t���N�u>K�V�2����2x6��v��P-�`����;ɹ3<��?�\� N�Ŵp��a�K�X�(J[�h��(�>��  �寻�9x�{>u����
Oư�D�w9<�� ��([*�]���u�l���c���n��O�� u��aSa+Y�7n�f�iQX$+�i9C+���#7����@PT��H�sa����m?f(r�!�ǚ)��w�+��1�Ģ{�!	�d!���:�Xt��8߈���V��Ap�� �/�OJPר3^��mQ]��_���WC����L���m�n��pO��РU���x�8�hǾ���PJ���b��,��AΥ�`��O���x񍊍�r['E\�Y�]�UX��aS��#��Ķ�uK�l�a%�	�
8�k�*r�p�`q~�ǯ���p��+��/�`��T���@�Om4�:S�zV
˂r��@��²��˧�{�����*!0`9��7�N=�`�=Pڢ
^�������d�z��-�)B�B��-�p�M����Z��PIR@������`�k[�fU�?�`%�)פku��|�R~zB���E�Y�ђ<=�L9-�����	S�il�7�a�X��q�� ��o�]`����\�dB\m���H!&��(�Hx�5r�7 �uc�tZ�!��C'F8U��İyC��`ax��8>��ռR�O�J��{�oO6�u����<�6�O��h}�P�'�%J	O5���_e�1F]?#T#��:��7�k��2�2.A�B쁎*��cbO�S&�=Xc��V���U�@�>��w@��Dw�U;��
��-�Ed�3R�n䖯���N��{��=sb��H�S�����[�Q4�FY�J"� .g�� M�@��D`5t�T�l-���G��:F��b�,�8���c�|�R5�L�� <4ր���iD��%���MR�iR>D�괿	tA�[�i1�y
�����"�e����[I�!v8�	A]���~�����|�LU�l0��Q�ؼ]��ڱX��9%ǣ���|�Fx{�D0F�G2'�lk�p�]je�Aq.��S���C�/���n��$�1� /I�����%r���}�B����3/lD�Qo�?�2K���>k�z*+%|:{=C�,(>P6�I�fg[�k�ω�t5�&��Ś 7W;nÅ��9��#�6�<�Y	NE׍���k^c��ʦ;V�:�W��Vɝ�߿��v8 T�[Z4?�w�Do1&��z}�Kur��%Q�J���V�h��p������s����+b��Z]ʈ��W�@�8�����.��lc:�ksX�8-�eI�D�^i:D�~5�����x� �E��ݑ�b�i���e
s���(!jK�%;j��UBM�,ʯ�lM�Cmvr��� �����+X�:�p�;e����P�����g���GZU�� ��� y�5L@_�}��[���̪B�!��oI��,�6<+������)�U�1��!��*λ�sd�r	��n
��U���-7�ܗ���� ݫ*����wo��[�};����E4���l_H�jɳ�R/:f+ui��Ք�]K�Ñ�3�Z����=u�;pP�tcλr�Bd�!��l�ۂ��㺔f���؈�q�74��FF��P�%�l�fYHt��/�Mx�:�Y�b��Ox>7}?R�!D�s����Y~��xK�*ǻ���(b���~bX�ǎ��Jm5�I��)���|�2t`���� ��Ɋ��0�&C�9�ݢ�jw���D��H( )���g��v|�@ϴ6Nz,�jK��D�Q��]�H>�(�����+��i'w���xz�Ϋ���:��UR򰍔���:c�B�2��):���G�,�����<�]1��U�{4�H�F3M�!��V��C�a��
m�5,/�!P "�#��;p�)?�]��(�KŰjr,/E��q�n�z
)���2Ч.�s����
6	�������ߖ!U��D� ʺ]�F;��ɺZ,b��	�,�/���P2����SG�;�A��� re��)M�Bt�\�)l�l}�Hy�|�:����}y��@	��_�C�ѧ�<�w<��F�5Щ��$iˬ�"�� ��
_��~:g��)ݡ`��V�i���]���eO�td�V���c)vv��MI�[ҟ�]@��\G#�~.H�k�S�h��0�ȇ�R�����f�㠢m�aw