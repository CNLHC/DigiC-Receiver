��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� �_���>h�7N��{�HD�M��3�9���a"aÿmK$�ݘog���
��)�K����#���6�292c������/�I �K����N��j� 5�����lK�.j2&ZT"v#��jQ��c?1���[�����fG�#�d���ρō����+�N�\F�o�y���Io�������y�q�I�Y��m3m��?��*�ω�CR#�M�6��d������qsd^ ��LH=9������;�L}:���I�Li,䅪E�A5I��٩��L�BJ�>�Օ�Z�7U������-3��}�z�1X�kZU��>�M{D�U�����A�m'm>�l��:$��52��O&"#տGtJ)to	�i<��Աhk�㣷�[.z�7+�yM�nyD��t6�Ԓ�Xe$�k���pq�i�r�9?��>k��*�\��7�����6#6u�F���{��:RS̜.|�lӉ�i�S��l����Ԃ��M�fF���3qB�r��02��{X�l�\��wY]r��´ӷo��Cׅ�g8t��gm�KO>��Ƨu�.��P6����Ep}r��W#�
�e7W��)pC�R�{��x��_�.tjM6����T���F3}��>|)G�^�s���/��cQ�
vaPDܡ54���aꎟCXC�$�S�U��?t�|�����W�Э���<�I�e>����m2���KΓ��	��[��`EWN�.�&�;�u�U�?}EO�_���['����L�z��yZ�����x�I�ͤ��	~Vt�eb�gG"OU-�W�8��*�����A��ꑵH���v��T�Iɼ�w�Cd���~+IO+����(�Ps�栍p<B����([D�[c��K1$xz��IFe���h�W��p�J�od^R�CTKP3a�_PRl�|�u,(��l�F�иqL���n�fk�J��n)��C:K�X���3e��oKϥ�J(��}��ThOW�_2/�M?pj���-���A�t
��[��1����i1\�=��d>�Z�W�<��6x�,sf�̧�'0o����@���=@�3��ʃ�b���Fk�P��"�z��,�_����D�����s�ia�{W҉��g���{*g����|�x����F���v�,s����mN���f�i����H�ADL'�r�f`f�.�:n+F��f;�gN�9din��L ������!%g�{}��<�?n�ӼP�l�+��H�۾�4����f��$����������tI���ゕ��Y6�T�F�ֲ����H�pse"�r�8�W�����%��#Lo�T���;��{�amҏT򧑡�li!\oR�U�ᘂ��k�����p����7 �5<]L6X�x[w7�K�K��+��Dܣ�r�w\O�����f�x�<�U��ߪ w[<�3�^X��>.
�o!�.�!��.��Jzz�ġ�ucw�s]����]G�N�t[r�N��υ�x��D�Z)MJ��v�P�yB��m$�I�B3/�F�!�D�c�U-%�:,l	6b5�o"���vv'qמ���ga%���$fҺ��o{��M��
 �M��7�J�U9�5��/>@4�c��1en@  4ޞ�,`M��F�2��Yj�K{\ ��pd�%quN�;!'K�(�X�0���H�=�p�.pKԷ�Fjk�toK����j5�cRGM���O�y�����zk���wK��H�vL%��3�ꇘzZB��~X\T�Q?\υ�n�M��W��%t"��1G/�$~�%�j�ns@�����Mm���Àe\i�+.���_��������b4n�5������E֓ᶸ���t�^��I>Y�[�:�>-C�-)Æ��Ҕ�]����A����OJ��`�D��D;'�Km���0���������&>}1b�ƑU*�� mԒ'H�>={��;F���v���g	.��8����ٟ7�qX&�X���m:��g�	�d�F�S�^�f,��몊W�ƚ��f�9��u+�xd�~v�f83��*��o�A�������tʨ?.,�����?�t�h��C,0t�i�ߙ��n9I�:E[,�T�Ȋ�ɣ6���Gq�E\�cg��z䠰RF����C=$�s����"�, |{j�㈧��`R��p� �`Z*u��HZ����ן��@}���,KI��/͊X�c��~���;�jL���n�k|L��T�Ĵ���tq��:%��vA��0�����t���YfM_�^��R����Ղ�,����j�� ��v�5|�:�]D�
�&�OH�"6��w��ӮF��|����$�H|o��N�)��Œ?r����5Y��Z�� �%򂐫9D�y�:_fra��	M�f�ot���I�l�H��r:�m!�� ����Ox4��r���F��йP�o������3�?�k摚��|D�����#�SIߦ�湱���]ǭ ����1a���@���y��|�Dp�o\��ɫX~|bC�\�q���q�s@�����W1./sr�>�tb���*�
	��̉�-%S�j�����06��/�PF�߶�ܤ~I��W��I�(�N��\5�*h�f�m��I��O��V]:r�
��[uQH*�)�U�%@�My����o�Hèe�C�.��V�E_��3�U�%�����/�?~�ms��q��4��umȌ�ϥ_�/�"6�F����s��eTe�$������~xW��2F��k���,�G����0h1��X'��g��2���^y[Y(���'��_q�f-���$\ԁ�EՅ-_�׉�wu,���Fn%2������r��uK��C�W5��e�H���Lľua8�u��ke��'kIe��h���!�߰@/��jx^����ȢD�kD��K~�16��+���zm���w-�꫞<I����󤋶𹩐���@*�h �R�������CzD��X�	���@]�J�����]�.@�N�se����N�5	�vՉ��fS5� ^�3?@�!7}���A:�P
آ0K)��)'�t��J��g��-`{�&~�QV~�Ma<��c8w���t�y�0!��Bu_�]�ߗO%GճM�~+��l�T��j�պJ<�
�+4�S]��!�1��"急�+#��D Nd�h������kC�8V�����O�B:^Ũ88�t����Ƀ�I�q;V�u
�����!�U{�	��;��w�oe�+�����&��g9,|ޤa����谍(�X^��d�6Bة�r@�)n�i��ѡ��R�9{�_�5��t��=�y��eykk^���#t���?L,,Mo�Lz4k�R�\�s�ʨ�M��	j�CG%�)_��N@5g�o�x7��6� $���tD�U��FA�UX��*M��5p�΃Rc�����6D1���7B,g9M��k.��)�� ��
���7�E���|�J�zAI������5�ǟҿZ:�g��	�D�c*]������g���.�:H�غ�)w�=j�=�1)�F����)P��H_��d�iG5�k�:$�gXd"�p�{�[�t|�ޑ5`�n����}�F���8�I/�őVZp@ب`r�`dm"Ha�#���z1d�?�e�O儷���qԛ|>E
�&R:����.w�TWjqf�.^���`���>[z$�d�F�o���o�-V"Y�9~j��Q�n��Е�ƞ����.�H�����(�� ����f��{��B�D���];�E|Q�
a�feB�x�����:��3�!l���%�~�r���PdOP�������I�y*�1����aV.��pp��]�$"�h�W0�<wɈ
���k#e��	s؎*��q�q��^��?�}w1������kЗg�W_0%�A���~�#;{ �pθ��Q���Vg笥��%q����(_��5B%�F_�J"���@�+�M�U�b�~JW���c)S@�P��n�Z��Ǒ����x�P�[�d���8������Ăy���b�x�*iIT�X��jO��G���/���y���9W�|q�`e��$�a�����a=��E���vfw#��}�j�>c��x�J'�\d�}F�!�Z��n�O�K�
o�h��G@y��� �$6*@W�18m|x��O����X�x��T���a�^v���'�$�����q��W�:v��J���K�����r�W��#�<w�V�veMԦ�;��g�k7Ouu$m����	�]��c}z�A�ofE%ce��D-_��Le��gO�K�Z�/�|S�^�o���F.�����=EpZxO
��t�Sv0'�i���&}Z-S;s��:�������/�O&"u��f�j�W`"��*U�f��-�8�,9������@_2X>��6TDe�����{*1��x����G�]��JkӢ��G�ؿ�ӧ���(�+C���K��s���ED���X�#�}��p��-7��Q�t�:k��GNA<.q	�e�i�?����A(��3<�?]A�Ȕ�'4G�����Q����-�:�/:�++��N��s���6|b+����^�ZwӜcs�Y����^�z7�c����W�Zr~;�?@'�n�� �u���F��'E�LV��@p�V�}\G�<7Z����z��D��+|��RA�wLJY�r����z�������'���c0�t���\���-�Oʲa��,�c,K	M��	��FN�����_�����1����\�?��z��MQ�pW�Q��:�`S1Y�Bd���|_�vK�{�0ݰH�J�%�a,i=���O��qB���pYqC��2״�(�7;�;��ȓxu����l��kM�=<�g��W�f��cC5s�U	������ԓ� �DZ��k�b�$�6�M���i1�=� .������� �j%xn��t)�#-�W���8�h_��W���w����Hϐ�i���w����&Y	�z�{J�ʸ0�1��;��!�D^���i�I=p��̷AtE��w�f�Fq�&aDX�JAh�lJ��⥟o� l�w91��hP�_E��`�	ϡb�K�o����1rhD���B�Ҿn��5F dB�0�&,-ˣF3v��k�7+;��k�f�t�O��	�8*z"��V��\e��Ɖ��B����Һj%�����<��VJx�<�0�����vso��~ͥІ0�7�F^��!��h��2��cn��in2���e2e�^�k��	���V`��i����v)�#$`VA��R�P�[e��R/+."}haK�A��nM�S�
^��/���_8���o/Z��U������q��X���$?η�XV	6m�1�em��:у7?�ԁ,�N��tp����q�Q��Jv��E>��S�����ui�C{��~_�V"W����;�����@��ʭh��͛"���)sh����\�'���2�LI�韽���N������Du�vُ�as���Q.�K�d�6�s���[�Re�TC�9�۠��g����'S#{1��ogH$`΋�8� ��g0���>=�7cB�.�
���>���?��K��ǿ���W���#`Kw8���D�w1�����t,�@�2rO��I~�Ki�Y������d"j݀�Vj�t�I�x8���~�95�<V��t����aR���eÄ�"��ER��/2_p�=�B76g�Z؝{��G��ק�����ᴦ����9<�-I�(ms���p2�&|�k�c��;Dy<Tx׹kz��ɓ��8�+C^0��٨$�}��O��B���i���L�Z�+��װ�v,��㿣���8�Z�_Z1�Fs�p@��-W��-_��#�^/L���p��"0��j�)J��U(�2�pRa�b��W�Ӿc�G7�jBK��f������lH����|)�lD)���?��Փ?1�d��%��#J+����m{�w��5�E�1��>-_��t�:5���W�)�c��OtW������I��һ�1�1d����6ѩ�JM�A��Ľ�m�-���$�}�8�n�J��HN�Q�{w�d��i��i�;y�O2�P�

�G�
�s!������:߁�� �:|\N2X�S�䤁�Jo�����h�6y��]0�d�S�Η6[߹1���$���i�����C�o��~�չC�g�辙�0�T^�B�v�n�Oµ������k��l�MJ��Np������Ɍ#�_'�#�!�k0�SCI�r���Y7_�K4��p��[3�p�t�dQF�U2\��>�W�{-�nk�+9�X0�e�%���|�$m�s.���8���1-�[߾��yy2��h�.��r���jԈ���O�s���4���n�ޝ��)���Y����C�)��(�So$@1GR