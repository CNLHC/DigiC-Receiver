��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����Ʋ������� =��f����>�%ʌX�]5I�Е��V�!��~�jK,&/��G�FA�zC�t��'w�ˌ�jP
��l	FE��ͪ�b,�&��k��vHZ�3�@j�C?����Ć���i�S�~2�D�U��&����� R�����cX%���@��p�x6��(UD�0UQ����i��@d��E�yЍZ'U�q���{��FPM@�5=P��߶��.��i�ے��9��kx�"�
嵀��*j	8�������.pY	�T�d"��G?/!7}ز�����	�z�F�hӻ[���������� .���aE��eP���]9I3��ט<g���m��	�Pނ_H%��А�L��n�X�~;FbT�W�n���~�_���`�3T��8���r�qsAp�n;J� �^��1��2&��Y�Bo��~tL.QKak*2�����٫*��@��K�L���93:�0|�$�h�x�c�[��8�g?]/�H���DV�A[Y:��ݗ���1���"ء�#'�R��m����� F -��̃����J�y���y��=�Ґ+=�<m,<��1�Х��Ņ4.�j�mMO[K�F��Mx~�_���.U)Q��/'ӗ2XI=�X��FbYyI�}Vܕ�߃����A/nO`C�*]\�)�k����@Jr���4 9����	_�R2����l������� 	X[����g%�� ٯ3���L���.
�5#�n����0"�I��0P��Θ8i*\�R2���V�`�K��g��O`=�%am� �T���?�iz7��b.05NLւ@V���?�m
�&wLz^�i/��$:& �*��:xZE��/���`�θv���i<��}���x��W�ƚ�u���)wB��62�(b,�C�P_�ēhಮ6�����\��'�[�����z!�-P���P�Ǚ��j,��A��,Hn��N��J��L�i�$V�{�(�f�>#H��cAY��CM8���tD��?��=�F0c�i8�<C����O��ӟL�̱���਑d��Po߲(� fUGkJ,�^��x
t��է�RY4�Ϡ-��Â�ۦf�����v�|D��z ��}�t�آDx�*��4 N��6N'J���]�c�o��b���(�F�֒�^t�0��oa}h�@ӄB0\V��^��E��[�%�>��>��G�H�E$���m��t�p�S��¡�*���u�eg}ŵٵ�K ��bcQ/w�MɁظY��&U��(gO�S><��u&�U+�,#�c���*�'�r����Z�"�(w���sv�ڏJTx�������W����BV��-�3�/�w���	���)�Ur��Q�{��*��gO$,���, $�Z������)Y.0o�X	��r�9M��E�d�Q�EY��q�k�s8h��0a�^B�gL�|�x?�p/��v�'c�(���+������N��Ej)����`�j�^�܃s1?�2�7�o���H�_,B�q�q8�Q�s"�]1+ H�����3���T���;R�q�i{����MO?M��+LF$���'��	�!&��*ޝj��X���ls�;gu�#0� ��4سj����a;��re�n���n�z>�h�]���ye�%L���U���dcq�F���ø��H�3\"x���$�n�8=� �\R4���P,&Vϰ+!B���7UbS 3�/7�AѬ�~��u{h4U���dٜ��*]�