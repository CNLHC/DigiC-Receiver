��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]Zɬf(�'4�o^d5��o5�V+�����YE�٘tv~Ҹ�5ѿ{fL5�+��򕰝���.�8�v�Ĉ䡹����>Q1͛���]�����6����G�W믬��RV��i��(�]Nxe�P'���IB]M��ֳs�]fd��=�23gQPn�i�p��5�_A�ZM�d΃44DV�j%F�0��W�A�ܴ���S�� ���v�e;4r��M6�z�;�5w0wGi�G�g�'�L�*��܀������*f�c`�2l�3��w8P08;�@�U҈�v�����&0��G��&DkJ����DMq��/�f\SswL2�X���hOi�g��!}�$wu��&	����H'+�'<2�l[��N`��X���Ua׵
>�#v���&�o����Y(�/C��>r�����r;pF�%0�U�R�%��o��Blvo���%�d�~5B�y�戆NM����6��{� \�`e���Kե��ccDfcd�EE�W�:�Xr
��|�G2@tT�������"��d/r��'F�����tt`��⫡ᚥ��$��@1��ێ'��y�}3�h[�j�7�� �#�&�c�����9�W �OJ�jI�����*N��������rSޥ���6�le���,"�s�<��͉F�B@��:���~�0���\c."���'mϲNo����������Q9��V}�ow.�QӋ��l�ԋ;]˥l���_�*71�_�\I����Bȷđ���|cg�E��k�����d�4���,����;j�$��\17J_�4���5���S��*;؎���.H:t�	���_0O����!�XR Y�N�3��$����m-��i
(� �ҷv�����U��
H4��>'n�u�K���5�r�P#�����@��� 4^Is���6A	��8M<3��ꎎ�[	>�R�!��;�
k��U�.OA���������B�]i̴���[�B��R��)���2t�����L�J/׎��?��3t�����)w�GϦ����?/X�"�7.���xȧk
t2�w|t�����Y�5 �0�yޥlg��@߶��O��]�@�ZRnw�U���"�AǿҎ�k����5�,�y����N+y� #� ⏭�3zj�}F����:�-���:��@�:�2��&5�܍���`/JO����@
���{#{�x9�Y/B�
�@�)B)$�U�c'�PF�����Y*����V�P��7{�;��2+IZ)�u�;r�p��2��4F��2��j{ߺU�J�^B��n3v�Ɨ�WE=�k~���m�/�E&ٱ4iMѐ5���JU�����N��P'��k�i�s�OŘ�2�+qI�%@�O�Gh�$�b.A.��)���ZT�.�C����Fuz�ߎ̕r�]y���m����_��_���e�א����oDz��%�Yv��R��'�7'���A�	�7!p��o����}S���M�zsd����ʏ|�7�0��RxS����yj���)�� ����-Bs��Fm-�2w'�r��	
XRoB�v_4l˓h=��d�-�m��&��cV�mWqQ~�s#�ݣ�z#C�)	ų-�:�������,%0"_`��{k���ه�4+��b�dۢ�O�+�^$Y\��'�9�#֊��Bi|M󄖘�8%ﭵ6ʚ�;�4X?&�%������f���E2�EXR�'�gxtu����� B"��܂��>��BW��B\�rW��I+a���~�{MBEI)�Qkb�@Pd9un���o?�>�����ڭ�m���i�w��S�}�,�4���U�淝,����d,��0��J{t��%IJ\0��IJ܇zw5m�e[�)=��?�/���Ao\?Hf�!�I��w�c�lqL��U�U�7��zr��e@(�ܕ��##�7i]c�S��yʃsJ�����$,�o�K��蜱��Kz����L|����Z��RM�j?,]�Ȯ��i��p�J���6s�R��*�W}{��#�� b��c�r�1E�"�`��i�t��=>z��̦DJ��a���}|��v�"iY4'j�a_�kp�T
P"i���	�RSݤLO'l�G�<fl��ҠT�	� ���Aj��La���=T)�����tQn��Zd�A�x�[%��ס��8�������Ș�7@������&"$j�tx�eO�r��ɨ����s-���  �B|�+K]�F���b���Qo�A��ꞟvF��'�_�L�+�*��۶���4m�:J�w^��Ƿ]�1�*�&r����[0�C���G�ܚA���5*���!����Q>n�����l�HV/Ѫ��0\��H��>� z��{O5���2m����?MG�,N��'DF*��y�?S�+� �7��?�wV����EP��!��eu ���ɖ74q��D�hu�-G��VR#�Zâ/ �K�ձg'�}�A���bԈ�^{K؅T�V�"߲��gB��P�U��@듄��X���t�!6ô9-l���ay��: ^�&T�*�����u�����ҬX.�s�}� g����m�!�ֆJ��g%-�cL��<�,�Pp�W"�"�O���i�:�M&
t��vĝֻ~�ҡ����Vھj�D����b\��*�I����臂%��R�K#I�<���g���ER����I����I$gd�v���c����Kjy�G�ku�6��B㿱�� ��S�g�Ʈ1=N�+�Io'�EJ��4��IG�~H�e8q�$���*~x�&�h^$.�y�7v�����Vw����"a����L�R_O���H�C��Ė�1r�iv�ק�&�k��3-��k������,�&�h�@������!i�6�� �����y���;%�7�rݍ�㫊ʊ"���.-�z�[W_�b#�iFΡ-N��d��	>�����ұ<SͶ;�|��*2�3a_��"��Bd.���㲜��^R��V�$is�<ur[��^(L�A��R�l�Q��q��Ƒ�}*n���+�#�����2[8$�P��I<yA�B;*6#G׉{�|D;���>�Kd�wX�e���b2�
�.�]����rI�7�bgT�E����s p� `��X�owDe��D1�C)%�A��2n�
o���%���\�	���&�"���f��Ӫ'uɡ����KL���o0�޲}�c/�'��ס��<��ݹ�qi:Y�YK~�d����f)�-M��ݦ��y�����	g�@�"p$�@4`��J�sn�fß�wg=V�B7Fsݷ"�L�(�9���"����w�Y�Ϲ�k�
����m�C���_��u_�;?��ُ+ЄP�Lz0��jU]m~}œ��s����:+!���ϑ��-�#bQ���H�&{Y��́8{uç*�֐U�U�Ki|�-�$Ĵ섻v�����$�Z�O!r�]֤�X]��٬��ms���v��t`��9�zh�x��C�Owv����G3�����o�f�qF��Kήzb[��gN:�MM΢������5�x�I�����j nj&��>���B&�5�%O�PQ'Ư�(����p"G���yl6��
�W�xB��+U{�cc�LW�����"i>%�,��>�M�r�~��:��'(36��Hf�^����6�W�avWr�+�h\Bi��DI�����)�h�`���&~`�^k���T��FM�"�]y����9�m,����2�%9HiU�e�=��Ȫ����F7���B	d���l~�����6����c�e�d�=Y�2+�Ceh�^�Bpo �I�����x�w$�ȝc��Gr7H)�{�1��TeD#o�����|.Wc�wW͒�����>B�@�\�,���N�����P�4����i9�9�m����\�o��T�qv�Ы3���.M9���Kz��{PM�1?���ݾw������lq�h����< 9UX�r����ncE_����U�(i�tC!�FC�M�4:�ͪ�x���qe;,�n��?���q<�+���"���6�#����;?���8�����6��hX#nމ8��+�94�pG���_��-0i ��X��_�e
�ف��2�����߼���݉���5R�/M��#'�J^Pk7���0\�[�% >[Owx��å�ow7�	��Sa�
`�X�>LY�����m��_S�x�s}sĐa�����Q?�3w��;,U��Zr�ƽh���襷{"�����}8�/��k�w4Fu �u"y�0��0��D`�9�I���y@�]E� ��������<H8�#J�;�i��#�Gʋ�O��0��b���~ %��\��Q:��/����z6�����4-.�b��5T��Fg��ǫ��Ӝ��k��@�_ =��2�F>�ֺ3�*Zt�zG��C]>ݷ��������޹��M71n�|�˵Ĉ))0�*"m��s�H��&���(4�5��������ޏ�F���6���Bb�X�^�U!�e�(�!)IH�sLA�,^C�X	U7�[���g�DHS.�0?�ы����«D\�����`6��)�J��~�֪4�Rz���+3U��@2���-�5�����&S�%x��ԋP)�<�N�yt��o$�]�T��K_����>
��>%��:�?�]�"�*A�M�H�!�|�pڸt��e~�����-B��9�-7����"� �#���<��)]����i$����D7����©� � �����&��#�:Cױ9l���Xg��qf���[Yg�Q�wa�t�oΡ�Y��g�6�y���v���5��_�^Px\ÿ�/+0?��#�|(sG �y-��[ &a�euJ�����xu�f���S��p5�/m]�g ���I�bL�|fo4��3
YZ}!ы�w[#;�>�iux'۬���)4"��np�k�OL�<A�3��Z��,֢8��Ʒ�g��	=\��@�����`!S��Pf�L^���!�����	��Ղ��-���i�NS�Y`�ɚH>����}S�1I�p]�Rp���{K���A����Dͳ�He"뛘��C�ra���[>���4��-���w1�>�_M���}9�!'��k�����J^+�*�8�!#^vҷ���9jb�^-OI x*G&T�	ۋ�������� ��Jo2_=��]Ң��~;ښS/�r��	�0G�/39��Ͽ�2>���O:�lwj��R�j�_ac�H����Wy	�|��)Z�BW���$�a7	����^�\#�F.�u��0��KM����9��>.g�J�b>���Y�z�j��2O�}�d6��7�P�oB�� �T��r#{I��߼��Rn��N�	�"j_`��6���#nN5���%hؗ=j�|r�.j�k�� ��+ޠu?poi��7%>~�	�,���HƋ�ī�2�}-�h@�%X���^�x�:3��8�j61lh���ߡ|z�w�th����F�p�lo��6#ߝ��kz[��ʫ3="P��#��I�ώg��e����x��u��BN��U��y�wˑ4̟-<�����<| Ӯ��2�F�b�K3�6�L�6��9g�Y�__u�&�lw4#\�B�ɨ[qw�������7����+A��ʹv.˦�����e���ˠݪ��@u��[��4|i� k��a�N�\uZ����P�[��Lܕz�v��h���X�A�?-#�#��2��Q�=���$&����A�67����B���.�g���)��_zP+����7�c]��8�@�
�;�)C�>,���ε��wp�����<��>���Y�­�q0�&�UA���BA��E�>�*����zk���t���Ͱ�woBE-���������#�_��#vQ��³�aOo�;�Bn�Q׼�N/��V#5�?um\˯a�����_q����.�X%�+��+��ҙp�7�V��#��d1L\鷄��a,����\�L{v�h��^�ٕ�B�/��nƌ'���و�N�����GO1;�`fXtq�$��Br={���B�ո>$�|�H���F�� `��G'��z��ԛA�>)��/±�$2R 93<��3�e2J��ۑL��9-�a�h����2�;)5�V�(ty<�qu�<0��8����U�[��A�C�%m���#-�?cP�2N���L�|�e7��EIY�)M�A�驶�(�q�Q�	R���v��ît���'��v.Ŷ8#;R���93�a��s�yW;��0U���K�p��������z;�/㦋r���v0+�	�hf����	�V{(<�� nZ�t����O�m�k"�n7����RȒ[^�3'�u2Ӏ�	mm2�vh��_X�L����*�D�~�����v�ӣ7�y
�8P�`�i�0����j��?=�/+
3^sN�2�%K�}v��ǚHL����X���V�R���9")���ȋ�E�S���l�	$��WN	��Rxwӎ�Y���_��:�z��W�q��4;F�Xt:��c�Dw�e�|v�FSK���:�-NG������uE�;�@��+y�R�)��֓��\4���"��_�� �F�e��*�P�z���״杻�.k�� J��ۢ�z�D�S$I9/_S�ou���94h(�9��i�jm@!�c
����.)�=�����L]N��P��d)f�lyٔ-xdA�uQ=�0q"׏��n�~<cb������Rv�U��,W�-P7��\B��MRc��+e>�_��*��;��y�h��Y PG|��-֓��/B���H�����>p��J�	!g�ӕ������x��+�?��� ����������O$�kn`,�Ĩd�M�o@,B�����F�<\��9v��	-��q1�\��f��K��K��6�X^���F>fR�3/G���?��j_=��y�#�L��{.U��������#P����B9Έ��G��|�DF|�<O17w���ݬ���䀈�� Hl:��4?��*�.t.�*�T��zŴ`,�����ѫF�A�ҭ:�.�er�=Iի^kTW�3j-h�t9 �zJr_�0�����I��+���Ԃ�uz*�����K�Y�����������z�Õ)��$h�s�c�v�\�b=}�m~�ʭk��	�<�;Z4���'�Z�KY\�\��U�/A�z��ٱ���p�<�M��Uh�0	!�\��9;�����<�L�
/ 7�'��e�A���W:F�*,�R�V5���6���ˁ"@#�R5���A�sX=���%�馅S/��eύW$D�ax�0/�%(�B��Ծi�x,��"��R۸S�I��0IKq�J�R���-BF�_(;:���X�#9Q�a��#��}��F�����y6���ۛ~hY&[#��ԏ�7�M��}��(��X��lpe����M
����H�X� ��s���9���q�?'MV,I�~�!�B��V��ߗ���r�p��/��BˁU�#�4x�A׮·(,�h�mf����ݰRT��k�[3N��%7�Y��$���պ��	��ȳ���=���L�5djv<�*����HdVz������K�툥���g����3�hp���2�+��z/�nU�m۟tn��4���p(����������Kʘn�����zF��;tm��E	�'�ِ����'��k;�k/Oz�����]�cH�#\��b8�dԫ���k�?��<��2�&fxRX�$�:�����U��鰀�o�LRjG�n�Y]���{]�詩�t<Ӻ�o����U�9S{�:P������a(-R�$(�CD�R������Ās�>,��ܶwjb�˶��[��Ux`,��3C�<m����/����c� ���v��ej���3U�����ߠ�5�$�t��g���!����5yɮ��e _"$6��Z�cL�>�G��hf>��q	�}%鑰7Mñ^�	BG�g&[ F���!~��<ZC����w�YW������
CW=�U���~����=�:��Lϵ���ٕ�i&�;i��)�H��st+���Y!ba�����aZO�ƁtW�u+���Of��~gd.�S{�&�z���_��:3�dU6��4�MÝ�Z��oz!~"/��� Y_1�R�)|���C���^ˣ���W 4�r�3�k�Wb,D��\�h$ۮ7l������������<<�G��7�-�/Ů����j{+ʓV�oK#�.���� uE�ɯ��[cad<Ժt,3UR1�0���?b)�t�Pt�6��PW���а���3R��������?���(�.\Ns�z ���'+���������Ǫ���^��i��s�<����Z�:Z�g��wo	��G�Q���{��U���ӓ��(�TP���E����bS�\�;m@�>A�=��t�'->��t�X�W]2������Ǩȗ����G!O�ҡA;*�uI=�t!�'lF��ME����B����G4[D;!�˷SV�O�^��x9TpQj��'��vB��>�',���23I���Fjs <�aXHsjKY�Z��*s��nH��"����⒱+��CmU!�h�(�)�{������Y�b�i���K�\I7ҷ�O7~�x���0#(�A������v������g�#iE�c�N{^��2x�!2(�:���H(�ᲘJ��+�U�s��+�`��/)��Jwc�ʦT�:!p��G�uWf\�J�x�~�	$���?[u[�lΖ��3�a�t�4.?�wFZ���{* �cA&�9��Z�R�S��>�F����^�X㠥Y�&ke:�Je.�[��\;�,i����X�z}��CZ���������1g��
�)�����bV.����:��H��#]2���-@��L6A�!s`qj���[�G��6YC���g�fc ���.���S@hn;#�5Z���G)xrw?��]q{y�Jo�W����F�^:�r��\�G�����?������pe������ȫlM����>���w]�x���K:a�\L��-��?/n����aM���$�to �Ӟdjbv�� 渪�e�`�y�A� �.�i1DO8����wq-�Yl`ky[/�oeIf�m �����Α��+Y���!�h7��7��d�9ȱj��6��5��;E.���&wE���@T�裧��E�}��t��mGuW��~v �mR�o��$�k��))19FSnE��o�'�Ȉ:��x��F��{�Ir)�7��k��_H,��NTx:kCKsk�Y���.�^̌'��AU�C���#l-��d��ھP �=��PtC�G��D4���g���M?��?�o���Xa�~�1` ��������ǘ�Y�|xԦw��!o�X���x}���0޾G�EQcΥ�%�|E JG�;'��S���.u |;!'�k�8���x�>�uyCa��h']�!��K�r���1CSj>Y�E����ĵ�C��^������ҍg�׻�-�z����F<o<�2kK�j�	����45�i|q�jÝRN�~2��H��L�/F']qz����lp�cHn�]�rœ���ïykJ�|o�`�|E���
n�^���ټ6���u����7�:�Ξ�.o����H��&�rȱ�u���*��%g����+��ϩ�t��2g��j�^8����ӊ�)	��,!|����Nb�l��'R��gK�-��e�u,UV���(�?�M��V^{@��RLZ�P4H\��t����I�Y� 6�ȷ-��TkN.�L٣.?1Otd0k��?{���)iz�Cazׄ�-�<��+��������_n�a�s.缉�8qC��D��#����Q���Mu׊���;ǗR-���$7��-�a�S���-�RY���?���Y��6e����D[9�_)A�jⷷ8��j�(�-ٱ��U�����-�n�Y� (�9LG�3�t�.$E��;i��n�Y�&�w�_`�����j��$x�t]N���|r�dpa�[6Ǉ{__���u𡐵7M�ZК����2�8sUD?���%�8H���o
&F�s��(T���0&�{��Ӻ�:�b#yjHEZ�cI�nU������xb>+�7���N���;]"����-��l��}�Iyh��%2����=�=d�xibA�.yh���,�����e�*v��K�?��6'����/:�ʧ��"sҍymG��%�2�:��S�@i�I�n�h��kH(+�ωt�!�[����BȾ�E��AWgg0��Pз�|��/�^="jW���#ѻ��Y�)
�c]Z����ŦS���-j^����g�����)��D(����.q������5��->�_��{���A��U�l��Eՙ����zv� ��|�p���)��+$�v���/��M�.=�ȑ�Ϣ�AHG�I���tB���
���r'=7�eĚ���<�0ۢ-�!&����r�C��&�z���8:b>�B�#e���>�Z@����Aq�	�;��c�n�X�_�;�q3|��Cl0�B����*MP�}I`Դ�B��~ s�'ΤX�����+��2��y#���_.Aj^�=���iϭ��ߝ���*�D�������5����R����\������%ǩWA��󩤳~��&D,����ٳ)@e4/skӵj�2���L��%R�i�۳�g���5��HU߁el�8� �����V���1��7^�*��C���IjC�fÃgh���0�N:��.FP�0�p�sW>�o̮ᜏA>�����wQ|�cT��M������15$E�=wO�|�-�����l��q�b8�]��,����NG�;\9թ�b��]&u�JSÂ{A���f-	Bq� ��n �#Ⳓ���?�t�(ki]B��=�1�S�-���u!+�"�=��P�e l�[9,�
9�#`v�?8}7��3�u�(�e�oE|~�f��A��[�LA�.[�a*�d^�!I�y&��fG�v =J�X�!LU���GrM1`h�/�6�ʙ���D&=���	��$O�A���c�}�C�΢�nY�\c(���Ւn��u6"� �БZ�6�M��-$���.�5��?f�C�(�L[Խ�JZ�V]`�-q��P��.�C$(��/ߡ�x| ��C�)��g,��:G橻����,�Gh'=�/<&O("F�(��q[R�jm�`�t�������n�-�g^�;�y��C9�1����!��4t��(��*�4���
��j&N������Q��'�J[�	����/�-�-P��e�J�Cp���ćP���EJzGg�<N^�7S�i���S��"@)ƀ�c�&N}`@\YP�f.=2ySf(J��\hQ$�Z7�"Q+I.p���0c	�� �w�P.SF�W�rJ 2��ib�Yf���(��bmr���"g�K�D�u\�� �IJMIXG�(ebeX�N�"s[\�z��0�N+�~���\�.б�}��J{\��	<���@�͚T��x�0���k��b���+��t�hr]p=���J �j��&�p�.�N���EQ�([�A��do�o�{��<�[:�e.9���OP��#"|�CF撖n�T��²$i"pi�(S���+��'^����"J���R��<00��=x��9���|Jz����,A�Q"5�L]z�zO�{����f!���N˼�TX�������'H�y!k" 8.�ӂ�D�w�N�w"
�4�𦛩�d�Κ�I��6I~�D݄ZP�o=lv�f5rP���Q���B7�a2θ��ռ��
S^j(�1�ZK��������宾��W�5XDK�!�[����w���x]�ӞW� i.h��+2~Vr<0P��n�I�v³��u���1W���ᤔ/��d��c5��1��ƺ���a��C���++Ii�B�Q�5D�#�A�eLXH�@ĺ��X$���2�h4��<*�S����V�E�̜h�S	{����ݺ^�/��AJ���.�4	�6V��Bpe�ib^g
j�����
���b����Ԥ��f������^��`�+��۩���_뼎��I�R�mA���M8Ek�q����/_Q��1����N��[�Ҽ�\� �05�@�������y��N��Mo��|��^8č������p��M@��	HyX�ik'�	���8��e���;O7�@�%��o�*?�P�h���7�Ȋ}e�;�R2_��l$����,-�<{��w(��;0���u�܃���l6�����jh4��N�s2���n�Ǎ�;
�O3w f��EO� brď$~��&���ې�U[�&�Z������j��M����5��H<��d�J���ϙ��p� �ĩL�HM�����Vp����<q�"�`���`'�v���V޼ㄤ����0 �mÁ�X����B˧2�����1�ἃ��K~?g��edꋣ{g��ɵ��{L�%��q�<b�E/"ytI���ʷDg���b��Bc D�A�@}�'1��X0�}�ߝ��i�����̺���\�PN������pu̽����aX�V��"n�aB���@�)j��|�BQ��=R`��¡$��~x�/o�9�3�d�؊oPE��9��~a�!y�����r�-���W���I�ÙS20���Z	����}��Ĩ��pA�t�3�2�I�!�?÷���#^��+�+{ja!�,"�m�?�=(w�1�N����B����$ck�������盂�����R�gW��֥�=z������?�fc
T���^!�*X�3�_V�YD��GOE��e�3Vq7�B����	T��|�9��3����^�҄p�z�Ӗ�����><i��W����>D��IҤ�ꨳnT5Aj`i�p���� ��M�@��a_b���To�2RJ�"�.*�YA�1x�SP��5��ir/�;5�4����w~Rv��F��+��5�����7濆�QsH#�Ǡ�lG���â�����W/�-F���hb^�SuRE���OߙM��N	 t�����?s���o9�9��559���b/��=���86x7��{����N�gW[svu��q�2k��k���ݥ�a��,Y��'�"�-t�G2e�Ԅ�m�bX���=Y6M�#UT�?�	3u��cr��x��Â�}\}�Z���Ih�T_�,����4ĕem(��^���[�8T��G��Y4ym���a:k���ֈ���7ZJ���e���IkG�)3I׻�T"Q|��+,�`9A�`3;J;7�E-��M�~��P*BNbI8m4�����C�A�6ҵ�
�֫� �/��%�/v?�.ڂ�x���6�V����Lr"�Pg�;�;��Y1���V�:��ײ8�2�n\U%�mv�[P9e�Gi�d�Vv��w�+���6=Y�l��f�x�,p�r����y���>T�Odc+$�db�'�^��c�[$��ʳ���wH�62�
��	��^�%?�TV$���z�-�:;9���&�0Ğ-��;r��n�s)�	e��Z�h��[.s�Ƥ�iy%��/�kS�7��=�(��<�˧^0�SiH�z���u �y�K���*f�c�D[�rDj>(�z��Z���
��/����41�?v�P�e�R�/�|��@ �-�)��/��L�G�@��>��8���}l��!��݊w�>�G��0��w���AUc�I��!)�/fA���5!;z��B����.x����m�hN'X�e�Z:h�;j��n�Aj�9:[�7sِ�H;�������nk���\��:��2ɿ�)T�vZx�����um��vW��4��E�,\Y� |`�]51�>c�G��6�>㑐;��U�'��ӗ�p���ND1B3;�D��
���8���T�%)�8��í�:̶byEw�K'WT��k�A�*:���c���VS˫_{�M���k�P�y�xaYGY�5 �8�˜D;�E �X��h�a9s��No�p1hZ[iw�R�K�i|]��|?ׂ�:�@�ؽ�4ы��zwr��R�!�fN��y]n%^�D��p��^{���z�5R���&��!M]ЀGE_�/TS�c��6����`j��j��)��x�s���,a\Ⱦ
���Kb���_2��ő.���ޢh�̧�3�<�"J}E~ͻ>���G�H�?����s��+M�4@g�2F�9^��eRS��!��bq+u�&aE�ۘrh炡���ӯ���is�k갲�uh���0��"	6��`�P����]~��k��5Qd��;����Җ��~0UI2�W2��7 ��>�Q��@�)[IUu�Wa��������;�����ǯi1�%
��na#5],5_O^��I���,�|��:gQ�����~4��<�t������+n�p�J�(ѥ^kҒgK���!��G]��6�ylHֶ��m��C�����0���A�c_�qaŎTʊ�i������9L���#Ԍ�a���%]�!~L^A�G.w>)�ɮ��������ː3X�������-ߔ���+8�!L�]�g�����/���YS2� ��!�R#����-�� �w�OK�p4��5n<�zΊ����H�g�1o�I����ר�U���\��X8�9�r���.��JJ�A�*<T�6�/l�"�*���{y�!'�\Tbј�!���y�2��ۧ��[�y���,��y��n���G6d6����vk�i����?N�9�g�UR
�A	j��cj�C���]�qY8B�C�x����E��k9zӹ���'�EG���4���{ν�2�sL�6Q/_���Ȟ/�h2��^��H����!��[������cp�<6%�RFi��B��ba�Z>�]h�$�F�(
�s��d�3� �t.�8!-��2��;�V�)������j�e}�
̃�l1c�Q����8�=��ʆ�-z�h�)�K��u��h��A;GN�e������LY�<νO�c����w&���R��� ��&&I��DӅ}*0�խ�sFf��PX��#!�@�%��k����h�_y�04�x�f��AJ�������r�o�$��礹1l��G�p�I6���T'%`��ӺT�L�vKlW���
E��.�cO���N$Zp���f�-Q��ߍ�;�8X�icI�q���q
Yh�]2�j���5H�C���
b��*���#@�ސ-�Z�G1�R �?}��B���	.퍦9'"�������/ ����G~�c����K;A$.@2�;���O۝N�p�v�Z����uۣ��,E�Dp#"U趚s�1�����%���oS;>]�-n�� �Ge���q��+���Z�[�Bh7�ꎜ�y;Q��j�7�<q�T]D�l�=O�
�=��bH��Y���y��1,�jaa��פ)�|
�&<'�0 �ʔE%Q����r�͕E�Be#H�oˊC���֪�}�؈�XH�G�E=]`����(���Ŀ����5�xMq���mQ1"��c�׋i�tF'����V[��u(��D���P�wގP�\-��w��äu�쎔/b�~���e��@�C�;ܖ��P+ڨP���ً�`�^�p�{��o��i�://��an��,Q���ö��D�3���F5bR;Gݨ줯�I������"{�xM�2��T/7~�kz��N/����e��9{ɓy�m�L;�GA2�ibd�'����KF�����8��&�J�%(��x@}��/ŐS�����Z,�����3�`����C~X�^�6���������>��E��F=�N�C<k�՚L!_sx�!��	���p�����N�S�y�8�@R�@�v��(n<����4XV�l $�v�U6�A�;ʘwǈ��	��s�L��:0e�]p����ע{�}.8��">�r)�0[.
Δ&{�:���(d>���|��nK�A_糁��e35��I�D��~�NqD����L��Wt<���ktP��"�5�m1��*�����e5ǔXq�<��X�2��ǌV7�fz�f���@W��R_���"��/?G�$%~
[XC�пl�
Ib�C@9|�4Ta�%<пpC�S�^x�\=쀺��`����<��.碗��2��~�~VPZ6k9��j^�cp��^(�煜)GRyd8Ԍݖ�M0+�c:9��� ������R�E���f:^�����4�/��o=DR���軔%��`�a��ToI5�!�}��:��-q+[�+���ڭv�k�}��[Dr�r6�����˼qZ�F�u,���*�q@�����Kn����T�p9u�b��8L"���R5J�/�;�b��CO�P�f�8���# ���c��k�v��*%�F5�Q"Jx����z�G�H,K��>$����Պ+�C.��c���seSN&���߽tF�@� #�o���v�N��pՓ���/G�q調§�ce�������S}I��uY��
m�h:�7��0��M���W�yM<~��:Ry"�f3Ra4܃5���R~�uo��M��vN�{�2����yÌZ�[��?QDss�*	V�Qt�(��,�/�&�k&�����n�.Ê���H�=���E�f+|%>(-���˽����倍��:�5��w����^�&/8ۈd��w���+O�@��P�ݿ�h*`,3� �1⥫"N����F������5�I�wj3[��۞�&vPnP���o��e,~9��J"��N:�>d������\��p7�nh�/)��r֞�M���6��J^T��~���vپ�f�zb�o�(���/z���!N"1�%c��wP:{��'�m>o�ޑ��\K��"��?��*��LK	��U{'�͞�O|��_Z��|�f[��8�'���iC��d�k���� ��X��26��Y���\�w#F�����^�:���u�QY��NBl�PZ;�#]���<�9��=H1u'����UX��*Je�׎Ǆ��	�b��M1��
��-9�I�f*TX�èv���y�U�8�i�Ԙ����g��䣇xM0E��ya�k��8�d��q�=��<���:�M~�YB~l?x��� ��O�����b�����揑�p�f'�5U��~�!�[;N�{U��P�T��#�-��ɧW2���aD��x}s��������N����J9ZP���ѴN� m��L�� �K>������2�����J���2;���vA���c:j�[�S|tnyՄ����צ��(j*:@�����xϓȱf��5N�\1��� <�V�^� y��PX��_�=�ĥ>[{O݂]���-��q�_������l�����q*��F�ե�9؏��	��O@��2r9P��
�,2��r��C8Q�f���ɋG��	&��⤜�$���K���e��|�R�+����)NuY5+g�(&��o�I��c���������aeݦxx���M+h# ,u��Ƥ��S�|�63�`~��\p/բ=}"�Zl�:� �I�=a���Jj�f�����Xf��]c��|���Ja!4t��"1��z`��A��{�ڏ�!�'}�&ϛ�Vl>���%�d@����/�0�)�2f�xH>��&pQ����W8B\�M���ESP�	,��j8��`��`�B��s�ڥ摫���(G�u�C ��c~�m�����ݍ�����G�_�+�����0�}N�;]Q���^ԝ"+S��U\o_i%MX�T����T�O"��D ��)���m��e�kyb&d_�Z�s�}��������4�P�t:�*?���P���n��z�[�t�.��l�����V�t�j�,��o@e���^4�� ��_l��}�'j����i����G u.|,K��t�ɳN�I�m�U:3r�/��7�J�t7![tx9�{��1?�&���%�%0�p��{��"�xK3��>�RihW�N��F& R�>�}��)"�O��k��D2�9<��Y�!������F'�s�������2cS??��I	�ً�n�F4�`M�������t���<� �	�B�����#�&NPC )�#=�hH���J3���������F6u�vo����&^+`�u���p%Ma��l�<�&�e�g��_�����aј�����N�\��j�+2�N���8/x�ݺ�ѡD!��E@��h�8��rQ��̯�K��ͮ��H������ɐ������`O ����TP����7}�r1����`���喲x�j<sK����J)�l?�^7PE/�q؍�C^�S��� ����Aln�[�z��dґ��]}�@[gg����@a��^@��*G�
*���\�!왶�Y�.�0]N瞈ʟ@+��n\8ˉ�~��!� ����ln����\��M[c0��G�����wB�j�!IY��7\4��N��cُ����̋;���~������9T�J�[i���w4���+iF�צ�}P�������Z�^M+lB�y��\�,w�}��f�/e ��>bٍ[;�8>쳥�Ռ䬐?��'Ӻ.B��z4]le���3�n4���y��7]&-�Hl���v�͊ i�jӐ����?9׌g��d�q^�c�bsNu����c�9�%�1�}vΊ"�a��K]�(�ix�����$JOÜ�2ͻ�cd�"�����Mb;6v�k�Z�?��p�L���n���J����NT��x<ՙ���&uEP��Th�L� ^'�R\lA.�ߨ�; 3c��bY�wAϫ!��-�d��b��	K��<�'�Y-f���@'��^�"v��ӑD�FW���t��c���e8)?0ہނ eZf9TX�ߘ</ f�U�Pe�P�uDJ`na�Ý;zB�m#�`6���MJ;1Wϲ-r������	��Ԃ,��(�W��4 FS�ʄ 匴8[�@o�ָ�c�!Q���`i�+�a�,�$�-��t��<m�	/�-jf��K*�ZO���c",�->q6�-m�����Z�-�='�ڑGհ'¢�'a'^^Z�1���Y��|���F�
R�ӘܬvW����ڋSy*%>
<X��W����,�ZU�hx�!S����u�oIA��m��^h�@�D!V�K�%������>�)�~¼S��9�<��&@���>��rgo[B��r
�Q��\%�F.�~N4Z�Z��9��V�(�+ .����gu��mI�>Uz��i:.w�B�����Zh�0ށP���X����6�7r�h'�G���\�%V�c�|��L������ʺ�Ł�.E������AD�ޗ��H˽Ȋ�H�l�?���֪�����Ob�ui�TVI��e��B����w�.N�0(�SS^���>����P˻;�N����iѮ�.����W3����{��a�p�+�Kŭ^J�p��<����U�����Ue�uHZ�脆����Y�9�J�|rw/��w0*������(1��Ĭ�@x�CN���y���TW����l�4�T>�?b_�=��u��/��'Z[��a�������^��1� �$�u|n��a�|���ʨs��ѭ]W|�}�v,�
̩KӴ�/����_�r"��0#Q�'2����P��9�x�����3�����gL]ihs�{�2K�`�3gt�oc����y)�};�LW{J�g��H]����B�xi�4ɓs[;�3L�Y����Ԝ�Z�N:g�4��vo��ÂDs�z���Gjy��n�ՅQ^)��I�y����l*����ğA�M�[���R�T!v������w6==W�;'�t���(]��Z�q��
�Z©�=����E�(̰�܁4�Ec�V���O��1�.7�+R{Tu��MhҸ{�:�Nj��tʪV��`,�͙4�HE���e�3����\֤S1/e����_�`�o$M��C��f:��X�Jwh�e��[��"����=���_JzaL�7*(ˀs�J�v�漑]�r��D<x����)����`WCmF�f]�6e�Ŵ�}ķ���Y'�w�є�>���8Ǐi��}�|�@&?g�J�X�(�y���/��� �:���H�<o�Z���s.l�� E$,�)�����ߔ��$��?��|��r=�g��H�ʆ��8��9��ˠN�#\�˶���x�?*VT�(_��y�����} ���f�����%=�%���8v�k	� 6�q| �L���d�t��
ԃ�-���x�����_������v�̴`�T�LƷZ%��7�oХk)] {��Ba�ɡ>1���( f���
�N��a�::��������v��N �I�U��YI�>�o�#T��`N9m�}����Ka|�铫�]}'&��w��6|>Vxw��?e��B7��)ëD��� ���*!��ڇA�O
�.�ڄ��.َ��'?9���g�dY�_%���Q(�j=E|�#]��9Oӛ�������:���;� _�p~' �tZM���<���Y�`b\���;��?#t�r�B,n�Z��qYN(L�t�G)[�b_GZ���n�͵�f�OR|H�4[��t$o��L>:��9«y�#9�Q-����U�l�da�~t�-mtr]A����P\uc��4�U6�xs�3<AĹ���G˄$�EO�Z��(�r���C	q�I���	 䏅Z8�C,���*��4�4���m��4�
3:��>�5ۥ��(r�7��`��r�LR��6K,M��=Q�B���G<Vd��r���nT`;�CD��i4Bz����B;�44��=w�b6*M$�+��Ĕ��[ �1��=E����zPh����+���[�22����_z_Qs����y����֦�������B�C���f�&t�����P�j���Qu,,+�ٟ�Z�:Ed�rH0i��B���cW���I��I2qnus?Z�����T���/mb���q��0$�&�2bD���d~��$������,��@1���dS�P�J\T��|6���ğf��uo\��KAů�ݩ�Ad<Tn:���8��\��vU�E׊�!*!�75м�^��n�V�FC�/��s��� 2���&�p��F�",3�/�'��H��}�M(��ۋ�����:x;s*�����$����V��RP��$�e�ߢy�m�LH�(�<�Bv�����g�i|�p��E ���i��� �4#9���&es Q����ܥq�N��[�iR�h��S_�����+̬�����䕞�c!P�DU\�N�]蒆C�U���4O���h�bؾm�#"�1�#�����C륖yH��������I}S!,�(#�U�u��]6�=`vV�����f�Q��7��`tX0U����Ŵ��Ȋ���kV�.��.�x@`���?�3��G<�+2S�@h΂i-��vk]e��@6.l)����3|�s[�x,{�A(/1���vN����[{-�[i�����:X�t�<�	��>4���n$�%���q�o���u�1g3��w�I�[�-	C�;'	�4�����p�wo�}hC��N��L`�����|��`�i�~M-��ts˴�U��<�Պ��Ȑ�u�@sp�+�l�0�F���d�A��dq�1�{�O1>yeS��}ّ�F7k0�3oeB�gʠ8j�ӣ[������M�L���݄3\�ޒT�r�"�E6NoD=��^�U�~�r��vλ������y��,;� �qOl�R��ܠ§��OO�ڙ��H'���<l��+Jr�{��\�{FF JG��2d�������M"��?������Qq�AY�~(��R�Jv�?Ŷ�jn���g4� �X��q�la�3tv!ڈV7{����@��}S*���b������_B��$_�Zv��S�F���ʂ�W����$���/���iڈ-X�q������t������8N�����WLҒ���"�������F�e���鯐��\%6��G�V�:�SӟC�1��`]G���Woʘ��Cv�Ns3�Q��wq������e�=���߆��ش�7��2�